//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 0 0 0 1 1 1 1 1 0 1 0 1 1 0 1 1 0 0 0 1 1 1 0 1 1 0 0 1 1 0 0 1 1 1 1 0 0 1 0 0 0 1 0 1 1 0 1 1 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n709_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n751_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n861_, new_n862_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n869_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n904_, new_n905_,
    new_n906_, new_n908_, new_n909_, new_n910_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n920_,
    new_n922_, new_n923_, new_n924_, new_n926_, new_n927_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(G141gat), .ZN(new_n203_));
  INV_X1    g002(.A(G148gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  OR2_X1    g004(.A1(new_n205_), .A2(KEYINPUT3), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT2), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n205_), .A2(KEYINPUT3), .ZN(new_n211_));
  NAND4_X1  g010(.A1(new_n206_), .A2(new_n209_), .A3(new_n210_), .A4(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G155gat), .B(G162gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT90), .ZN(new_n214_));
  OR2_X1    g013(.A1(new_n213_), .A2(KEYINPUT90), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n212_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(G155gat), .ZN(new_n217_));
  INV_X1    g016(.A(G162gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT1), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n219_), .B1(G155gat), .B2(G162gat), .ZN(new_n220_));
  NOR3_X1   g019(.A1(new_n217_), .A2(new_n218_), .A3(KEYINPUT1), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n207_), .B(new_n205_), .C1(new_n220_), .C2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n216_), .A2(new_n222_), .ZN(new_n223_));
  XOR2_X1   g022(.A(G127gat), .B(G134gat), .Z(new_n224_));
  XOR2_X1   g023(.A(G113gat), .B(G120gat), .Z(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n223_), .A2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n216_), .A2(new_n226_), .A3(new_n222_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n228_), .A2(KEYINPUT4), .A3(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G225gat), .A2(G233gat), .ZN(new_n231_));
  XOR2_X1   g030(.A(new_n231_), .B(KEYINPUT95), .Z(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n226_), .B1(new_n216_), .B2(new_n222_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT4), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n233_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n230_), .A2(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n228_), .A2(new_n229_), .A3(new_n233_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G1gat), .B(G29gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G57gat), .B(G85gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n239_), .A2(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n237_), .A2(new_n238_), .A3(new_n244_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT23), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n249_), .A2(G183gat), .A3(G190gat), .ZN(new_n250_));
  OR2_X1    g049(.A1(new_n250_), .A2(KEYINPUT83), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(KEYINPUT83), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n249_), .B1(G183gat), .B2(G190gat), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(G169gat), .A2(G176gat), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n256_), .B(KEYINPUT84), .C1(KEYINPUT24), .C2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT25), .B(G183gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT26), .B(G190gat), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT24), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n262_), .B1(G169gat), .B2(G176gat), .ZN(new_n263_));
  AOI22_X1  g062(.A1(new_n260_), .A2(new_n261_), .B1(new_n263_), .B2(new_n258_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT82), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT84), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n254_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n258_), .A2(KEYINPUT24), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n266_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n259_), .A2(new_n265_), .A3(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT22), .B(G169gat), .ZN(new_n271_));
  INV_X1    g070(.A(G176gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G169gat), .A2(G176gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  OR2_X1    g074(.A1(new_n275_), .A2(KEYINPUT85), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(KEYINPUT85), .ZN(new_n277_));
  AND2_X1   g076(.A1(new_n255_), .A2(new_n250_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(G183gat), .A2(G190gat), .ZN(new_n279_));
  OAI211_X1 g078(.A(new_n276_), .B(new_n277_), .C1(new_n278_), .C2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n270_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT30), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT88), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT30), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n281_), .B(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT88), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n284_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G227gat), .A2(G233gat), .ZN(new_n289_));
  INV_X1    g088(.A(G15gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(G71gat), .ZN(new_n292_));
  INV_X1    g091(.A(G99gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  XOR2_X1   g093(.A(KEYINPUT86), .B(G43gat), .Z(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT87), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n294_), .B(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n288_), .A2(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n298_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  XOR2_X1   g100(.A(new_n226_), .B(KEYINPUT31), .Z(new_n302_));
  NAND3_X1  g101(.A1(new_n299_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n302_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n297_), .B1(new_n284_), .B2(new_n287_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n304_), .B1(new_n305_), .B2(new_n300_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n248_), .B1(new_n303_), .B2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT102), .B(KEYINPUT27), .ZN(new_n308_));
  XOR2_X1   g107(.A(G197gat), .B(G204gat), .Z(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT21), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G211gat), .B(G218gat), .ZN(new_n311_));
  OR2_X1    g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G197gat), .B(G204gat), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT21), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n310_), .A2(new_n315_), .A3(new_n311_), .ZN(new_n316_));
  AND2_X1   g115(.A1(new_n312_), .A2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n270_), .A2(new_n317_), .A3(new_n280_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n261_), .B(KEYINPUT92), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(new_n260_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n263_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT93), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n257_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n323_), .B1(new_n322_), .B2(new_n321_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n278_), .A2(new_n268_), .ZN(new_n325_));
  AND3_X1   g124(.A1(new_n320_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  OAI211_X1 g125(.A(new_n274_), .B(new_n273_), .C1(new_n267_), .C2(new_n279_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT94), .ZN(new_n328_));
  INV_X1    g127(.A(new_n279_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n275_), .B1(new_n256_), .B2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT94), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n326_), .B1(new_n328_), .B2(new_n332_), .ZN(new_n333_));
  OAI211_X1 g132(.A(KEYINPUT20), .B(new_n318_), .C1(new_n333_), .C2(new_n317_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G226gat), .A2(G233gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT19), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n336_), .B1(new_n333_), .B2(new_n317_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT20), .ZN(new_n339_));
  INV_X1    g138(.A(new_n317_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n339_), .B1(new_n281_), .B2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n338_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n337_), .A2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G8gat), .B(G36gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT18), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G64gat), .B(G92gat), .ZN(new_n346_));
  XOR2_X1   g145(.A(new_n345_), .B(new_n346_), .Z(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n343_), .A2(new_n348_), .ZN(new_n349_));
  AOI22_X1  g148(.A1(new_n334_), .A2(new_n336_), .B1(new_n338_), .B2(new_n341_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(new_n347_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n308_), .B1(new_n349_), .B2(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(KEYINPUT101), .B1(new_n334_), .B2(new_n336_), .ZN(new_n353_));
  OR2_X1    g152(.A1(new_n333_), .A2(new_n317_), .ZN(new_n354_));
  AND2_X1   g153(.A1(new_n318_), .A2(KEYINPUT20), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT101), .ZN(new_n356_));
  INV_X1    g155(.A(new_n336_), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n354_), .A2(new_n355_), .A3(new_n356_), .A4(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT100), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n359_), .B1(new_n326_), .B2(new_n330_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n320_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n361_), .A2(KEYINPUT100), .A3(new_n327_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n360_), .A2(new_n317_), .A3(new_n362_), .ZN(new_n363_));
  AND2_X1   g162(.A1(new_n341_), .A2(new_n363_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n353_), .B(new_n358_), .C1(new_n357_), .C2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(new_n348_), .ZN(new_n366_));
  AND2_X1   g165(.A1(new_n351_), .A2(KEYINPUT27), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n352_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n317_), .B1(new_n223_), .B2(KEYINPUT29), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G228gat), .A2(G233gat), .ZN(new_n370_));
  AND2_X1   g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n369_), .A2(new_n370_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G78gat), .B(G106gat), .ZN(new_n373_));
  OR3_X1    g172(.A1(new_n371_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n373_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n223_), .A2(KEYINPUT29), .ZN(new_n376_));
  XOR2_X1   g175(.A(G22gat), .B(G50gat), .Z(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT28), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n376_), .B(new_n378_), .ZN(new_n379_));
  AND4_X1   g178(.A1(KEYINPUT91), .A2(new_n374_), .A3(new_n375_), .A4(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT91), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n375_), .A2(new_n381_), .ZN(new_n382_));
  AOI22_X1  g181(.A1(new_n382_), .A2(new_n379_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n380_), .A2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n307_), .A2(new_n368_), .A3(new_n384_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n237_), .A2(KEYINPUT33), .A3(new_n238_), .A4(new_n244_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n228_), .A2(new_n229_), .A3(new_n232_), .ZN(new_n387_));
  AND3_X1   g186(.A1(new_n228_), .A2(KEYINPUT4), .A3(new_n229_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n233_), .B1(new_n228_), .B2(KEYINPUT4), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n245_), .B(new_n387_), .C1(new_n388_), .C2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n386_), .A2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT98), .B(KEYINPUT33), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n392_), .B1(new_n247_), .B2(KEYINPUT97), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT97), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n237_), .A2(new_n394_), .A3(new_n238_), .A4(new_n244_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n391_), .B1(new_n393_), .B2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n396_), .A2(new_n349_), .A3(new_n351_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT99), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n396_), .A2(new_n349_), .A3(KEYINPUT99), .A4(new_n351_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n347_), .A2(KEYINPUT32), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n365_), .A2(new_n402_), .ZN(new_n403_));
  AOI22_X1  g202(.A1(new_n350_), .A2(new_n401_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n399_), .A2(new_n400_), .A3(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n384_), .A2(new_n248_), .ZN(new_n407_));
  AOI22_X1  g206(.A1(new_n406_), .A2(new_n384_), .B1(new_n368_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT89), .ZN(new_n409_));
  INV_X1    g208(.A(new_n306_), .ZN(new_n410_));
  NOR3_X1   g209(.A1(new_n305_), .A2(new_n300_), .A3(new_n304_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n409_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n303_), .A2(new_n306_), .A3(KEYINPUT89), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n385_), .B1(new_n408_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT8), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G85gat), .B(G92gat), .ZN(new_n417_));
  OAI21_X1  g216(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NOR3_X1   g218(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G99gat), .A2(G106gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT6), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT6), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n424_), .A2(G99gat), .A3(G106gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n423_), .A2(new_n425_), .ZN(new_n426_));
  AOI211_X1 g225(.A(new_n416_), .B(new_n417_), .C1(new_n421_), .C2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT7), .ZN(new_n428_));
  INV_X1    g227(.A(G106gat), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n428_), .A2(new_n293_), .A3(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n424_), .B1(G99gat), .B2(G106gat), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n422_), .A2(KEYINPUT6), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n418_), .B(new_n430_), .C1(new_n431_), .C2(new_n432_), .ZN(new_n433_));
  AND2_X1   g232(.A1(G85gat), .A2(G92gat), .ZN(new_n434_));
  NOR2_X1   g233(.A1(G85gat), .A2(G92gat), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(KEYINPUT8), .B1(new_n433_), .B2(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n427_), .A2(new_n437_), .ZN(new_n438_));
  OR2_X1    g237(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n439_), .A2(new_n429_), .A3(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n441_), .B1(new_n417_), .B2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT9), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n434_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n426_), .A2(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(KEYINPUT65), .B1(new_n443_), .B2(new_n446_), .ZN(new_n447_));
  XOR2_X1   g246(.A(KEYINPUT64), .B(KEYINPUT9), .Z(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(new_n436_), .ZN(new_n449_));
  AOI22_X1  g248(.A1(new_n423_), .A2(new_n425_), .B1(new_n434_), .B2(new_n444_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT65), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n449_), .A2(new_n450_), .A3(new_n451_), .A4(new_n441_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n447_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n438_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G29gat), .B(G36gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G43gat), .B(G50gat), .ZN(new_n457_));
  OR2_X1    g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n456_), .A2(new_n457_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n455_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G232gat), .A2(G233gat), .ZN(new_n462_));
  XOR2_X1   g261(.A(new_n462_), .B(KEYINPUT34), .Z(new_n463_));
  INV_X1    g262(.A(KEYINPUT35), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n461_), .A2(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n463_), .A2(new_n464_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n460_), .B(KEYINPUT15), .ZN(new_n468_));
  AND2_X1   g267(.A1(new_n454_), .A2(new_n468_), .ZN(new_n469_));
  NOR3_X1   g268(.A1(new_n466_), .A2(new_n467_), .A3(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT73), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n466_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n461_), .A2(KEYINPUT73), .A3(new_n465_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT72), .ZN(new_n474_));
  OR2_X1    g273(.A1(new_n469_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n469_), .A2(new_n474_), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n472_), .A2(new_n473_), .A3(new_n475_), .A4(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n470_), .B1(new_n477_), .B2(new_n467_), .ZN(new_n478_));
  XOR2_X1   g277(.A(G190gat), .B(G218gat), .Z(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(KEYINPUT74), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G134gat), .B(G162gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT36), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(KEYINPUT76), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n478_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n482_), .A2(new_n483_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(KEYINPUT75), .ZN(new_n488_));
  AOI211_X1 g287(.A(new_n470_), .B(new_n488_), .C1(new_n477_), .C2(new_n467_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n486_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n415_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(KEYINPUT77), .B(G15gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(G22gat), .ZN(new_n494_));
  XOR2_X1   g293(.A(G1gat), .B(G8gat), .Z(new_n495_));
  INV_X1    g294(.A(G8gat), .ZN(new_n496_));
  OAI21_X1  g295(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n494_), .A2(new_n495_), .A3(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n495_), .B1(new_n494_), .B2(new_n497_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G57gat), .B(G64gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT11), .ZN(new_n503_));
  XOR2_X1   g302(.A(G71gat), .B(G78gat), .Z(new_n504_));
  OR2_X1    g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n503_), .A2(new_n504_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n502_), .A2(KEYINPUT11), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n505_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n501_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n500_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(new_n498_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n508_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  AND2_X1   g312(.A1(G231gat), .A2(G233gat), .ZN(new_n514_));
  OR3_X1    g313(.A1(new_n509_), .A2(new_n513_), .A3(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n514_), .B1(new_n509_), .B2(new_n513_), .ZN(new_n516_));
  XOR2_X1   g315(.A(G127gat), .B(G155gat), .Z(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT16), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G183gat), .B(G211gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT17), .ZN(new_n521_));
  OR2_X1    g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(new_n521_), .ZN(new_n523_));
  AOI22_X1  g322(.A1(new_n515_), .A2(new_n516_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT78), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n515_), .A2(new_n522_), .A3(new_n516_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n525_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n527_), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT78), .B1(new_n529_), .B2(new_n524_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G113gat), .B(G141gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G169gat), .B(G197gat), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n533_), .B(new_n534_), .Z(new_n535_));
  NAND2_X1  g334(.A1(G229gat), .A2(G233gat), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  AND3_X1   g336(.A1(new_n458_), .A2(KEYINPUT79), .A3(new_n459_), .ZN(new_n538_));
  AOI21_X1  g337(.A(KEYINPUT79), .B1(new_n458_), .B2(new_n459_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n537_), .B1(new_n501_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT80), .ZN(new_n543_));
  AND3_X1   g342(.A1(new_n511_), .A2(new_n543_), .A3(new_n468_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n543_), .B1(new_n511_), .B2(new_n468_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n542_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n501_), .A2(new_n541_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n511_), .A2(new_n540_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(new_n537_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n535_), .B1(new_n546_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n546_), .A2(new_n550_), .A3(new_n535_), .ZN(new_n553_));
  AOI21_X1  g352(.A(KEYINPUT81), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n553_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT81), .ZN(new_n556_));
  NOR3_X1   g355(.A1(new_n555_), .A2(new_n556_), .A3(new_n551_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n554_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT67), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n508_), .B1(new_n438_), .B2(new_n453_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT68), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n559_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  OAI21_X1  g361(.A(KEYINPUT12), .B1(new_n560_), .B2(new_n559_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G230gat), .A2(G233gat), .ZN(new_n565_));
  OAI211_X1 g364(.A(new_n559_), .B(KEYINPUT12), .C1(new_n560_), .C2(new_n561_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n455_), .A2(new_n508_), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n564_), .A2(new_n565_), .A3(new_n566_), .A4(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n565_), .B1(new_n560_), .B2(KEYINPUT66), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT66), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n567_), .A2(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n569_), .B1(new_n571_), .B2(new_n560_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G120gat), .B(G148gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT5), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G176gat), .B(G204gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n568_), .A2(new_n572_), .A3(new_n576_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n568_), .A2(new_n572_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n576_), .B(KEYINPUT69), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n577_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT13), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n581_), .A2(KEYINPUT70), .ZN(new_n582_));
  OR2_X1    g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n581_), .A2(KEYINPUT70), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n580_), .B1(new_n584_), .B2(new_n582_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n558_), .B1(new_n583_), .B2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NOR3_X1   g386(.A1(new_n492_), .A2(new_n532_), .A3(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n202_), .B1(new_n588_), .B2(new_n248_), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n589_), .B(KEYINPUT103), .Z(new_n590_));
  AND3_X1   g389(.A1(new_n307_), .A2(new_n368_), .A3(new_n384_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n406_), .A2(new_n384_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n368_), .A2(new_n407_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n412_), .A2(new_n413_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n591_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n583_), .A2(new_n585_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT71), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT37), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n599_), .B1(new_n486_), .B2(new_n489_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n488_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n478_), .A2(new_n601_), .ZN(new_n602_));
  OAI211_X1 g401(.A(new_n602_), .B(KEYINPUT37), .C1(new_n478_), .C2(new_n485_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n600_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(new_n531_), .ZN(new_n606_));
  NOR4_X1   g405(.A1(new_n596_), .A2(new_n598_), .A3(new_n558_), .A4(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n607_), .A2(new_n202_), .A3(new_n248_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT38), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n590_), .A2(new_n609_), .ZN(G1324gat));
  INV_X1    g409(.A(new_n368_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n607_), .A2(new_n496_), .A3(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT39), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n596_), .A2(new_n490_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n587_), .A2(new_n532_), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n614_), .A2(KEYINPUT104), .A3(new_n611_), .A4(new_n615_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n616_), .A2(G8gat), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n614_), .A2(new_n611_), .A3(new_n615_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT104), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n613_), .B1(new_n617_), .B2(new_n620_), .ZN(new_n621_));
  AND4_X1   g420(.A1(new_n613_), .A2(new_n620_), .A3(G8gat), .A4(new_n616_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n612_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT40), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  OAI211_X1 g424(.A(KEYINPUT40), .B(new_n612_), .C1(new_n621_), .C2(new_n622_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(G1325gat));
  NAND3_X1  g426(.A1(new_n607_), .A2(new_n290_), .A3(new_n414_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n588_), .A2(new_n414_), .ZN(new_n629_));
  AND3_X1   g428(.A1(new_n629_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n630_));
  AOI21_X1  g429(.A(KEYINPUT41), .B1(new_n629_), .B2(G15gat), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n628_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT105), .ZN(G1326gat));
  INV_X1    g432(.A(G22gat), .ZN(new_n634_));
  INV_X1    g433(.A(new_n384_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n634_), .B1(new_n588_), .B2(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n607_), .A2(new_n634_), .A3(new_n635_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(G1327gat));
  INV_X1    g439(.A(new_n248_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n558_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n597_), .A2(new_n642_), .A3(new_n532_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(KEYINPUT107), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT107), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n586_), .A2(new_n645_), .A3(new_n532_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n644_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT44), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(KEYINPUT109), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT43), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n415_), .A2(new_n651_), .A3(new_n604_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n651_), .B1(new_n415_), .B2(new_n604_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n650_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(KEYINPUT109), .B1(new_n648_), .B2(KEYINPUT108), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(KEYINPUT43), .B1(new_n596_), .B2(new_n605_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n415_), .A2(new_n651_), .A3(new_n604_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n655_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n659_), .A2(new_n650_), .A3(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n641_), .B1(new_n656_), .B2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(G29gat), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n491_), .A2(new_n531_), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n664_), .A2(new_n597_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n415_), .A2(new_n642_), .A3(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT110), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n415_), .A2(KEYINPUT110), .A3(new_n642_), .A4(new_n665_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n248_), .A2(new_n663_), .ZN(new_n671_));
  OAI22_X1  g470(.A1(new_n662_), .A2(new_n663_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT111), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  OAI221_X1 g473(.A(KEYINPUT111), .B1(new_n670_), .B2(new_n671_), .C1(new_n662_), .C2(new_n663_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(G1328gat));
  INV_X1    g475(.A(KEYINPUT46), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n368_), .A2(G36gat), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n668_), .A2(new_n669_), .A3(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(KEYINPUT112), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT112), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n668_), .A2(new_n681_), .A3(new_n669_), .A4(new_n678_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n680_), .A2(KEYINPUT45), .A3(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n368_), .B1(new_n656_), .B2(new_n661_), .ZN(new_n684_));
  INV_X1    g483(.A(G36gat), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n683_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(KEYINPUT45), .B1(new_n680_), .B2(new_n682_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n677_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n654_), .A2(new_n655_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n660_), .B1(new_n659_), .B2(new_n650_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n611_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(G36gat), .ZN(new_n692_));
  INV_X1    g491(.A(new_n687_), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n692_), .A2(KEYINPUT46), .A3(new_n693_), .A4(new_n683_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n688_), .A2(new_n694_), .ZN(G1329gat));
  INV_X1    g494(.A(KEYINPUT47), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n410_), .A2(new_n411_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n698_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(G43gat), .ZN(new_n700_));
  INV_X1    g499(.A(new_n670_), .ZN(new_n701_));
  INV_X1    g500(.A(G43gat), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n701_), .A2(new_n702_), .A3(new_n414_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n696_), .B1(new_n700_), .B2(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n697_), .B1(new_n656_), .B2(new_n661_), .ZN(new_n705_));
  OAI211_X1 g504(.A(new_n696_), .B(new_n703_), .C1(new_n705_), .C2(new_n702_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n704_), .A2(new_n707_), .ZN(G1330gat));
  AOI21_X1  g507(.A(G50gat), .B1(new_n701_), .B2(new_n635_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n656_), .A2(new_n661_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n635_), .A2(G50gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n709_), .B1(new_n710_), .B2(new_n711_), .ZN(G1331gat));
  NOR2_X1   g511(.A1(new_n596_), .A2(new_n642_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n606_), .A2(new_n597_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT113), .ZN(new_n716_));
  AOI211_X1 g515(.A(G57gat), .B(new_n641_), .C1(new_n715_), .C2(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n717_), .B1(new_n716_), .B2(new_n715_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n598_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n558_), .A2(new_n531_), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n492_), .A2(new_n719_), .A3(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(new_n248_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(G57gat), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n718_), .A2(new_n723_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT114), .ZN(G1332gat));
  INV_X1    g524(.A(G64gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n726_), .B1(new_n721_), .B2(new_n611_), .ZN(new_n727_));
  XOR2_X1   g526(.A(new_n727_), .B(KEYINPUT48), .Z(new_n728_));
  INV_X1    g527(.A(new_n715_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n729_), .A2(new_n726_), .A3(new_n611_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(G1333gat));
  INV_X1    g530(.A(G71gat), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n732_), .B1(new_n721_), .B2(new_n414_), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n733_), .B(KEYINPUT49), .Z(new_n734_));
  NAND3_X1  g533(.A1(new_n729_), .A2(new_n732_), .A3(new_n414_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(G1334gat));
  INV_X1    g535(.A(G78gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n737_), .B1(new_n721_), .B2(new_n635_), .ZN(new_n738_));
  XOR2_X1   g537(.A(new_n738_), .B(KEYINPUT50), .Z(new_n739_));
  NAND3_X1  g538(.A1(new_n729_), .A2(new_n737_), .A3(new_n635_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(G1335gat));
  AND2_X1   g540(.A1(new_n598_), .A2(new_n664_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n713_), .A2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(G85gat), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n744_), .A2(new_n745_), .A3(new_n248_), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n597_), .A2(new_n642_), .A3(new_n531_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n659_), .A2(new_n747_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n748_), .A2(new_n248_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n746_), .B1(new_n749_), .B2(new_n745_), .ZN(G1336gat));
  AOI21_X1  g549(.A(G92gat), .B1(new_n744_), .B2(new_n611_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n611_), .A2(G92gat), .ZN(new_n752_));
  XOR2_X1   g551(.A(new_n752_), .B(KEYINPUT115), .Z(new_n753_));
  AOI21_X1  g552(.A(new_n751_), .B1(new_n748_), .B2(new_n753_), .ZN(G1337gat));
  NAND2_X1  g553(.A1(new_n748_), .A2(new_n414_), .ZN(new_n755_));
  AND3_X1   g554(.A1(new_n698_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n756_));
  AOI22_X1  g555(.A1(new_n755_), .A2(G99gat), .B1(new_n744_), .B2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT51), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n757_), .B(new_n758_), .ZN(G1338gat));
  NAND3_X1  g558(.A1(new_n659_), .A2(new_n635_), .A3(new_n747_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(G106gat), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT52), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n760_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n713_), .A2(new_n742_), .A3(new_n429_), .A4(new_n635_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT116), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n765_), .B(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n763_), .A2(new_n764_), .A3(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(KEYINPUT53), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT53), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n763_), .A2(new_n770_), .A3(new_n764_), .A4(new_n767_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n769_), .A2(new_n771_), .ZN(G1339gat));
  INV_X1    g571(.A(new_n597_), .ZN(new_n773_));
  NOR4_X1   g572(.A1(new_n773_), .A2(new_n604_), .A3(KEYINPUT54), .A4(new_n720_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT54), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n604_), .A2(new_n720_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n776_), .B2(new_n597_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n774_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT120), .ZN(new_n779_));
  INV_X1    g578(.A(new_n577_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n557_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n556_), .B1(new_n555_), .B2(new_n551_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n780_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT56), .ZN(new_n784_));
  AOI22_X1  g583(.A1(new_n562_), .A2(new_n563_), .B1(new_n455_), .B2(new_n508_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n565_), .B1(new_n785_), .B2(new_n566_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n568_), .A2(KEYINPUT117), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n787_), .B2(KEYINPUT55), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT55), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n568_), .A2(KEYINPUT117), .A3(new_n789_), .ZN(new_n790_));
  AOI211_X1 g589(.A(new_n784_), .B(new_n579_), .C1(new_n788_), .C2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n787_), .A2(KEYINPUT55), .ZN(new_n792_));
  INV_X1    g591(.A(new_n786_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n792_), .A2(new_n790_), .A3(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n579_), .ZN(new_n795_));
  AOI21_X1  g594(.A(KEYINPUT56), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n783_), .B1(new_n791_), .B2(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n535_), .B1(new_n549_), .B2(new_n536_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n536_), .B1(new_n501_), .B2(new_n541_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n799_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n798_), .A2(new_n800_), .A3(KEYINPUT118), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(new_n553_), .ZN(new_n802_));
  AOI21_X1  g601(.A(KEYINPUT118), .B1(new_n798_), .B2(new_n800_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n580_), .A2(KEYINPUT119), .A3(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT119), .B1(new_n580_), .B2(new_n804_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n490_), .B1(new_n797_), .B2(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n779_), .B1(new_n809_), .B2(KEYINPUT57), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n577_), .B1(new_n554_), .B2(new_n557_), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n568_), .A2(KEYINPUT117), .A3(new_n789_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n789_), .B1(new_n568_), .B2(KEYINPUT117), .ZN(new_n813_));
  NOR3_X1   g612(.A1(new_n812_), .A2(new_n813_), .A3(new_n786_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n784_), .B1(new_n814_), .B2(new_n579_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n794_), .A2(KEYINPUT56), .A3(new_n795_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n811_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n580_), .A2(new_n804_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT119), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n805_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n491_), .B1(new_n817_), .B2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT57), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n822_), .A2(KEYINPUT120), .A3(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n809_), .A2(KEYINPUT57), .ZN(new_n825_));
  NOR3_X1   g624(.A1(new_n780_), .A2(new_n802_), .A3(new_n803_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(new_n791_), .B2(new_n796_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT58), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  OAI211_X1 g628(.A(KEYINPUT58), .B(new_n826_), .C1(new_n791_), .C2(new_n796_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n829_), .A2(new_n830_), .A3(new_n604_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n810_), .A2(new_n824_), .A3(new_n825_), .A4(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n778_), .B1(new_n832_), .B2(new_n532_), .ZN(new_n833_));
  NOR4_X1   g632(.A1(new_n611_), .A2(new_n697_), .A3(new_n641_), .A4(new_n635_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n833_), .A2(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(G113gat), .B1(new_n836_), .B2(new_n642_), .ZN(new_n837_));
  OAI21_X1  g636(.A(KEYINPUT59), .B1(new_n833_), .B2(new_n835_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT121), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n835_), .A2(KEYINPUT59), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n822_), .A2(new_n823_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n841_), .A2(new_n825_), .A3(new_n831_), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n842_), .A2(new_n532_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n840_), .B1(new_n843_), .B2(new_n778_), .ZN(new_n844_));
  AND3_X1   g643(.A1(new_n838_), .A2(new_n839_), .A3(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n839_), .B1(new_n838_), .B2(new_n844_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n642_), .A2(G113gat), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n837_), .B1(new_n847_), .B2(new_n848_), .ZN(G1340gat));
  AND3_X1   g648(.A1(new_n838_), .A2(new_n598_), .A3(new_n844_), .ZN(new_n850_));
  INV_X1    g649(.A(G120gat), .ZN(new_n851_));
  INV_X1    g650(.A(new_n836_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n851_), .B1(new_n597_), .B2(KEYINPUT60), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n851_), .A2(KEYINPUT60), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n853_), .B1(KEYINPUT122), .B2(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n855_), .B1(KEYINPUT122), .B2(new_n853_), .ZN(new_n856_));
  OAI22_X1  g655(.A1(new_n850_), .A2(new_n851_), .B1(new_n852_), .B2(new_n856_), .ZN(G1341gat));
  AOI21_X1  g656(.A(G127gat), .B1(new_n836_), .B2(new_n531_), .ZN(new_n858_));
  AND2_X1   g657(.A1(new_n531_), .A2(G127gat), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n858_), .B1(new_n847_), .B2(new_n859_), .ZN(G1342gat));
  AOI21_X1  g659(.A(G134gat), .B1(new_n836_), .B2(new_n490_), .ZN(new_n861_));
  AND2_X1   g660(.A1(new_n604_), .A2(G134gat), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n861_), .B1(new_n847_), .B2(new_n862_), .ZN(G1343gat));
  INV_X1    g662(.A(new_n833_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n611_), .A2(new_n641_), .A3(new_n384_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n864_), .A2(new_n595_), .A3(new_n865_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n866_), .A2(new_n558_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(new_n203_), .ZN(G1344gat));
  NOR2_X1   g667(.A1(new_n866_), .A2(new_n719_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(new_n204_), .ZN(G1345gat));
  NOR2_X1   g669(.A1(new_n866_), .A2(new_n532_), .ZN(new_n871_));
  XOR2_X1   g670(.A(KEYINPUT61), .B(G155gat), .Z(new_n872_));
  XNOR2_X1  g671(.A(new_n871_), .B(new_n872_), .ZN(G1346gat));
  OAI21_X1  g672(.A(G162gat), .B1(new_n866_), .B2(new_n605_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n490_), .A2(new_n218_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n866_), .B2(new_n875_), .ZN(G1347gat));
  INV_X1    g675(.A(KEYINPUT124), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n595_), .A2(new_n248_), .A3(new_n368_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n384_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  OAI211_X1 g679(.A(new_n877_), .B(new_n880_), .C1(new_n843_), .C2(new_n778_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n778_), .B1(new_n842_), .B2(new_n532_), .ZN(new_n882_));
  OAI21_X1  g681(.A(KEYINPUT124), .B1(new_n882_), .B2(new_n879_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n881_), .A2(new_n883_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n884_), .A2(new_n271_), .A3(new_n642_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n882_), .A2(new_n558_), .A3(new_n879_), .ZN(new_n886_));
  INV_X1    g685(.A(G169gat), .ZN(new_n887_));
  OAI21_X1  g686(.A(KEYINPUT123), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n642_), .B(new_n880_), .C1(new_n843_), .C2(new_n778_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT123), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n889_), .A2(new_n890_), .A3(G169gat), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT62), .ZN(new_n892_));
  AND3_X1   g691(.A1(new_n888_), .A2(new_n891_), .A3(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n892_), .B1(new_n888_), .B2(new_n891_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n885_), .B1(new_n893_), .B2(new_n894_), .ZN(G1348gat));
  NAND3_X1  g694(.A1(new_n878_), .A2(G176gat), .A3(new_n598_), .ZN(new_n896_));
  NOR3_X1   g695(.A1(new_n833_), .A2(new_n635_), .A3(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n884_), .A2(new_n773_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n898_), .A2(KEYINPUT125), .A3(new_n272_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT125), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n597_), .B1(new_n881_), .B2(new_n883_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(G176gat), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n897_), .B1(new_n899_), .B2(new_n902_), .ZN(G1349gat));
  NOR2_X1   g702(.A1(new_n532_), .A2(new_n260_), .ZN(new_n904_));
  NAND4_X1  g703(.A1(new_n864_), .A2(new_n384_), .A3(new_n531_), .A4(new_n878_), .ZN(new_n905_));
  INV_X1    g704(.A(G183gat), .ZN(new_n906_));
  AOI22_X1  g705(.A1(new_n884_), .A2(new_n904_), .B1(new_n905_), .B2(new_n906_), .ZN(G1350gat));
  NAND3_X1  g706(.A1(new_n884_), .A2(new_n490_), .A3(new_n319_), .ZN(new_n908_));
  INV_X1    g707(.A(G190gat), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n605_), .B1(new_n881_), .B2(new_n883_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n908_), .B1(new_n909_), .B2(new_n910_), .ZN(G1351gat));
  NAND3_X1  g710(.A1(new_n595_), .A2(new_n407_), .A3(new_n611_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n833_), .A2(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(KEYINPUT126), .A2(G197gat), .ZN(new_n914_));
  OR2_X1    g713(.A1(KEYINPUT126), .A2(G197gat), .ZN(new_n915_));
  AOI22_X1  g714(.A1(new_n913_), .A2(new_n642_), .B1(new_n914_), .B2(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n913_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n917_), .A2(new_n558_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n916_), .B1(new_n918_), .B2(new_n915_), .ZN(G1352gat));
  NAND2_X1  g718(.A1(new_n913_), .A2(new_n598_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g720(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n913_), .A2(new_n531_), .A3(new_n922_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n924_));
  XOR2_X1   g723(.A(new_n923_), .B(new_n924_), .Z(G1354gat));
  OR3_X1    g724(.A1(new_n917_), .A2(G218gat), .A3(new_n491_), .ZN(new_n926_));
  OAI21_X1  g725(.A(G218gat), .B1(new_n917_), .B2(new_n605_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n926_), .A2(new_n927_), .ZN(G1355gat));
endmodule


