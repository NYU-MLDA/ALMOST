//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 1 1 0 0 1 1 1 1 1 0 1 1 0 0 1 1 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 0 0 1 0 1 0 1 1 0 0 0 1 0 0 0 0 1 1 0 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n713_, new_n714_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n766_,
    new_n767_, new_n768_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n890_, new_n891_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n916_, new_n917_,
    new_n919_, new_n920_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n928_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n936_, new_n937_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT23), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT23), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n204_), .A2(G183gat), .A3(G190gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n205_), .A3(KEYINPUT81), .ZN(new_n206_));
  OR3_X1    g005(.A1(new_n202_), .A2(KEYINPUT81), .A3(KEYINPUT23), .ZN(new_n207_));
  INV_X1    g006(.A(G183gat), .ZN(new_n208_));
  INV_X1    g007(.A(G190gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n206_), .A2(new_n207_), .A3(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(KEYINPUT80), .A2(G169gat), .ZN(new_n212_));
  AOI21_X1  g011(.A(G176gat), .B1(new_n212_), .B2(KEYINPUT22), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT22), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(KEYINPUT80), .A3(G169gat), .ZN(new_n215_));
  AOI22_X1  g014(.A1(new_n213_), .A2(new_n215_), .B1(G169gat), .B2(G176gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n211_), .A2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT26), .B(G190gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT25), .B1(new_n208_), .B2(KEYINPUT79), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT25), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(G183gat), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n218_), .B(new_n219_), .C1(KEYINPUT79), .C2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(G169gat), .ZN(new_n223_));
  INV_X1    g022(.A(G176gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(KEYINPUT24), .A3(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT24), .ZN(new_n228_));
  NOR2_X1   g027(.A1(G169gat), .A2(G176gat), .ZN(new_n229_));
  AOI22_X1  g028(.A1(new_n203_), .A2(new_n205_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n222_), .A2(new_n227_), .A3(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n217_), .A2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G197gat), .B(G204gat), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT21), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(G218gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(G211gat), .ZN(new_n237_));
  INV_X1    g036(.A(G211gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(G218gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(G204gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(G197gat), .ZN(new_n243_));
  INV_X1    g042(.A(G197gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(G204gat), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT88), .ZN(new_n246_));
  AND3_X1   g045(.A1(new_n243_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n242_), .A2(KEYINPUT88), .A3(G197gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT21), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n235_), .B(new_n241_), .C1(new_n247_), .C2(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n233_), .A2(new_n234_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(new_n240_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT20), .B1(new_n232_), .B2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n203_), .A2(new_n205_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(new_n210_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT22), .B(G169gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(new_n224_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n256_), .A2(new_n226_), .A3(new_n258_), .ZN(new_n259_));
  AND2_X1   g058(.A1(KEYINPUT91), .A2(KEYINPUT24), .ZN(new_n260_));
  NOR2_X1   g059(.A1(KEYINPUT91), .A2(KEYINPUT24), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n229_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n225_), .A2(new_n226_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT91), .B(KEYINPUT24), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n262_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n208_), .A2(KEYINPUT25), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n220_), .A2(G183gat), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT90), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n208_), .A2(KEYINPUT25), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT90), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n221_), .A2(new_n269_), .A3(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n268_), .A2(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n265_), .B1(new_n272_), .B2(new_n218_), .ZN(new_n273_));
  AND2_X1   g072(.A1(new_n206_), .A2(new_n207_), .ZN(new_n274_));
  AOI21_X1  g073(.A(KEYINPUT92), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  AND3_X1   g074(.A1(new_n221_), .A2(new_n269_), .A3(new_n270_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n270_), .B1(new_n221_), .B2(new_n269_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n218_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  OR2_X1    g077(.A1(KEYINPUT91), .A2(KEYINPUT24), .ZN(new_n279_));
  NAND2_X1  g078(.A1(KEYINPUT91), .A2(KEYINPUT24), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n279_), .A2(new_n225_), .A3(new_n226_), .A4(new_n280_), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n281_), .A2(new_n262_), .ZN(new_n282_));
  AND4_X1   g081(.A1(KEYINPUT92), .A2(new_n278_), .A3(new_n282_), .A4(new_n274_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n259_), .B1(new_n275_), .B2(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n254_), .B1(new_n284_), .B2(new_n253_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G226gat), .A2(G233gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT19), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT89), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT20), .ZN(new_n290_));
  AND3_X1   g089(.A1(new_n250_), .A2(new_n259_), .A3(new_n252_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n278_), .A2(new_n282_), .A3(new_n274_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n290_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n229_), .A2(new_n228_), .ZN(new_n294_));
  AND3_X1   g093(.A1(new_n255_), .A2(new_n227_), .A3(new_n294_), .ZN(new_n295_));
  AOI22_X1  g094(.A1(new_n295_), .A2(new_n222_), .B1(new_n211_), .B2(new_n216_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n240_), .B1(new_n234_), .B2(new_n233_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n243_), .A2(new_n245_), .ZN(new_n298_));
  OAI211_X1 g097(.A(KEYINPUT21), .B(new_n248_), .C1(new_n298_), .C2(KEYINPUT88), .ZN(new_n299_));
  AOI22_X1  g098(.A1(new_n297_), .A2(new_n299_), .B1(new_n240_), .B2(new_n251_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT93), .ZN(new_n301_));
  NOR3_X1   g100(.A1(new_n296_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(KEYINPUT93), .B1(new_n232_), .B2(new_n253_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n293_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  AOI22_X1  g103(.A1(new_n285_), .A2(new_n289_), .B1(new_n287_), .B2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G8gat), .B(G36gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT18), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G64gat), .B(G92gat), .ZN(new_n308_));
  XOR2_X1   g107(.A(new_n307_), .B(new_n308_), .Z(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT27), .B1(new_n305_), .B2(new_n309_), .ZN(new_n310_));
  OAI211_X1 g109(.A(new_n300_), .B(new_n259_), .C1(new_n275_), .C2(new_n283_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n301_), .B1(new_n296_), .B2(new_n300_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n232_), .A2(KEYINPUT93), .A3(new_n253_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n287_), .A2(new_n290_), .ZN(new_n315_));
  AND3_X1   g114(.A1(new_n311_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT94), .ZN(new_n317_));
  INV_X1    g116(.A(new_n254_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n259_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT92), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n292_), .A2(new_n320_), .ZN(new_n321_));
  NAND4_X1  g120(.A1(new_n278_), .A2(new_n282_), .A3(new_n274_), .A4(KEYINPUT92), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n319_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n318_), .B1(new_n323_), .B2(new_n300_), .ZN(new_n324_));
  AOI22_X1  g123(.A1(new_n316_), .A2(new_n317_), .B1(new_n324_), .B2(new_n288_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n311_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(KEYINPUT94), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n325_), .A2(KEYINPUT100), .A3(new_n327_), .A4(new_n309_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n324_), .A2(new_n288_), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n311_), .A2(new_n314_), .A3(new_n317_), .A4(new_n315_), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n327_), .A2(new_n329_), .A3(new_n330_), .A4(new_n309_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT100), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n310_), .B1(new_n328_), .B2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT101), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n327_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n309_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(KEYINPUT27), .B1(new_n338_), .B2(new_n331_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n335_), .A2(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(G155gat), .A2(G162gat), .ZN(new_n342_));
  AND2_X1   g141(.A1(G155gat), .A2(G162gat), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT1), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n342_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT84), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n346_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G155gat), .A2(G162gat), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n348_), .A2(KEYINPUT84), .A3(KEYINPUT1), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n345_), .A2(new_n347_), .A3(new_n349_), .ZN(new_n350_));
  XOR2_X1   g149(.A(G141gat), .B(G148gat), .Z(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT3), .ZN(new_n353_));
  INV_X1    g152(.A(G141gat), .ZN(new_n354_));
  INV_X1    g153(.A(G148gat), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n353_), .A2(new_n354_), .A3(new_n355_), .A4(KEYINPUT85), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT85), .ZN(new_n357_));
  OAI22_X1  g156(.A1(new_n357_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G141gat), .A2(G148gat), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT2), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n356_), .A2(new_n358_), .A3(new_n361_), .A4(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT86), .ZN(new_n364_));
  OR3_X1    g163(.A1(new_n343_), .A2(new_n342_), .A3(new_n364_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n364_), .B1(new_n343_), .B2(new_n342_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n363_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n352_), .A2(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n368_), .A2(KEYINPUT29), .ZN(new_n369_));
  XOR2_X1   g168(.A(G22gat), .B(G50gat), .Z(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G228gat), .A2(G233gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(G78gat), .ZN(new_n373_));
  INV_X1    g172(.A(G106gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  AND2_X1   g174(.A1(new_n371_), .A2(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n371_), .A2(new_n375_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n300_), .B1(new_n368_), .B2(KEYINPUT29), .ZN(new_n378_));
  XNOR2_X1  g177(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n379_));
  XOR2_X1   g178(.A(new_n378_), .B(new_n379_), .Z(new_n380_));
  OR3_X1    g179(.A1(new_n376_), .A2(new_n377_), .A3(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n380_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G1gat), .B(G29gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(G85gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT0), .B(G57gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n386_), .B(new_n387_), .ZN(new_n388_));
  XOR2_X1   g187(.A(G127gat), .B(G134gat), .Z(new_n389_));
  INV_X1    g188(.A(G120gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(G113gat), .ZN(new_n391_));
  INV_X1    g190(.A(G113gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(G120gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n391_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n389_), .A2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G127gat), .B(G134gat), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n396_), .A2(new_n391_), .A3(new_n393_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n395_), .A2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n352_), .A2(new_n367_), .A3(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n398_), .B1(new_n352_), .B2(new_n367_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G225gat), .A2(G233gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n403_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n398_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n368_), .A2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n407_), .A2(KEYINPUT4), .A3(new_n399_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT95), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT4), .ZN(new_n410_));
  AND4_X1   g209(.A1(new_n409_), .A2(new_n368_), .A3(new_n410_), .A4(new_n406_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n409_), .B1(new_n401_), .B2(new_n410_), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n405_), .B(new_n408_), .C1(new_n411_), .C2(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n404_), .B1(new_n413_), .B2(KEYINPUT96), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT96), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n403_), .B1(new_n402_), .B2(KEYINPUT4), .ZN(new_n416_));
  OAI21_X1  g215(.A(KEYINPUT95), .B1(new_n407_), .B2(KEYINPUT4), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n401_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n415_), .B1(new_n416_), .B2(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n388_), .B1(new_n414_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT99), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n413_), .A2(KEYINPUT96), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n416_), .A2(new_n415_), .A3(new_n419_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n388_), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n423_), .A2(new_n424_), .A3(new_n425_), .A4(new_n404_), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n421_), .A2(new_n422_), .A3(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n422_), .B1(new_n421_), .B2(new_n426_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(G227gat), .A2(G233gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n431_), .B(KEYINPUT83), .ZN(new_n432_));
  XOR2_X1   g231(.A(G71gat), .B(G99gat), .Z(new_n433_));
  XNOR2_X1  g232(.A(new_n432_), .B(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n296_), .B(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(new_n398_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G15gat), .B(G43gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(KEYINPUT82), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(KEYINPUT30), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(KEYINPUT31), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n436_), .A2(new_n440_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n436_), .A2(new_n440_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n430_), .A2(new_n443_), .ZN(new_n444_));
  OR3_X1    g243(.A1(new_n341_), .A2(new_n384_), .A3(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n421_), .A2(new_n426_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n309_), .A2(KEYINPUT32), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n325_), .A2(new_n327_), .A3(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n304_), .A2(new_n287_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n449_), .B1(new_n324_), .B2(new_n288_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n450_), .A2(KEYINPUT32), .A3(new_n309_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n446_), .A2(new_n448_), .A3(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT98), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n446_), .A2(KEYINPUT98), .A3(new_n448_), .A4(new_n451_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n419_), .A2(new_n403_), .A3(new_n408_), .ZN(new_n456_));
  OR3_X1    g255(.A1(new_n400_), .A2(new_n401_), .A3(KEYINPUT97), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT97), .B1(new_n400_), .B2(new_n401_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n457_), .A2(new_n405_), .A3(new_n458_), .ZN(new_n459_));
  AND3_X1   g258(.A1(new_n456_), .A2(new_n388_), .A3(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT33), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n460_), .B1(new_n426_), .B2(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n414_), .A2(new_n420_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n463_), .A2(KEYINPUT33), .A3(new_n425_), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n462_), .A2(new_n464_), .A3(new_n331_), .A4(new_n338_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n454_), .A2(new_n455_), .A3(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(new_n383_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n446_), .A2(KEYINPUT99), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n421_), .A2(new_n426_), .A3(new_n422_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n383_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n328_), .A2(new_n333_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n310_), .ZN(new_n472_));
  AOI21_X1  g271(.A(KEYINPUT101), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT101), .ZN(new_n474_));
  AOI211_X1 g273(.A(new_n474_), .B(new_n310_), .C1(new_n328_), .C2(new_n333_), .ZN(new_n475_));
  OAI211_X1 g274(.A(new_n340_), .B(new_n470_), .C1(new_n473_), .C2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n467_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n443_), .ZN(new_n478_));
  AOI21_X1  g277(.A(KEYINPUT102), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT102), .ZN(new_n480_));
  AOI211_X1 g279(.A(new_n480_), .B(new_n443_), .C1(new_n467_), .C2(new_n476_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n445_), .B1(new_n479_), .B2(new_n481_), .ZN(new_n482_));
  XOR2_X1   g281(.A(G15gat), .B(G22gat), .Z(new_n483_));
  NAND2_X1  g282(.A1(G1gat), .A2(G8gat), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n483_), .B1(KEYINPUT14), .B2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT74), .ZN(new_n486_));
  XOR2_X1   g285(.A(G1gat), .B(G8gat), .Z(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n486_), .B(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G29gat), .B(G36gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G43gat), .B(G50gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n489_), .A2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n486_), .B(new_n487_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n492_), .B(KEYINPUT15), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G229gat), .A2(G233gat), .ZN(new_n497_));
  AND3_X1   g296(.A1(new_n493_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT77), .ZN(new_n499_));
  INV_X1    g298(.A(new_n492_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n494_), .A2(new_n500_), .ZN(new_n501_));
  OR2_X1    g300(.A1(new_n486_), .A2(new_n487_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n486_), .A2(new_n487_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n492_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n499_), .B1(new_n501_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n497_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n494_), .A2(new_n500_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n493_), .A2(new_n507_), .A3(KEYINPUT77), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n505_), .A2(new_n506_), .A3(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT78), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT78), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n505_), .A2(new_n511_), .A3(new_n508_), .A4(new_n506_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n498_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n513_));
  XOR2_X1   g312(.A(G113gat), .B(G141gat), .Z(new_n514_));
  XNOR2_X1  g313(.A(G169gat), .B(G197gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  AND2_X1   g315(.A1(new_n513_), .A2(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n513_), .A2(new_n516_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G230gat), .A2(G233gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT64), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G85gat), .B(G92gat), .ZN(new_n523_));
  OR2_X1    g322(.A1(new_n523_), .A2(KEYINPUT66), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(KEYINPUT66), .ZN(new_n525_));
  NOR2_X1   g324(.A1(G99gat), .A2(G106gat), .ZN(new_n526_));
  XOR2_X1   g325(.A(new_n526_), .B(KEYINPUT7), .Z(new_n527_));
  NAND2_X1  g326(.A1(G99gat), .A2(G106gat), .ZN(new_n528_));
  XOR2_X1   g327(.A(new_n528_), .B(KEYINPUT6), .Z(new_n529_));
  OAI211_X1 g328(.A(new_n524_), .B(new_n525_), .C1(new_n527_), .C2(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT8), .ZN(new_n531_));
  INV_X1    g330(.A(G92gat), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n523_), .B1(KEYINPUT9), .B2(new_n532_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n533_), .B1(KEYINPUT9), .B2(new_n523_), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n534_), .A2(KEYINPUT65), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(KEYINPUT65), .ZN(new_n536_));
  XOR2_X1   g335(.A(KEYINPUT10), .B(G99gat), .Z(new_n537_));
  AOI21_X1  g336(.A(new_n529_), .B1(new_n374_), .B2(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n535_), .A2(new_n536_), .A3(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n531_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT67), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G57gat), .B(G64gat), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT11), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT68), .ZN(new_n545_));
  XOR2_X1   g344(.A(G71gat), .B(G78gat), .Z(new_n546_));
  OAI21_X1  g345(.A(new_n546_), .B1(KEYINPUT11), .B2(new_n543_), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n545_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n545_), .A2(new_n547_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n542_), .A2(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n540_), .B(KEYINPUT67), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(new_n550_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n522_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT69), .ZN(new_n556_));
  OR2_X1    g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n540_), .A2(new_n551_), .A3(KEYINPUT12), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n554_), .A2(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(KEYINPUT12), .B1(new_n542_), .B2(new_n551_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(new_n522_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n555_), .A2(new_n556_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n557_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(G120gat), .B(G148gat), .Z(new_n565_));
  XNOR2_X1  g364(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  XOR2_X1   g366(.A(G176gat), .B(G204gat), .Z(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT71), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n564_), .A2(new_n571_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n557_), .A2(new_n562_), .A3(new_n569_), .A4(new_n563_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(KEYINPUT13), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT13), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n572_), .A2(new_n576_), .A3(new_n573_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n575_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n553_), .A2(new_n492_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n540_), .A2(new_n495_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(KEYINPUT72), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G232gat), .A2(G233gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT34), .ZN(new_n584_));
  AND3_X1   g383(.A1(new_n582_), .A2(KEYINPUT35), .A3(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n581_), .A2(new_n586_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n584_), .A2(KEYINPUT35), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n579_), .B(new_n580_), .C1(new_n585_), .C2(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(G134gat), .B(G162gat), .Z(new_n590_));
  XNOR2_X1  g389(.A(G190gat), .B(G218gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT36), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n587_), .A2(new_n589_), .A3(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n595_), .A2(new_n593_), .A3(new_n592_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n592_), .A2(new_n593_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n587_), .A2(new_n589_), .A3(new_n597_), .A4(new_n594_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(KEYINPUT73), .B(KEYINPUT37), .ZN(new_n599_));
  AND3_X1   g398(.A1(new_n596_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(KEYINPUT73), .A2(KEYINPUT37), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n601_), .B1(new_n596_), .B2(new_n598_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G231gat), .A2(G233gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n550_), .B(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(new_n489_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G127gat), .B(G155gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G183gat), .B(G211gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT17), .Z(new_n612_));
  OR2_X1    g411(.A1(new_n606_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(KEYINPUT17), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n606_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n613_), .A2(new_n615_), .ZN(new_n616_));
  OR2_X1    g415(.A1(new_n616_), .A2(KEYINPUT76), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(KEYINPUT76), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n603_), .A2(new_n620_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n482_), .A2(new_n520_), .A3(new_n578_), .A4(new_n621_), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n622_), .B(KEYINPUT103), .Z(new_n623_));
  INV_X1    g422(.A(G1gat), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n429_), .A2(KEYINPUT104), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n429_), .A2(KEYINPUT104), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n623_), .A2(new_n624_), .A3(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT38), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n578_), .A2(new_n520_), .A3(new_n619_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT105), .ZN(new_n633_));
  NOR3_X1   g432(.A1(new_n341_), .A2(new_n384_), .A3(new_n444_), .ZN(new_n634_));
  NOR3_X1   g433(.A1(new_n429_), .A2(new_n383_), .A3(new_n339_), .ZN(new_n635_));
  AOI22_X1  g434(.A1(new_n335_), .A2(new_n635_), .B1(new_n466_), .B2(new_n383_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n480_), .B1(new_n636_), .B2(new_n443_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n477_), .A2(KEYINPUT102), .A3(new_n478_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n634_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n596_), .A2(new_n598_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n633_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n640_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n482_), .A2(KEYINPUT105), .A3(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n632_), .B1(new_n641_), .B2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(G1gat), .B1(new_n645_), .B2(new_n430_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n629_), .A2(new_n630_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n631_), .A2(new_n646_), .A3(new_n647_), .ZN(G1324gat));
  INV_X1    g447(.A(G8gat), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n623_), .A2(new_n649_), .A3(new_n341_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT39), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n644_), .A2(new_n341_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n651_), .B1(new_n652_), .B2(G8gat), .ZN(new_n653_));
  AOI211_X1 g452(.A(KEYINPUT39), .B(new_n649_), .C1(new_n644_), .C2(new_n341_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n650_), .B1(new_n653_), .B2(new_n654_), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n655_), .B(KEYINPUT40), .Z(G1325gat));
  OR3_X1    g455(.A1(new_n622_), .A2(G15gat), .A3(new_n478_), .ZN(new_n657_));
  OAI21_X1  g456(.A(G15gat), .B1(new_n645_), .B2(new_n478_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT41), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n658_), .A2(new_n659_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n657_), .B1(new_n660_), .B2(new_n661_), .ZN(G1326gat));
  OR3_X1    g461(.A1(new_n622_), .A2(G22gat), .A3(new_n383_), .ZN(new_n663_));
  OAI21_X1  g462(.A(G22gat), .B1(new_n645_), .B2(new_n383_), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n664_), .A2(KEYINPUT42), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n664_), .A2(KEYINPUT42), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n663_), .B1(new_n665_), .B2(new_n666_), .ZN(G1327gat));
  INV_X1    g466(.A(new_n578_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n642_), .A2(new_n619_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  NOR4_X1   g469(.A1(new_n639_), .A2(new_n668_), .A3(new_n670_), .A4(new_n519_), .ZN(new_n671_));
  INV_X1    g470(.A(G29gat), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n671_), .A2(new_n672_), .A3(new_n429_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT43), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n674_), .B1(new_n603_), .B2(KEYINPUT106), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n596_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n676_), .B1(new_n640_), .B2(new_n601_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n675_), .B1(new_n639_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT106), .ZN(new_n679_));
  OAI21_X1  g478(.A(KEYINPUT43), .B1(new_n677_), .B2(new_n679_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n482_), .A2(new_n603_), .A3(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n678_), .A2(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n578_), .A2(new_n520_), .A3(new_n620_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(KEYINPUT44), .B1(new_n682_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n686_));
  AOI211_X1 g485(.A(new_n686_), .B(new_n683_), .C1(new_n678_), .C2(new_n681_), .ZN(new_n687_));
  NOR3_X1   g486(.A1(new_n685_), .A2(new_n687_), .A3(new_n627_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n673_), .B1(new_n688_), .B2(new_n672_), .ZN(G1328gat));
  INV_X1    g488(.A(G36gat), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n671_), .A2(new_n690_), .A3(new_n341_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT45), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n685_), .A2(new_n687_), .ZN(new_n693_));
  AOI21_X1  g492(.A(KEYINPUT107), .B1(new_n693_), .B2(new_n341_), .ZN(new_n694_));
  NOR3_X1   g493(.A1(new_n639_), .A2(new_n675_), .A3(new_n677_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n680_), .B1(new_n482_), .B2(new_n603_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n684_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(new_n686_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n682_), .A2(KEYINPUT44), .A3(new_n684_), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n698_), .A2(KEYINPUT107), .A3(new_n341_), .A4(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(G36gat), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n692_), .B1(new_n694_), .B2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT108), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n703_), .A2(KEYINPUT46), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n704_), .ZN(new_n705_));
  OAI221_X1 g504(.A(new_n692_), .B1(new_n703_), .B2(KEYINPUT46), .C1(new_n694_), .C2(new_n701_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(G1329gat));
  NAND3_X1  g506(.A1(new_n693_), .A2(G43gat), .A3(new_n443_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n671_), .A2(new_n443_), .ZN(new_n709_));
  OR2_X1    g508(.A1(new_n709_), .A2(G43gat), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(new_n710_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g511(.A(G50gat), .B1(new_n671_), .B2(new_n384_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n384_), .A2(G50gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n693_), .B2(new_n714_), .ZN(G1331gat));
  NAND3_X1  g514(.A1(new_n668_), .A2(new_n519_), .A3(new_n619_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n716_), .B1(new_n641_), .B2(new_n643_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(G57gat), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n718_), .A2(new_n719_), .A3(new_n430_), .ZN(new_n720_));
  AOI21_X1  g519(.A(KEYINPUT109), .B1(new_n482_), .B2(new_n519_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n721_), .A2(new_n578_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n482_), .A2(KEYINPUT109), .A3(new_n519_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  NOR3_X1   g523(.A1(new_n724_), .A2(new_n620_), .A3(new_n603_), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n725_), .A2(KEYINPUT110), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(KEYINPUT110), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n726_), .A2(new_n628_), .A3(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n720_), .B1(new_n728_), .B2(new_n719_), .ZN(G1332gat));
  INV_X1    g528(.A(new_n341_), .ZN(new_n730_));
  OAI21_X1  g529(.A(G64gat), .B1(new_n718_), .B2(new_n730_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n731_), .A2(KEYINPUT48), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n731_), .A2(KEYINPUT48), .ZN(new_n733_));
  INV_X1    g532(.A(new_n725_), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n730_), .A2(G64gat), .ZN(new_n735_));
  OAI22_X1  g534(.A1(new_n732_), .A2(new_n733_), .B1(new_n734_), .B2(new_n735_), .ZN(G1333gat));
  OR2_X1    g535(.A1(new_n478_), .A2(G71gat), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n717_), .A2(new_n443_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(KEYINPUT111), .B(KEYINPUT49), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n738_), .A2(G71gat), .A3(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n738_), .B2(G71gat), .ZN(new_n741_));
  OAI22_X1  g540(.A1(new_n734_), .A2(new_n737_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT112), .ZN(G1334gat));
  OAI21_X1  g542(.A(G78gat), .B1(new_n718_), .B2(new_n383_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n744_), .A2(KEYINPUT50), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n744_), .A2(KEYINPUT50), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n383_), .A2(G78gat), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT113), .ZN(new_n748_));
  OAI22_X1  g547(.A1(new_n745_), .A2(new_n746_), .B1(new_n734_), .B2(new_n748_), .ZN(G1335gat));
  NAND4_X1  g548(.A1(new_n575_), .A2(new_n519_), .A3(new_n577_), .A4(new_n620_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT114), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n682_), .A2(new_n751_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n752_), .A2(KEYINPUT115), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT115), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n754_), .B1(new_n682_), .B2(new_n751_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n753_), .A2(new_n755_), .ZN(new_n756_));
  OAI21_X1  g555(.A(G85gat), .B1(new_n756_), .B2(new_n430_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n722_), .A2(new_n669_), .A3(new_n723_), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n758_), .A2(G85gat), .A3(new_n627_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n757_), .A2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT116), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n757_), .A2(KEYINPUT116), .A3(new_n760_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(G1336gat));
  OAI21_X1  g564(.A(G92gat), .B1(new_n756_), .B2(new_n730_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n758_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n767_), .A2(new_n532_), .A3(new_n341_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(G1337gat));
  INV_X1    g568(.A(KEYINPUT117), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT51), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n443_), .A2(new_n537_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n771_), .B1(new_n758_), .B2(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n443_), .B1(new_n753_), .B2(new_n755_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n773_), .B1(new_n774_), .B2(G99gat), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n770_), .A2(KEYINPUT51), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n775_), .B(new_n776_), .ZN(G1338gat));
  NAND3_X1  g576(.A1(new_n767_), .A2(new_n374_), .A3(new_n384_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n752_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n384_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT52), .ZN(new_n781_));
  OAI21_X1  g580(.A(G106gat), .B1(new_n781_), .B2(KEYINPUT118), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  AOI22_X1  g582(.A1(new_n780_), .A2(new_n783_), .B1(KEYINPUT118), .B2(new_n781_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n781_), .A2(KEYINPUT118), .ZN(new_n785_));
  AOI211_X1 g584(.A(new_n785_), .B(new_n782_), .C1(new_n779_), .C2(new_n384_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n778_), .B1(new_n784_), .B2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(KEYINPUT53), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT53), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n778_), .B(new_n789_), .C1(new_n784_), .C2(new_n786_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n790_), .ZN(G1339gat));
  NAND3_X1  g590(.A1(new_n621_), .A2(new_n519_), .A3(new_n578_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n792_), .B(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT121), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n505_), .A2(new_n497_), .A3(new_n508_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n501_), .A2(new_n497_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n516_), .B1(new_n797_), .B2(new_n496_), .ZN(new_n798_));
  AOI22_X1  g597(.A1(new_n513_), .A2(new_n516_), .B1(new_n796_), .B2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n573_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT120), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT120), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n573_), .A2(new_n799_), .A3(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n553_), .A2(new_n550_), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n554_), .B(new_n558_), .C1(new_n805_), .C2(KEYINPUT12), .ZN(new_n806_));
  INV_X1    g605(.A(new_n522_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n804_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n561_), .A2(KEYINPUT55), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n522_), .A2(KEYINPUT119), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n808_), .A2(new_n809_), .A3(new_n811_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n806_), .A2(new_n804_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n570_), .B1(new_n813_), .B2(new_n810_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n812_), .A2(new_n814_), .A3(KEYINPUT56), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(KEYINPUT56), .B1(new_n812_), .B2(new_n814_), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n801_), .B(new_n803_), .C1(new_n816_), .C2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT58), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n812_), .A2(new_n814_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT56), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n815_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT58), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n823_), .A2(new_n824_), .A3(new_n801_), .A4(new_n803_), .ZN(new_n825_));
  AND2_X1   g624(.A1(new_n819_), .A2(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n795_), .B1(new_n826_), .B2(new_n677_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n573_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n828_), .B1(new_n822_), .B2(new_n815_), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n574_), .A2(new_n799_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n642_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT57), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  OAI211_X1 g632(.A(KEYINPUT57), .B(new_n642_), .C1(new_n829_), .C2(new_n830_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n677_), .B1(new_n819_), .B2(new_n825_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT121), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n827_), .A2(new_n835_), .A3(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n794_), .B1(new_n838_), .B2(new_n620_), .ZN(new_n839_));
  NOR4_X1   g638(.A1(new_n341_), .A2(new_n627_), .A3(new_n384_), .A4(new_n478_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(KEYINPUT122), .B1(new_n839_), .B2(new_n841_), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n833_), .B(new_n834_), .C1(new_n836_), .C2(KEYINPUT121), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n836_), .A2(KEYINPUT121), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n620_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n794_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT122), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n847_), .A2(new_n848_), .A3(new_n840_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n842_), .A2(new_n849_), .A3(new_n520_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n847_), .A2(new_n840_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n833_), .A2(new_n834_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n620_), .B1(new_n852_), .B2(new_n836_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n794_), .B1(new_n853_), .B2(KEYINPUT123), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT123), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n855_), .B(new_n620_), .C1(new_n852_), .C2(new_n836_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n854_), .A2(new_n856_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n841_), .A2(KEYINPUT59), .ZN(new_n858_));
  AOI22_X1  g657(.A1(new_n851_), .A2(KEYINPUT59), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n520_), .A2(G113gat), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(KEYINPUT124), .ZN(new_n861_));
  AOI22_X1  g660(.A1(new_n392_), .A2(new_n850_), .B1(new_n859_), .B2(new_n861_), .ZN(G1340gat));
  XNOR2_X1  g661(.A(KEYINPUT125), .B(G120gat), .ZN(new_n863_));
  OR2_X1    g662(.A1(new_n863_), .A2(KEYINPUT60), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n578_), .B2(KEYINPUT60), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n842_), .A2(new_n849_), .A3(new_n864_), .A4(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n867_), .B1(new_n847_), .B2(new_n840_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n858_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n869_), .B1(new_n854_), .B2(new_n856_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n868_), .A2(new_n870_), .A3(new_n578_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n866_), .B1(new_n871_), .B2(new_n863_), .ZN(G1341gat));
  INV_X1    g671(.A(G127gat), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n842_), .A2(new_n849_), .A3(new_n619_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n620_), .A2(KEYINPUT126), .ZN(new_n875_));
  MUX2_X1   g674(.A(KEYINPUT126), .B(new_n875_), .S(G127gat), .Z(new_n876_));
  AOI22_X1  g675(.A1(new_n873_), .A2(new_n874_), .B1(new_n859_), .B2(new_n876_), .ZN(G1342gat));
  INV_X1    g676(.A(G134gat), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n842_), .A2(new_n849_), .A3(new_n640_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(KEYINPUT127), .B(G134gat), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n677_), .A2(new_n880_), .ZN(new_n881_));
  AOI22_X1  g680(.A1(new_n878_), .A2(new_n879_), .B1(new_n859_), .B2(new_n881_), .ZN(G1343gat));
  NAND2_X1  g681(.A1(new_n384_), .A2(new_n478_), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n341_), .A2(new_n627_), .A3(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n847_), .A2(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n886_), .A2(new_n354_), .A3(new_n520_), .ZN(new_n887_));
  OAI21_X1  g686(.A(G141gat), .B1(new_n885_), .B2(new_n519_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(G1344gat));
  NAND3_X1  g688(.A1(new_n886_), .A2(new_n355_), .A3(new_n668_), .ZN(new_n890_));
  OAI21_X1  g689(.A(G148gat), .B1(new_n885_), .B2(new_n578_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(G1345gat));
  XNOR2_X1  g691(.A(KEYINPUT61), .B(G155gat), .ZN(new_n893_));
  OR3_X1    g692(.A1(new_n885_), .A2(new_n620_), .A3(new_n893_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n885_), .B2(new_n620_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1346gat));
  OR3_X1    g695(.A1(new_n885_), .A2(G162gat), .A3(new_n642_), .ZN(new_n897_));
  OAI21_X1  g696(.A(G162gat), .B1(new_n885_), .B2(new_n677_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(G1347gat));
  INV_X1    g698(.A(KEYINPUT62), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n628_), .A2(new_n478_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n341_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n902_), .A2(new_n384_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n903_), .ZN(new_n904_));
  AOI211_X1 g703(.A(new_n519_), .B(new_n904_), .C1(new_n854_), .C2(new_n856_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n900_), .B1(new_n905_), .B2(new_n223_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n257_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n857_), .A2(new_n520_), .A3(new_n903_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n908_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n906_), .A2(new_n907_), .A3(new_n909_), .ZN(G1348gat));
  AOI21_X1  g709(.A(new_n904_), .B1(new_n854_), .B2(new_n856_), .ZN(new_n911_));
  AOI21_X1  g710(.A(G176gat), .B1(new_n911_), .B2(new_n668_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n839_), .A2(new_n384_), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n902_), .A2(new_n578_), .A3(new_n224_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n912_), .B1(new_n913_), .B2(new_n914_), .ZN(G1349gat));
  NAND4_X1  g714(.A1(new_n913_), .A2(new_n341_), .A3(new_n619_), .A4(new_n901_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n620_), .A2(new_n272_), .ZN(new_n917_));
  AOI22_X1  g716(.A1(new_n916_), .A2(new_n208_), .B1(new_n911_), .B2(new_n917_), .ZN(G1350gat));
  NAND3_X1  g717(.A1(new_n911_), .A2(new_n218_), .A3(new_n640_), .ZN(new_n919_));
  AND2_X1   g718(.A1(new_n911_), .A2(new_n603_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n919_), .B1(new_n920_), .B2(new_n209_), .ZN(G1351gat));
  NOR3_X1   g720(.A1(new_n730_), .A2(new_n429_), .A3(new_n883_), .ZN(new_n922_));
  AND2_X1   g721(.A1(new_n847_), .A2(new_n922_), .ZN(new_n923_));
  AOI21_X1  g722(.A(G197gat), .B1(new_n923_), .B2(new_n520_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n847_), .A2(new_n922_), .ZN(new_n925_));
  NOR3_X1   g724(.A1(new_n925_), .A2(new_n244_), .A3(new_n519_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n924_), .A2(new_n926_), .ZN(G1352gat));
  NAND3_X1  g726(.A1(new_n923_), .A2(new_n242_), .A3(new_n668_), .ZN(new_n928_));
  OAI21_X1  g727(.A(G204gat), .B1(new_n925_), .B2(new_n578_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(G1353gat));
  OR2_X1    g729(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n620_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n932_));
  AND3_X1   g731(.A1(new_n923_), .A2(new_n931_), .A3(new_n932_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n931_), .B1(new_n923_), .B2(new_n932_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n933_), .A2(new_n934_), .ZN(G1354gat));
  NAND3_X1  g734(.A1(new_n923_), .A2(new_n236_), .A3(new_n640_), .ZN(new_n936_));
  OAI21_X1  g735(.A(G218gat), .B1(new_n925_), .B2(new_n677_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n936_), .A2(new_n937_), .ZN(G1355gat));
endmodule


