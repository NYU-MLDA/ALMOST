//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 0 1 0 1 0 0 1 1 0 0 1 0 1 1 1 0 1 1 1 1 1 1 1 1 1 1 0 1 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n800_, new_n801_, new_n803_,
    new_n804_, new_n805_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n883_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n909_, new_n911_, new_n912_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n933_, new_n934_,
    new_n936_, new_n937_, new_n939_, new_n940_, new_n941_, new_n943_,
    new_n944_, new_n946_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n953_, new_n954_, new_n955_;
  XNOR2_X1  g000(.A(KEYINPUT81), .B(G183gat), .ZN(new_n202_));
  INV_X1    g001(.A(G190gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G183gat), .A2(G190gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT23), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT87), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n205_), .A2(KEYINPUT87), .A3(KEYINPUT23), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT83), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT83), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT23), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n205_), .B1(new_n212_), .B2(new_n214_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n204_), .B1(new_n210_), .B2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(G176gat), .ZN(new_n217_));
  AND2_X1   g016(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n219_));
  OAI211_X1 g018(.A(KEYINPUT85), .B(new_n217_), .C1(new_n218_), .C2(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(KEYINPUT85), .A2(KEYINPUT22), .ZN(new_n221_));
  OAI21_X1  g020(.A(G169gat), .B1(new_n221_), .B2(G176gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT86), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n220_), .A2(KEYINPUT86), .A3(new_n222_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n216_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT82), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G169gat), .A2(G176gat), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n229_), .A2(new_n230_), .A3(KEYINPUT24), .A4(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(KEYINPUT24), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT82), .B1(new_n233_), .B2(new_n228_), .ZN(new_n234_));
  AND2_X1   g033(.A1(new_n232_), .A2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT26), .B(G190gat), .ZN(new_n236_));
  AND2_X1   g035(.A1(KEYINPUT81), .A2(G183gat), .ZN(new_n237_));
  NOR2_X1   g036(.A1(KEYINPUT81), .A2(G183gat), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT25), .ZN(new_n239_));
  NOR3_X1   g038(.A1(new_n237_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n236_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n229_), .A2(KEYINPUT24), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n212_), .A2(new_n214_), .A3(new_n205_), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT84), .B1(new_n205_), .B2(KEYINPUT23), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT84), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n247_), .A2(new_n211_), .A3(G183gat), .A4(G190gat), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n245_), .A2(new_n246_), .A3(new_n248_), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n235_), .A2(new_n242_), .A3(new_n244_), .A4(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n227_), .A2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT30), .ZN(new_n252_));
  XOR2_X1   g051(.A(G71gat), .B(G99gat), .Z(new_n253_));
  XNOR2_X1  g052(.A(new_n252_), .B(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT88), .ZN(new_n255_));
  AND2_X1   g054(.A1(G127gat), .A2(G134gat), .ZN(new_n256_));
  NOR2_X1   g055(.A1(G127gat), .A2(G134gat), .ZN(new_n257_));
  OAI21_X1  g056(.A(G113gat), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(G127gat), .ZN(new_n259_));
  INV_X1    g058(.A(G134gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(G113gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G127gat), .A2(G134gat), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n261_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  AND3_X1   g063(.A1(new_n258_), .A2(new_n264_), .A3(G120gat), .ZN(new_n265_));
  AOI21_X1  g064(.A(G120gat), .B1(new_n258_), .B2(new_n264_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n255_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(G120gat), .ZN(new_n268_));
  NOR3_X1   g067(.A1(new_n256_), .A2(new_n257_), .A3(G113gat), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n262_), .B1(new_n261_), .B2(new_n263_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n268_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n258_), .A2(new_n264_), .A3(G120gat), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(KEYINPUT88), .A3(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n267_), .A2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT31), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n254_), .B(new_n275_), .ZN(new_n276_));
  XOR2_X1   g075(.A(G15gat), .B(G43gat), .Z(new_n277_));
  NAND2_X1  g076(.A1(G227gat), .A2(G233gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  OR2_X1    g078(.A1(new_n276_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n276_), .A2(new_n279_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  AND2_X1   g082(.A1(G155gat), .A2(G162gat), .ZN(new_n284_));
  NOR2_X1   g083(.A1(G155gat), .A2(G162gat), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT1), .ZN(new_n287_));
  INV_X1    g086(.A(G141gat), .ZN(new_n288_));
  INV_X1    g087(.A(G148gat), .ZN(new_n289_));
  AOI22_X1  g088(.A1(new_n286_), .A2(new_n287_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  AOI22_X1  g089(.A1(new_n284_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT2), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n292_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT3), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n294_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n296_));
  NAND3_X1  g095(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n293_), .A2(new_n295_), .A3(new_n296_), .A4(new_n297_), .ZN(new_n298_));
  AOI22_X1  g097(.A1(new_n290_), .A2(new_n291_), .B1(new_n298_), .B2(new_n286_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n299_), .B1(new_n267_), .B2(new_n273_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n290_), .A2(new_n291_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n298_), .A2(new_n286_), .ZN(new_n302_));
  AND4_X1   g101(.A1(new_n301_), .A2(new_n302_), .A3(new_n272_), .A4(new_n271_), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT4), .B1(new_n300_), .B2(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n304_), .B1(KEYINPUT4), .B2(new_n300_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G225gat), .A2(G233gat), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n299_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n274_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n303_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n310_), .A2(new_n306_), .A3(new_n311_), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n308_), .A2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT0), .B(G57gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(G85gat), .ZN(new_n315_));
  XOR2_X1   g114(.A(G1gat), .B(G29gat), .Z(new_n316_));
  XOR2_X1   g115(.A(new_n315_), .B(new_n316_), .Z(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n313_), .B(new_n318_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n283_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT20), .ZN(new_n321_));
  AND3_X1   g120(.A1(new_n220_), .A2(KEYINPUT86), .A3(new_n222_), .ZN(new_n322_));
  AOI21_X1  g121(.A(KEYINPUT86), .B1(new_n220_), .B2(new_n222_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  AND3_X1   g123(.A1(new_n249_), .A2(new_n234_), .A3(new_n232_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n241_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n326_), .B1(new_n202_), .B2(new_n239_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n243_), .B1(new_n327_), .B2(new_n236_), .ZN(new_n328_));
  AOI22_X1  g127(.A1(new_n216_), .A2(new_n324_), .B1(new_n325_), .B2(new_n328_), .ZN(new_n329_));
  XOR2_X1   g128(.A(G211gat), .B(G218gat), .Z(new_n330_));
  INV_X1    g129(.A(G204gat), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n331_), .A2(G197gat), .ZN(new_n332_));
  INV_X1    g131(.A(G197gat), .ZN(new_n333_));
  OAI21_X1  g132(.A(KEYINPUT91), .B1(new_n333_), .B2(G204gat), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT91), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n335_), .A2(new_n331_), .A3(G197gat), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n332_), .B1(new_n334_), .B2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT21), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n330_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n333_), .A2(KEYINPUT90), .A3(G204gat), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n340_), .B1(new_n333_), .B2(G204gat), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n332_), .A2(KEYINPUT90), .ZN(new_n342_));
  OAI21_X1  g141(.A(KEYINPUT21), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n334_), .A2(new_n336_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n332_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n338_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  AOI22_X1  g145(.A1(new_n339_), .A2(new_n343_), .B1(new_n346_), .B2(new_n330_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n321_), .B1(new_n329_), .B2(new_n347_), .ZN(new_n348_));
  OR2_X1    g147(.A1(G183gat), .A2(G190gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n249_), .A2(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n217_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n351_));
  AOI21_X1  g150(.A(KEYINPUT96), .B1(new_n351_), .B2(new_n231_), .ZN(new_n352_));
  AND3_X1   g151(.A1(new_n351_), .A2(KEYINPUT96), .A3(new_n231_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n350_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(KEYINPUT97), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT96), .ZN(new_n356_));
  OR2_X1    g155(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n358_));
  AOI21_X1  g157(.A(G176gat), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n231_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n356_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n351_), .A2(KEYINPUT96), .A3(new_n231_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT97), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n363_), .A2(new_n364_), .A3(new_n350_), .ZN(new_n365_));
  AND3_X1   g164(.A1(new_n205_), .A2(KEYINPUT87), .A3(KEYINPUT23), .ZN(new_n366_));
  AOI21_X1  g165(.A(KEYINPUT87), .B1(new_n205_), .B2(KEYINPUT23), .ZN(new_n367_));
  NOR3_X1   g166(.A1(new_n215_), .A2(new_n366_), .A3(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(KEYINPUT95), .B1(new_n368_), .B2(new_n243_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(KEYINPUT83), .B(KEYINPUT23), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n208_), .B(new_n209_), .C1(new_n370_), .C2(new_n205_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT95), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n371_), .A2(new_n372_), .A3(new_n244_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n369_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT93), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n233_), .A2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n231_), .A2(KEYINPUT93), .A3(KEYINPUT24), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n376_), .A2(new_n229_), .A3(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(KEYINPUT25), .B(G183gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n236_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT94), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n378_), .A2(KEYINPUT94), .A3(new_n380_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  AOI22_X1  g184(.A1(new_n355_), .A2(new_n365_), .B1(new_n374_), .B2(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n348_), .B1(new_n386_), .B2(new_n347_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G226gat), .A2(G233gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(KEYINPUT19), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT106), .B1(new_n387_), .B2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n389_), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n371_), .A2(new_n372_), .A3(new_n244_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n372_), .B1(new_n371_), .B2(new_n244_), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n378_), .A2(KEYINPUT94), .A3(new_n380_), .ZN(new_n394_));
  AOI21_X1  g193(.A(KEYINPUT94), .B1(new_n378_), .B2(new_n380_), .ZN(new_n395_));
  OAI22_X1  g194(.A1(new_n392_), .A2(new_n393_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n396_), .A2(new_n347_), .A3(new_n354_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n347_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n321_), .B1(new_n251_), .B2(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n391_), .B1(new_n397_), .B2(new_n399_), .ZN(new_n400_));
  MUX2_X1   g199(.A(new_n390_), .B(KEYINPUT106), .S(new_n400_), .Z(new_n401_));
  XNOR2_X1  g200(.A(KEYINPUT18), .B(G64gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(G92gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G8gat), .B(G36gat), .ZN(new_n404_));
  XOR2_X1   g203(.A(new_n403_), .B(new_n404_), .Z(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n401_), .A2(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n364_), .B1(new_n363_), .B2(new_n350_), .ZN(new_n408_));
  AND3_X1   g207(.A1(new_n363_), .A2(new_n364_), .A3(new_n350_), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n396_), .B(new_n347_), .C1(new_n408_), .C2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n410_), .A2(new_n391_), .A3(new_n399_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT99), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n347_), .A2(new_n227_), .A3(new_n250_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT20), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n396_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n415_), .B1(new_n416_), .B2(new_n398_), .ZN(new_n417_));
  OAI21_X1  g216(.A(KEYINPUT98), .B1(new_n417_), .B2(new_n391_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT98), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n355_), .A2(new_n365_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n347_), .B1(new_n420_), .B2(new_n396_), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n419_), .B(new_n389_), .C1(new_n421_), .C2(new_n415_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n418_), .A2(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n413_), .A2(new_n423_), .A3(new_n405_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n407_), .A2(KEYINPUT27), .A3(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT27), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n413_), .A2(new_n405_), .A3(new_n423_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n405_), .B1(new_n413_), .B2(new_n423_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n426_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n425_), .A2(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n347_), .B1(KEYINPUT29), .B2(new_n309_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G228gat), .A2(G233gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n431_), .B(new_n432_), .ZN(new_n433_));
  XOR2_X1   g232(.A(G78gat), .B(G106gat), .Z(new_n434_));
  OR2_X1    g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(KEYINPUT89), .B1(new_n433_), .B2(new_n434_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n309_), .A2(KEYINPUT29), .ZN(new_n438_));
  XOR2_X1   g237(.A(G22gat), .B(G50gat), .Z(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(KEYINPUT28), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n438_), .B(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT92), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n441_), .B1(new_n442_), .B2(new_n434_), .ZN(new_n443_));
  AOI22_X1  g242(.A1(new_n437_), .A2(new_n441_), .B1(new_n436_), .B2(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n435_), .B1(new_n442_), .B2(new_n441_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n430_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n320_), .A2(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(KEYINPUT101), .A2(KEYINPUT33), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n300_), .A2(KEYINPUT4), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n310_), .A2(new_n311_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n450_), .B1(new_n451_), .B2(KEYINPUT4), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n312_), .B(new_n318_), .C1(new_n452_), .C2(new_n306_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(KEYINPUT101), .A2(KEYINPUT33), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n308_), .A2(new_n312_), .A3(new_n318_), .A4(new_n454_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT103), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n458_), .B1(new_n452_), .B2(new_n307_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT102), .ZN(new_n460_));
  NOR3_X1   g259(.A1(new_n300_), .A2(new_n306_), .A3(new_n303_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n460_), .B1(new_n461_), .B2(new_n318_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n310_), .A2(new_n307_), .A3(new_n311_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n463_), .A2(KEYINPUT102), .A3(new_n317_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n305_), .A2(KEYINPUT103), .A3(new_n306_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n459_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT104), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT104), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n459_), .A2(new_n465_), .A3(new_n469_), .A4(new_n466_), .ZN(new_n470_));
  AOI221_X4 g269(.A(new_n449_), .B1(new_n456_), .B2(new_n457_), .C1(new_n468_), .C2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT100), .ZN(new_n472_));
  NOR3_X1   g271(.A1(new_n427_), .A2(new_n428_), .A3(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n422_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n419_), .B1(new_n387_), .B2(new_n389_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n411_), .B(KEYINPUT99), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n406_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(KEYINPUT100), .B1(new_n478_), .B2(new_n424_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n471_), .B1(new_n473_), .B2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT105), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n401_), .A2(KEYINPUT32), .A3(new_n405_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n405_), .A2(KEYINPUT32), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n413_), .A2(new_n423_), .A3(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n483_), .A2(new_n319_), .A3(new_n485_), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n471_), .B(KEYINPUT105), .C1(new_n473_), .C2(new_n479_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n482_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n446_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n489_), .A2(new_n319_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n430_), .ZN(new_n491_));
  AOI22_X1  g290(.A1(new_n488_), .A2(new_n489_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n448_), .B1(new_n492_), .B2(new_n282_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT7), .ZN(new_n494_));
  INV_X1    g293(.A(G99gat), .ZN(new_n495_));
  INV_X1    g294(.A(G106gat), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n494_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G99gat), .A2(G106gat), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT6), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n497_), .A2(new_n500_), .A3(new_n501_), .A4(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT8), .ZN(new_n504_));
  OR2_X1    g303(.A1(G85gat), .A2(G92gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G85gat), .A2(G92gat), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  AND3_X1   g306(.A1(new_n503_), .A2(new_n504_), .A3(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n504_), .B1(new_n503_), .B2(new_n507_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(KEYINPUT10), .B(G99gat), .ZN(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT64), .B1(new_n510_), .B2(G106gat), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT64), .ZN(new_n512_));
  AND2_X1   g311(.A1(new_n495_), .A2(KEYINPUT10), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n495_), .A2(KEYINPUT10), .ZN(new_n514_));
  OAI211_X1 g313(.A(new_n512_), .B(new_n496_), .C1(new_n513_), .C2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n511_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT65), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT9), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n505_), .A2(new_n519_), .A3(new_n506_), .A4(new_n520_), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n517_), .A2(new_n518_), .A3(G85gat), .A4(G92gat), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n521_), .A2(new_n500_), .A3(new_n501_), .A4(new_n522_), .ZN(new_n523_));
  OAI22_X1  g322(.A1(new_n508_), .A2(new_n509_), .B1(new_n516_), .B2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT66), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  AND3_X1   g325(.A1(new_n522_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n511_), .A2(new_n527_), .A3(new_n515_), .A4(new_n521_), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n528_), .B(KEYINPUT66), .C1(new_n508_), .C2(new_n509_), .ZN(new_n529_));
  XOR2_X1   g328(.A(G57gat), .B(G64gat), .Z(new_n530_));
  INV_X1    g329(.A(KEYINPUT11), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G57gat), .B(G64gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT11), .ZN(new_n534_));
  XOR2_X1   g333(.A(G71gat), .B(G78gat), .Z(new_n535_));
  NAND3_X1  g334(.A1(new_n532_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n534_), .A2(new_n535_), .ZN(new_n537_));
  AND2_X1   g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n526_), .A2(new_n529_), .A3(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT12), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n524_), .A2(new_n538_), .A3(KEYINPUT12), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT67), .ZN(new_n543_));
  OR2_X1    g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(new_n543_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n541_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT68), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n538_), .B1(new_n526_), .B2(new_n529_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G230gat), .A2(G233gat), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n547_), .B1(new_n548_), .B2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n526_), .A2(new_n529_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n538_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n554_), .A2(KEYINPUT68), .A3(new_n549_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n546_), .B1(new_n551_), .B2(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n549_), .B1(new_n554_), .B2(new_n539_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G120gat), .B(G148gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(new_n331_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT5), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(new_n217_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n558_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(KEYINPUT69), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n564_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  XOR2_X1   g365(.A(KEYINPUT70), .B(KEYINPUT13), .Z(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT13), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n563_), .B(new_n565_), .C1(KEYINPUT70), .C2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(KEYINPUT71), .B(G43gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(G50gat), .ZN(new_n574_));
  XOR2_X1   g373(.A(G29gat), .B(G36gat), .Z(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n574_), .B(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT79), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(KEYINPUT76), .B(G22gat), .ZN(new_n580_));
  INV_X1    g379(.A(G15gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(G1gat), .ZN(new_n583_));
  INV_X1    g382(.A(G8gat), .ZN(new_n584_));
  OAI21_X1  g383(.A(KEYINPUT14), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n582_), .A2(new_n585_), .ZN(new_n586_));
  XOR2_X1   g385(.A(G1gat), .B(G8gat), .Z(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n586_), .B(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n579_), .A2(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n577_), .B(KEYINPUT15), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(new_n589_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G229gat), .A2(G233gat), .ZN(new_n594_));
  AND3_X1   g393(.A1(new_n591_), .A2(new_n593_), .A3(new_n594_), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n577_), .A2(KEYINPUT79), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n577_), .A2(KEYINPUT79), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(new_n589_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n594_), .B1(new_n599_), .B2(new_n591_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G113gat), .B(G141gat), .ZN(new_n601_));
  INV_X1    g400(.A(G169gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(new_n333_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n605_), .A2(KEYINPUT80), .ZN(new_n606_));
  NOR3_X1   g405(.A1(new_n595_), .A2(new_n600_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n606_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n594_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n598_), .A2(new_n589_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n579_), .A2(new_n590_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n609_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n591_), .A2(new_n593_), .A3(new_n594_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n608_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n607_), .A2(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n572_), .A2(new_n615_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n493_), .A2(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n589_), .B(new_n538_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(G231gat), .A2(G233gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  XOR2_X1   g419(.A(G127gat), .B(G155gat), .Z(new_n621_));
  XNOR2_X1  g420(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  XOR2_X1   g422(.A(G183gat), .B(G211gat), .Z(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  AND3_X1   g424(.A1(new_n620_), .A2(KEYINPUT17), .A3(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(KEYINPUT17), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n620_), .A2(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n626_), .A2(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT78), .ZN(new_n630_));
  NAND2_X1  g429(.A1(G232gat), .A2(G233gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT34), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n632_), .A2(KEYINPUT35), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n633_), .B1(new_n592_), .B2(new_n524_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n632_), .A2(KEYINPUT73), .A3(KEYINPUT35), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT72), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n636_), .B1(new_n552_), .B2(new_n577_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n552_), .A2(new_n577_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n638_), .A2(KEYINPUT72), .ZN(new_n639_));
  OAI211_X1 g438(.A(new_n634_), .B(new_n635_), .C1(new_n637_), .C2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n632_), .A2(KEYINPUT35), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT73), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n640_), .A2(new_n644_), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n639_), .A2(new_n637_), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n646_), .A2(new_n643_), .A3(new_n635_), .A4(new_n634_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(G190gat), .B(G218gat), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(G134gat), .ZN(new_n649_));
  INV_X1    g448(.A(G162gat), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT36), .ZN(new_n652_));
  AND3_X1   g451(.A1(new_n645_), .A2(new_n647_), .A3(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT36), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n651_), .A2(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n655_), .B1(new_n645_), .B2(new_n647_), .ZN(new_n656_));
  OAI21_X1  g455(.A(KEYINPUT74), .B1(new_n653_), .B2(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n645_), .A2(new_n647_), .A3(new_n652_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT74), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n657_), .A2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(KEYINPUT37), .ZN(new_n662_));
  INV_X1    g461(.A(new_n645_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n640_), .A2(new_n644_), .ZN(new_n664_));
  OAI21_X1  g463(.A(KEYINPUT75), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT75), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n645_), .A2(new_n647_), .A3(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n665_), .A2(new_n652_), .A3(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT37), .ZN(new_n669_));
  INV_X1    g468(.A(new_n656_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n668_), .A2(new_n669_), .A3(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n630_), .B1(new_n662_), .B2(new_n671_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n617_), .A2(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n673_), .A2(new_n583_), .A3(new_n319_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT38), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n668_), .A2(new_n670_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n617_), .A2(new_n676_), .A3(new_n629_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n319_), .ZN(new_n678_));
  OAI21_X1  g477(.A(G1gat), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n675_), .A2(new_n679_), .ZN(G1324gat));
  INV_X1    g479(.A(KEYINPUT107), .ZN(new_n681_));
  OR3_X1    g480(.A1(new_n677_), .A2(new_n681_), .A3(new_n491_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n681_), .B1(new_n677_), .B2(new_n491_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n682_), .A2(G8gat), .A3(new_n683_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT39), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n673_), .A2(new_n584_), .A3(new_n430_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT40), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n685_), .A2(KEYINPUT40), .A3(new_n686_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(G1325gat));
  OAI21_X1  g490(.A(G15gat), .B1(new_n677_), .B2(new_n283_), .ZN(new_n692_));
  XOR2_X1   g491(.A(new_n692_), .B(KEYINPUT41), .Z(new_n693_));
  NAND3_X1  g492(.A1(new_n673_), .A2(new_n581_), .A3(new_n282_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(G1326gat));
  OAI21_X1  g494(.A(G22gat), .B1(new_n677_), .B2(new_n489_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT42), .ZN(new_n697_));
  INV_X1    g496(.A(G22gat), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n673_), .A2(new_n698_), .A3(new_n446_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n697_), .A2(new_n699_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT108), .ZN(G1327gat));
  INV_X1    g500(.A(KEYINPUT78), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n629_), .B(new_n702_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n703_), .A2(new_n676_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n617_), .A2(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(G29gat), .B1(new_n705_), .B2(new_n319_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT43), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n668_), .A2(new_n669_), .A3(new_n670_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n669_), .B1(new_n657_), .B2(new_n660_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n488_), .A2(new_n489_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n491_), .A2(new_n490_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n282_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n448_), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n707_), .B(new_n710_), .C1(new_n713_), .C2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT109), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n711_), .A2(new_n712_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n714_), .B1(new_n718_), .B2(new_n283_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n710_), .ZN(new_n720_));
  OAI21_X1  g519(.A(KEYINPUT43), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n493_), .A2(KEYINPUT109), .A3(new_n707_), .A4(new_n710_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n717_), .A2(new_n721_), .A3(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n723_), .A2(new_n616_), .A3(new_n630_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n723_), .A2(KEYINPUT44), .A3(new_n616_), .A4(new_n630_), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n726_), .A2(new_n319_), .A3(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n706_), .B1(new_n728_), .B2(G29gat), .ZN(G1328gat));
  NAND3_X1  g528(.A1(new_n726_), .A2(new_n430_), .A3(new_n727_), .ZN(new_n730_));
  INV_X1    g529(.A(G36gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n705_), .A2(new_n731_), .A3(new_n430_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(KEYINPUT45), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n732_), .A2(KEYINPUT45), .ZN(new_n734_));
  AOI22_X1  g533(.A1(new_n730_), .A2(G36gat), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT46), .ZN(new_n736_));
  OR2_X1    g535(.A1(new_n736_), .A2(KEYINPUT110), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(KEYINPUT110), .ZN(new_n738_));
  AND3_X1   g537(.A1(new_n735_), .A2(new_n737_), .A3(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n737_), .B1(new_n735_), .B2(new_n738_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n739_), .A2(new_n740_), .ZN(G1329gat));
  INV_X1    g540(.A(G43gat), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n283_), .A2(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n726_), .A2(new_n727_), .A3(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT111), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT111), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n726_), .A2(new_n746_), .A3(new_n727_), .A4(new_n743_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n705_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n742_), .B1(new_n749_), .B2(new_n283_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT47), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT47), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n748_), .A2(new_n753_), .A3(new_n750_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n752_), .A2(new_n754_), .ZN(G1330gat));
  AND4_X1   g554(.A1(G50gat), .A2(new_n726_), .A3(new_n446_), .A4(new_n727_), .ZN(new_n756_));
  AOI21_X1  g555(.A(G50gat), .B1(new_n705_), .B2(new_n446_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n756_), .A2(new_n757_), .ZN(G1331gat));
  INV_X1    g557(.A(new_n672_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n759_), .A2(KEYINPUT112), .A3(new_n571_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n615_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(KEYINPUT112), .B1(new_n759_), .B2(new_n571_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n762_), .A2(new_n493_), .A3(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(G57gat), .B1(new_n765_), .B2(new_n319_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n571_), .A2(new_n761_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n493_), .A2(new_n767_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n768_), .A2(new_n676_), .A3(new_n703_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT113), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n770_), .A2(new_n319_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n766_), .B1(new_n771_), .B2(G57gat), .ZN(G1332gat));
  INV_X1    g571(.A(G64gat), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n765_), .A2(new_n773_), .A3(new_n430_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT48), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n770_), .A2(new_n430_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n776_), .B2(G64gat), .ZN(new_n777_));
  AOI211_X1 g576(.A(KEYINPUT48), .B(new_n773_), .C1(new_n770_), .C2(new_n430_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n774_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT114), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT114), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n781_), .B(new_n774_), .C1(new_n777_), .C2(new_n778_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(G1333gat));
  INV_X1    g582(.A(G71gat), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n784_), .B1(new_n770_), .B2(new_n282_), .ZN(new_n785_));
  XOR2_X1   g584(.A(new_n785_), .B(KEYINPUT49), .Z(new_n786_));
  NAND3_X1  g585(.A1(new_n765_), .A2(new_n784_), .A3(new_n282_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(G1334gat));
  INV_X1    g587(.A(G78gat), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n789_), .B1(new_n770_), .B2(new_n446_), .ZN(new_n790_));
  XOR2_X1   g589(.A(new_n790_), .B(KEYINPUT50), .Z(new_n791_));
  NAND3_X1  g590(.A1(new_n765_), .A2(new_n789_), .A3(new_n446_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(G1335gat));
  NAND2_X1  g592(.A1(new_n768_), .A2(new_n704_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(G85gat), .B1(new_n795_), .B2(new_n319_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n723_), .A2(new_n630_), .A3(new_n767_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n797_), .A2(new_n678_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n796_), .B1(new_n798_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g598(.A(G92gat), .B1(new_n795_), .B2(new_n430_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n797_), .A2(new_n491_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n800_), .B1(new_n801_), .B2(G92gat), .ZN(G1337gat));
  OAI21_X1  g601(.A(G99gat), .B1(new_n797_), .B2(new_n283_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n282_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n803_), .B1(new_n794_), .B2(new_n804_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n805_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g605(.A1(new_n795_), .A2(new_n496_), .A3(new_n446_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n723_), .A2(new_n446_), .A3(new_n630_), .A4(new_n767_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT52), .ZN(new_n809_));
  AND3_X1   g608(.A1(new_n808_), .A2(new_n809_), .A3(G106gat), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n809_), .B1(new_n808_), .B2(G106gat), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n807_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n812_), .B(KEYINPUT53), .ZN(G1339gat));
  OAI211_X1 g612(.A(new_n615_), .B(new_n703_), .C1(new_n708_), .C2(new_n709_), .ZN(new_n814_));
  OAI21_X1  g613(.A(KEYINPUT54), .B1(new_n814_), .B2(new_n572_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n672_), .A2(new_n816_), .A3(new_n615_), .A4(new_n571_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n815_), .A2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n609_), .B1(new_n599_), .B2(new_n591_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT117), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n820_), .A2(new_n821_), .A3(new_n604_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n591_), .A2(new_n593_), .A3(new_n609_), .ZN(new_n823_));
  OAI21_X1  g622(.A(KEYINPUT117), .B1(new_n819_), .B2(new_n605_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n822_), .A2(new_n823_), .A3(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n612_), .A2(new_n605_), .A3(new_n613_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT118), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n827_), .B(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(KEYINPUT55), .B1(new_n556_), .B2(KEYINPUT115), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT115), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT55), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n555_), .A2(new_n551_), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n831_), .B(new_n832_), .C1(new_n833_), .C2(new_n546_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n550_), .B1(new_n546_), .B2(new_n548_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n830_), .A2(new_n834_), .A3(new_n835_), .ZN(new_n836_));
  AND3_X1   g635(.A1(new_n836_), .A2(KEYINPUT56), .A3(new_n564_), .ZN(new_n837_));
  AOI21_X1  g636(.A(KEYINPUT56), .B1(new_n836_), .B2(new_n564_), .ZN(new_n838_));
  OR2_X1    g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n829_), .A2(new_n839_), .A3(new_n563_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT58), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n829_), .A2(new_n839_), .A3(KEYINPUT58), .A4(new_n563_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n842_), .A2(new_n710_), .A3(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n615_), .B1(new_n558_), .B2(new_n562_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n845_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(KEYINPUT116), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n827_), .A2(new_n828_), .ZN(new_n848_));
  AOI21_X1  g647(.A(KEYINPUT118), .B1(new_n825_), .B2(new_n826_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n566_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT116), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n845_), .B(new_n851_), .C1(new_n837_), .C2(new_n838_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n847_), .A2(new_n850_), .A3(new_n852_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(KEYINPUT119), .A2(KEYINPUT57), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n853_), .A2(new_n676_), .A3(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n854_), .B1(new_n853_), .B2(new_n676_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n844_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n629_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n818_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n447_), .A2(new_n319_), .A3(new_n282_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(G113gat), .B1(new_n864_), .B2(new_n761_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT121), .ZN(new_n866_));
  OAI21_X1  g665(.A(KEYINPUT59), .B1(new_n859_), .B2(new_n861_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(KEYINPUT120), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT120), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n869_), .B(KEYINPUT59), .C1(new_n859_), .C2(new_n861_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n868_), .A2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n857_), .A2(new_n630_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n818_), .ZN(new_n873_));
  AOI211_X1 g672(.A(KEYINPUT59), .B(new_n861_), .C1(new_n872_), .C2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n866_), .B1(new_n871_), .B2(new_n875_), .ZN(new_n876_));
  AOI211_X1 g675(.A(KEYINPUT121), .B(new_n874_), .C1(new_n868_), .C2(new_n870_), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n876_), .A2(new_n877_), .A3(new_n615_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n865_), .B1(new_n878_), .B2(G113gat), .ZN(G1340gat));
  NAND2_X1  g678(.A1(new_n871_), .A2(new_n875_), .ZN(new_n880_));
  OAI21_X1  g679(.A(G120gat), .B1(new_n880_), .B2(new_n571_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n268_), .B1(new_n571_), .B2(KEYINPUT60), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n864_), .B(new_n882_), .C1(KEYINPUT60), .C2(new_n268_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n881_), .A2(new_n883_), .ZN(G1341gat));
  INV_X1    g683(.A(KEYINPUT122), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n858_), .A2(new_n259_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n876_), .A2(new_n877_), .A3(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(G127gat), .B1(new_n864_), .B2(new_n703_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n885_), .B1(new_n888_), .B2(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n880_), .A2(KEYINPUT121), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n871_), .A2(new_n866_), .A3(new_n875_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n891_), .A2(new_n892_), .A3(new_n886_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n889_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n893_), .A2(KEYINPUT122), .A3(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n890_), .A2(new_n895_), .ZN(G1342gat));
  INV_X1    g695(.A(new_n676_), .ZN(new_n897_));
  AOI21_X1  g696(.A(G134gat), .B1(new_n864_), .B2(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n876_), .A2(new_n877_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n720_), .A2(new_n260_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n898_), .B1(new_n899_), .B2(new_n900_), .ZN(G1343gat));
  NOR4_X1   g700(.A1(new_n282_), .A2(new_n430_), .A3(new_n489_), .A4(new_n678_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(KEYINPUT123), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n860_), .A2(new_n903_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(KEYINPUT124), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(new_n761_), .ZN(new_n906_));
  XOR2_X1   g705(.A(KEYINPUT125), .B(G141gat), .Z(new_n907_));
  XNOR2_X1  g706(.A(new_n906_), .B(new_n907_), .ZN(G1344gat));
  NAND2_X1  g707(.A1(new_n905_), .A2(new_n572_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g709(.A1(new_n905_), .A2(new_n703_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(KEYINPUT61), .B(G155gat), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n911_), .B(new_n912_), .ZN(G1346gat));
  INV_X1    g712(.A(KEYINPUT126), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n905_), .A2(new_n650_), .A3(new_n897_), .ZN(new_n915_));
  AND2_X1   g714(.A1(new_n905_), .A2(new_n710_), .ZN(new_n916_));
  OAI211_X1 g715(.A(new_n914_), .B(new_n915_), .C1(new_n916_), .C2(new_n650_), .ZN(new_n917_));
  AND3_X1   g716(.A1(new_n905_), .A2(new_n650_), .A3(new_n897_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n650_), .B1(new_n905_), .B2(new_n710_), .ZN(new_n919_));
  OAI21_X1  g718(.A(KEYINPUT126), .B1(new_n918_), .B2(new_n919_), .ZN(new_n920_));
  AND2_X1   g719(.A1(new_n917_), .A2(new_n920_), .ZN(G1347gat));
  AOI21_X1  g720(.A(new_n446_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n320_), .A2(new_n430_), .ZN(new_n923_));
  INV_X1    g722(.A(new_n923_), .ZN(new_n924_));
  AND2_X1   g723(.A1(new_n922_), .A2(new_n924_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n602_), .B1(new_n925_), .B2(new_n761_), .ZN(new_n926_));
  OR2_X1    g725(.A1(new_n926_), .A2(KEYINPUT62), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n926_), .A2(KEYINPUT62), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n218_), .A2(new_n219_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n925_), .A2(new_n761_), .ZN(new_n930_));
  OAI211_X1 g729(.A(new_n927_), .B(new_n928_), .C1(new_n929_), .C2(new_n930_), .ZN(G1348gat));
  AOI21_X1  g730(.A(G176gat), .B1(new_n925_), .B2(new_n572_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n859_), .A2(new_n446_), .ZN(new_n933_));
  NOR3_X1   g732(.A1(new_n923_), .A2(new_n571_), .A3(new_n217_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n932_), .B1(new_n933_), .B2(new_n934_), .ZN(G1349gat));
  NOR2_X1   g734(.A1(new_n858_), .A2(new_n379_), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n933_), .A2(new_n703_), .A3(new_n924_), .ZN(new_n937_));
  AOI22_X1  g736(.A1(new_n925_), .A2(new_n936_), .B1(new_n937_), .B2(new_n202_), .ZN(G1350gat));
  INV_X1    g737(.A(new_n925_), .ZN(new_n939_));
  OAI21_X1  g738(.A(G190gat), .B1(new_n939_), .B2(new_n720_), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n925_), .A2(new_n897_), .A3(new_n236_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n940_), .A2(new_n941_), .ZN(G1351gat));
  AND4_X1   g741(.A1(new_n490_), .A2(new_n860_), .A3(new_n430_), .A4(new_n283_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n943_), .A2(new_n761_), .ZN(new_n944_));
  XNOR2_X1  g743(.A(new_n944_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g744(.A1(new_n943_), .A2(new_n572_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g746(.A1(new_n943_), .A2(new_n629_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n949_));
  AND2_X1   g748(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n950_));
  NOR3_X1   g749(.A1(new_n948_), .A2(new_n949_), .A3(new_n950_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n951_), .B1(new_n948_), .B2(new_n949_), .ZN(G1354gat));
  AOI21_X1  g751(.A(G218gat), .B1(new_n943_), .B2(new_n897_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n710_), .A2(G218gat), .ZN(new_n954_));
  XOR2_X1   g753(.A(new_n954_), .B(KEYINPUT127), .Z(new_n955_));
  AOI21_X1  g754(.A(new_n953_), .B1(new_n943_), .B2(new_n955_), .ZN(G1355gat));
endmodule


