//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 0 0 0 0 1 0 0 1 0 1 0 0 0 1 1 1 1 0 0 1 0 1 1 1 0 1 1 0 0 1 1 0 1 0 0 0 0 1 0 0 1 1 1 0 0 1 1 1 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n631_, new_n632_, new_n633_, new_n634_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n808_, new_n809_, new_n811_, new_n812_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n821_, new_n823_,
    new_n824_, new_n826_, new_n827_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n838_,
    new_n839_, new_n840_, new_n842_, new_n843_, new_n845_, new_n846_,
    new_n847_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n870_, new_n871_;
  NAND2_X1  g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT81), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT81), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n204_), .A2(G169gat), .A3(G176gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G183gat), .ZN(new_n207_));
  INV_X1    g006(.A(G190gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT23), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT86), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n207_), .A2(KEYINPUT23), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n210_), .B1(new_n211_), .B2(G190gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT23), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n213_), .A2(G183gat), .A3(G190gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n214_), .A2(KEYINPUT86), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n209_), .B1(new_n212_), .B2(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(G183gat), .A2(G190gat), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n206_), .B1(new_n216_), .B2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(G169gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT22), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT84), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(G176gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT22), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(G169gat), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n222_), .B1(new_n221_), .B2(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT85), .B1(new_n225_), .B2(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(G176gat), .B1(new_n221_), .B2(new_n222_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT85), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT22), .B(G169gat), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n230_), .B(new_n231_), .C1(new_n222_), .C2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n229_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT82), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n209_), .B(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT83), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n214_), .B(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n236_), .A2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(KEYINPUT25), .B(G183gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT26), .B(G190gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n220_), .A2(new_n224_), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n243_), .A2(KEYINPUT24), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n203_), .A2(new_n205_), .A3(new_n243_), .A4(KEYINPUT24), .ZN(new_n245_));
  AND3_X1   g044(.A1(new_n242_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  AOI22_X1  g045(.A1(new_n219_), .A2(new_n234_), .B1(new_n239_), .B2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT30), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G227gat), .A2(G233gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT87), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G71gat), .B(G99gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n250_), .B(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n248_), .B(new_n252_), .ZN(new_n253_));
  XOR2_X1   g052(.A(KEYINPUT88), .B(KEYINPUT31), .Z(new_n254_));
  XNOR2_X1  g053(.A(new_n253_), .B(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(G134gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(G127gat), .ZN(new_n257_));
  INV_X1    g056(.A(G127gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(G134gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(G120gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(G113gat), .ZN(new_n262_));
  INV_X1    g061(.A(G113gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(G120gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n260_), .A2(new_n265_), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n257_), .A2(new_n259_), .A3(new_n262_), .A4(new_n264_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  XOR2_X1   g067(.A(G15gat), .B(G43gat), .Z(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  XOR2_X1   g069(.A(new_n255_), .B(new_n270_), .Z(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT27), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G226gat), .A2(G233gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT19), .ZN(new_n275_));
  AND2_X1   g074(.A1(KEYINPUT90), .A2(G204gat), .ZN(new_n276_));
  NOR2_X1   g075(.A1(KEYINPUT90), .A2(G204gat), .ZN(new_n277_));
  OAI21_X1  g076(.A(G197gat), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n278_), .B1(G197gat), .B2(G204gat), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT21), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G211gat), .B(G218gat), .ZN(new_n281_));
  NOR3_X1   g080(.A1(new_n279_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n281_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n284_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT91), .ZN(new_n286_));
  NOR3_X1   g085(.A1(new_n276_), .A2(new_n277_), .A3(G197gat), .ZN(new_n287_));
  INV_X1    g086(.A(G197gat), .ZN(new_n288_));
  INV_X1    g087(.A(G204gat), .ZN(new_n289_));
  OAI21_X1  g088(.A(KEYINPUT21), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n286_), .B1(new_n287_), .B2(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n280_), .B1(G197gat), .B2(G204gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT90), .B(G204gat), .ZN(new_n293_));
  OAI211_X1 g092(.A(KEYINPUT91), .B(new_n292_), .C1(new_n293_), .C2(G197gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n291_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT92), .ZN(new_n296_));
  AND3_X1   g095(.A1(new_n285_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n296_), .B1(new_n285_), .B2(new_n295_), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n247_), .B(new_n283_), .C1(new_n297_), .C2(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n299_), .A2(KEYINPUT95), .A3(KEYINPUT20), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n283_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n239_), .A2(new_n218_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n206_), .B1(new_n224_), .B2(new_n232_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n243_), .A2(KEYINPUT24), .A3(new_n202_), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n216_), .A2(new_n242_), .A3(new_n244_), .A4(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n301_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n300_), .A2(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(KEYINPUT95), .B1(new_n299_), .B2(KEYINPUT20), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n275_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(KEYINPUT20), .B1(new_n301_), .B2(new_n307_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n285_), .A2(new_n295_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT92), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n285_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n282_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n316_), .A2(new_n247_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n312_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n275_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G8gat), .B(G36gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT18), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(G64gat), .ZN(new_n323_));
  INV_X1    g122(.A(G92gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n311_), .A2(new_n320_), .A3(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n325_), .B1(new_n311_), .B2(new_n320_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n326_), .B1(new_n327_), .B2(KEYINPUT96), .ZN(new_n328_));
  NOR3_X1   g127(.A1(new_n312_), .A2(new_n317_), .A3(new_n275_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n299_), .A2(KEYINPUT20), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT95), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n332_), .A2(new_n308_), .A3(new_n300_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n329_), .B1(new_n333_), .B2(new_n275_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT96), .ZN(new_n335_));
  NOR3_X1   g134(.A1(new_n334_), .A2(new_n335_), .A3(new_n325_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n273_), .B1(new_n328_), .B2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G78gat), .B(G106gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT94), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  AND2_X1   g139(.A1(G228gat), .A2(G233gat), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n341_), .B1(new_n316_), .B2(KEYINPUT93), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G155gat), .B(G162gat), .ZN(new_n343_));
  NOR3_X1   g142(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n344_));
  AND3_X1   g143(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n345_));
  AOI21_X1  g144(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n346_));
  NOR3_X1   g145(.A1(new_n344_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT89), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  OAI211_X1 g149(.A(KEYINPUT89), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n343_), .B1(new_n347_), .B2(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n343_), .A2(KEYINPUT1), .ZN(new_n354_));
  INV_X1    g153(.A(G141gat), .ZN(new_n355_));
  INV_X1    g154(.A(G148gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G141gat), .A2(G148gat), .ZN(new_n358_));
  NAND3_X1  g157(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n357_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n354_), .A2(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n353_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT29), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G22gat), .B(G50gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT28), .ZN(new_n365_));
  AND3_X1   g164(.A1(new_n362_), .A2(new_n363_), .A3(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n365_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n342_), .A2(new_n369_), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n368_), .B(new_n341_), .C1(new_n316_), .C2(KEYINPUT93), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n301_), .B1(new_n363_), .B2(new_n362_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n370_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n372_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n340_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n370_), .A2(new_n371_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n372_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n379_), .A2(new_n339_), .A3(new_n373_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n376_), .A2(new_n380_), .ZN(new_n381_));
  AND2_X1   g180(.A1(new_n357_), .A2(new_n358_), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n382_), .B(new_n359_), .C1(KEYINPUT1), .C2(new_n343_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT3), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n384_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT2), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n358_), .A2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n385_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n389_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n268_), .B(new_n383_), .C1(new_n390_), .C2(new_n343_), .ZN(new_n391_));
  AND2_X1   g190(.A1(new_n266_), .A2(new_n267_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n392_), .B1(new_n353_), .B2(new_n361_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n391_), .A2(new_n393_), .A3(KEYINPUT97), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT97), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n362_), .A2(new_n395_), .A3(new_n268_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n394_), .A2(KEYINPUT4), .A3(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G225gat), .A2(G233gat), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT4), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n393_), .A2(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n397_), .A2(new_n399_), .A3(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n394_), .A2(new_n398_), .A3(new_n396_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G1gat), .B(G29gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(KEYINPUT0), .ZN(new_n406_));
  INV_X1    g205(.A(G57gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(G85gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n408_), .B(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n404_), .A2(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n402_), .A2(new_n410_), .A3(new_n403_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n381_), .A2(new_n414_), .ZN(new_n415_));
  MUX2_X1   g214(.A(new_n318_), .B(new_n333_), .S(new_n319_), .Z(new_n416_));
  OAI211_X1 g215(.A(KEYINPUT27), .B(new_n326_), .C1(new_n416_), .C2(new_n325_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n337_), .A2(new_n415_), .A3(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n381_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n335_), .B1(new_n334_), .B2(new_n325_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n404_), .A2(KEYINPUT33), .A3(new_n411_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n397_), .A2(new_n401_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(new_n398_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n394_), .A2(new_n396_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(KEYINPUT99), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT99), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n394_), .A2(new_n426_), .A3(new_n396_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n425_), .A2(new_n399_), .A3(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n423_), .A2(new_n428_), .A3(new_n410_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n421_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT98), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n410_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n431_), .B1(new_n432_), .B2(KEYINPUT33), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT33), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n412_), .A2(KEYINPUT98), .A3(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n430_), .B1(new_n433_), .B2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n311_), .A2(new_n320_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n325_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n437_), .A2(KEYINPUT96), .A3(new_n438_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n420_), .A2(new_n436_), .A3(new_n439_), .A4(new_n326_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n325_), .A2(KEYINPUT32), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(KEYINPUT100), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n334_), .A2(new_n442_), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n443_), .B(new_n414_), .C1(new_n416_), .C2(new_n441_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n419_), .B1(new_n440_), .B2(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n418_), .B1(new_n445_), .B2(KEYINPUT101), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT101), .ZN(new_n447_));
  AOI211_X1 g246(.A(new_n447_), .B(new_n419_), .C1(new_n440_), .C2(new_n444_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n272_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT102), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT102), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n451_), .B(new_n272_), .C1(new_n446_), .C2(new_n448_), .ZN(new_n452_));
  AND2_X1   g251(.A1(new_n337_), .A2(new_n417_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n381_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n414_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n271_), .A2(new_n455_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n454_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n450_), .A2(new_n452_), .A3(new_n458_), .ZN(new_n459_));
  XOR2_X1   g258(.A(G29gat), .B(G36gat), .Z(new_n460_));
  XOR2_X1   g259(.A(G43gat), .B(G50gat), .Z(new_n461_));
  XNOR2_X1  g260(.A(new_n460_), .B(new_n461_), .ZN(new_n462_));
  XOR2_X1   g261(.A(new_n462_), .B(KEYINPUT80), .Z(new_n463_));
  XNOR2_X1  g262(.A(G15gat), .B(G22gat), .ZN(new_n464_));
  INV_X1    g263(.A(G1gat), .ZN(new_n465_));
  INV_X1    g264(.A(G8gat), .ZN(new_n466_));
  OAI21_X1  g265(.A(KEYINPUT14), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n464_), .A2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G1gat), .B(G8gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n468_), .B(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n463_), .B(new_n470_), .ZN(new_n471_));
  AND3_X1   g270(.A1(new_n471_), .A2(G229gat), .A3(G233gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G229gat), .A2(G233gat), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n463_), .A2(new_n470_), .ZN(new_n474_));
  XOR2_X1   g273(.A(new_n462_), .B(KEYINPUT76), .Z(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT15), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n474_), .B1(new_n476_), .B2(new_n470_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n472_), .B1(new_n473_), .B2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G113gat), .B(G141gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(G169gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(new_n288_), .ZN(new_n481_));
  AND2_X1   g280(.A1(new_n478_), .A2(new_n481_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n478_), .A2(new_n481_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n459_), .A2(new_n485_), .ZN(new_n486_));
  XOR2_X1   g285(.A(new_n486_), .B(KEYINPUT103), .Z(new_n487_));
  INV_X1    g286(.A(KEYINPUT37), .ZN(new_n488_));
  XOR2_X1   g287(.A(KEYINPUT70), .B(KEYINPUT6), .Z(new_n489_));
  NAND2_X1  g288(.A1(G99gat), .A2(G106gat), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  OR2_X1    g290(.A1(new_n489_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT7), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(KEYINPUT66), .ZN(new_n494_));
  NOR2_X1   g293(.A1(G99gat), .A2(G106gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n489_), .A2(new_n491_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n492_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  XOR2_X1   g297(.A(G85gat), .B(G92gat), .Z(new_n499_));
  AND2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT8), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  AND2_X1   g301(.A1(new_n501_), .A2(KEYINPUT68), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n501_), .A2(KEYINPUT68), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(new_n499_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(KEYINPUT65), .B(KEYINPUT6), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(new_n490_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n509_), .A2(KEYINPUT67), .A3(new_n496_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(KEYINPUT67), .B1(new_n509_), .B2(new_n496_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n507_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(KEYINPUT69), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n509_), .A2(new_n496_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT67), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(new_n510_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT69), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n518_), .A2(new_n519_), .A3(new_n507_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n502_), .B1(new_n514_), .B2(new_n520_), .ZN(new_n521_));
  XOR2_X1   g320(.A(KEYINPUT10), .B(G99gat), .Z(new_n522_));
  INV_X1    g321(.A(G106gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NOR3_X1   g323(.A1(new_n409_), .A2(new_n324_), .A3(KEYINPUT9), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n525_), .B1(new_n499_), .B2(KEYINPUT9), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n509_), .A2(new_n524_), .A3(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n521_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(new_n462_), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n527_), .B(KEYINPUT72), .Z(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n476_), .B1(new_n521_), .B2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G232gat), .A2(G233gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT75), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT34), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n536_), .A2(KEYINPUT35), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n530_), .A2(new_n533_), .A3(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n538_), .A2(KEYINPUT35), .A3(new_n536_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n536_), .A2(KEYINPUT35), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n530_), .A2(new_n533_), .A3(new_n540_), .A4(new_n537_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G190gat), .B(G218gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G134gat), .B(G162gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  XOR2_X1   g344(.A(new_n545_), .B(KEYINPUT36), .Z(new_n546_));
  NAND2_X1  g345(.A1(new_n542_), .A2(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n488_), .B1(new_n547_), .B2(KEYINPUT77), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n545_), .A2(KEYINPUT36), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n547_), .B1(new_n550_), .B2(new_n542_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n548_), .A2(new_n551_), .ZN(new_n552_));
  OAI221_X1 g351(.A(new_n547_), .B1(KEYINPUT77), .B2(new_n488_), .C1(new_n550_), .C2(new_n542_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  XOR2_X1   g354(.A(KEYINPUT74), .B(KEYINPUT13), .Z(new_n556_));
  NAND2_X1  g355(.A1(G230gat), .A2(G233gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT64), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n519_), .B1(new_n518_), .B2(new_n507_), .ZN(new_n560_));
  AOI211_X1 g359(.A(KEYINPUT69), .B(new_n506_), .C1(new_n517_), .C2(new_n510_), .ZN(new_n561_));
  OAI22_X1  g360(.A1(new_n560_), .A2(new_n561_), .B1(new_n501_), .B2(new_n500_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G57gat), .B(G64gat), .ZN(new_n563_));
  AND2_X1   g362(.A1(new_n563_), .A2(KEYINPUT11), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n563_), .A2(KEYINPUT11), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G71gat), .B(G78gat), .ZN(new_n566_));
  OR3_X1    g365(.A1(new_n564_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n563_), .A2(new_n566_), .A3(KEYINPUT11), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n569_), .B(KEYINPUT71), .Z(new_n570_));
  NAND3_X1  g369(.A1(new_n562_), .A2(new_n527_), .A3(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n570_), .B1(new_n562_), .B2(new_n527_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n559_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT12), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n569_), .A2(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n576_), .B1(new_n521_), .B2(new_n532_), .ZN(new_n577_));
  OAI211_X1 g376(.A(new_n577_), .B(new_n571_), .C1(new_n573_), .C2(KEYINPUT12), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n574_), .B1(new_n578_), .B2(new_n559_), .ZN(new_n579_));
  XOR2_X1   g378(.A(G120gat), .B(G148gat), .Z(new_n580_));
  XNOR2_X1  g379(.A(KEYINPUT73), .B(G204gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(KEYINPUT5), .B(G176gat), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n582_), .B(new_n583_), .Z(new_n584_));
  AND2_X1   g383(.A1(new_n579_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n584_), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n574_), .B(new_n586_), .C1(new_n578_), .C2(new_n559_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n556_), .B1(new_n585_), .B2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n579_), .A2(new_n584_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT13), .ZN(new_n591_));
  OAI211_X1 g390(.A(new_n590_), .B(new_n587_), .C1(KEYINPUT74), .C2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n589_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  AND2_X1   g393(.A1(G231gat), .A2(G233gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n470_), .B(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n570_), .B(new_n596_), .ZN(new_n597_));
  XOR2_X1   g396(.A(G183gat), .B(G211gat), .Z(new_n598_));
  XNOR2_X1  g397(.A(G127gat), .B(G155gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  XOR2_X1   g399(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n602_), .A2(KEYINPUT17), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n602_), .A2(KEYINPUT17), .ZN(new_n604_));
  OR3_X1    g403(.A1(new_n597_), .A2(new_n603_), .A3(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n596_), .ZN(new_n606_));
  AOI22_X1  g405(.A1(new_n603_), .A2(KEYINPUT79), .B1(new_n606_), .B2(new_n569_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n596_), .A2(new_n568_), .A3(new_n567_), .ZN(new_n608_));
  OAI211_X1 g407(.A(new_n607_), .B(new_n608_), .C1(KEYINPUT79), .C2(new_n603_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n605_), .A2(new_n609_), .ZN(new_n610_));
  NOR3_X1   g409(.A1(new_n555_), .A2(new_n594_), .A3(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n487_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n613_), .A2(new_n465_), .A3(new_n414_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT38), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n551_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n457_), .B1(new_n449_), .B2(KEYINPUT102), .ZN(new_n618_));
  AOI211_X1 g417(.A(new_n610_), .B(new_n617_), .C1(new_n618_), .C2(new_n452_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n594_), .A2(new_n484_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(G1gat), .B1(new_n621_), .B2(new_n455_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n614_), .A2(new_n615_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n616_), .A2(new_n622_), .A3(new_n623_), .ZN(G1324gat));
  OAI21_X1  g423(.A(G8gat), .B1(new_n621_), .B2(new_n453_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT39), .ZN(new_n626_));
  INV_X1    g425(.A(new_n453_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(new_n466_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n626_), .B1(new_n612_), .B2(new_n628_), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n629_), .B(KEYINPUT40), .Z(G1325gat));
  OR3_X1    g429(.A1(new_n612_), .A2(G15gat), .A3(new_n272_), .ZN(new_n631_));
  OAI21_X1  g430(.A(G15gat), .B1(new_n621_), .B2(new_n272_), .ZN(new_n632_));
  XOR2_X1   g431(.A(new_n632_), .B(KEYINPUT41), .Z(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n633_), .ZN(new_n634_));
  XOR2_X1   g433(.A(new_n634_), .B(KEYINPUT104), .Z(G1326gat));
  OAI21_X1  g434(.A(G22gat), .B1(new_n621_), .B2(new_n381_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT42), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n381_), .A2(G22gat), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n637_), .B1(new_n612_), .B2(new_n638_), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n639_), .B(KEYINPUT105), .Z(G1327gat));
  AOI211_X1 g439(.A(KEYINPUT43), .B(new_n554_), .C1(new_n618_), .C2(new_n452_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT43), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n642_), .B1(new_n459_), .B2(new_n555_), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n610_), .B(new_n620_), .C1(new_n641_), .C2(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(KEYINPUT44), .B1(new_n644_), .B2(KEYINPUT106), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n641_), .A2(new_n643_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT106), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n646_), .A2(new_n647_), .A3(new_n610_), .A4(new_n620_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n645_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT44), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n644_), .A2(new_n650_), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n649_), .A2(G29gat), .A3(new_n414_), .A4(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n610_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n551_), .A2(new_n653_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n654_), .A2(new_n593_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n487_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(new_n414_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n652_), .B1(new_n658_), .B2(G29gat), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT107), .ZN(G1328gat));
  NOR2_X1   g459(.A1(new_n453_), .A2(G36gat), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n487_), .A2(new_n655_), .A3(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT45), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n627_), .B1(new_n644_), .B2(new_n650_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n664_), .B1(new_n648_), .B2(new_n645_), .ZN(new_n665_));
  OAI21_X1  g464(.A(G36gat), .B1(new_n665_), .B2(KEYINPUT108), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT108), .ZN(new_n667_));
  AOI211_X1 g466(.A(new_n667_), .B(new_n664_), .C1(new_n648_), .C2(new_n645_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n663_), .B1(new_n666_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT46), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  OAI211_X1 g470(.A(new_n663_), .B(KEYINPUT46), .C1(new_n666_), .C2(new_n668_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1329gat));
  NAND4_X1  g472(.A1(new_n649_), .A2(G43gat), .A3(new_n271_), .A4(new_n651_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n656_), .A2(new_n271_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n674_), .B1(new_n676_), .B2(G43gat), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g477(.A(G50gat), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n419_), .A2(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT109), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n656_), .A2(new_n681_), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n649_), .A2(new_n419_), .A3(new_n651_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n682_), .B1(new_n683_), .B2(new_n679_), .ZN(G1331gat));
  NOR2_X1   g483(.A1(new_n593_), .A2(new_n485_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n619_), .A2(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(G57gat), .B1(new_n686_), .B2(new_n455_), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n459_), .A2(new_n653_), .A3(new_n554_), .A4(new_n685_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT110), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n414_), .A2(new_n407_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n687_), .B1(new_n690_), .B2(new_n691_), .ZN(G1332gat));
  OAI21_X1  g491(.A(G64gat), .B1(new_n686_), .B2(new_n453_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT48), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n453_), .A2(G64gat), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n694_), .B1(new_n690_), .B2(new_n695_), .ZN(G1333gat));
  OAI21_X1  g495(.A(G71gat), .B1(new_n686_), .B2(new_n272_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT49), .ZN(new_n698_));
  OR2_X1    g497(.A1(new_n272_), .A2(G71gat), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n698_), .B1(new_n690_), .B2(new_n699_), .ZN(G1334gat));
  OAI21_X1  g499(.A(G78gat), .B1(new_n686_), .B2(new_n381_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT50), .ZN(new_n702_));
  OR2_X1    g501(.A1(new_n381_), .A2(G78gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n702_), .B1(new_n690_), .B2(new_n703_), .ZN(G1335gat));
  NOR2_X1   g503(.A1(new_n641_), .A2(new_n643_), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n705_), .A2(KEYINPUT111), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(KEYINPUT111), .ZN(new_n707_));
  NOR3_X1   g506(.A1(new_n593_), .A2(new_n485_), .A3(new_n653_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n706_), .A2(new_n707_), .A3(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(G85gat), .B1(new_n709_), .B2(new_n455_), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n459_), .A2(new_n654_), .A3(new_n685_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n711_), .A2(new_n409_), .A3(new_n414_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT112), .ZN(G1336gat));
  NOR3_X1   g513(.A1(new_n709_), .A2(new_n324_), .A3(new_n453_), .ZN(new_n715_));
  AOI21_X1  g514(.A(G92gat), .B1(new_n711_), .B2(new_n627_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT113), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n715_), .A2(new_n717_), .ZN(G1337gat));
  INV_X1    g517(.A(KEYINPUT114), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n719_), .A2(KEYINPUT51), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n706_), .A2(new_n271_), .A3(new_n707_), .A4(new_n708_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(G99gat), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n711_), .A2(new_n271_), .A3(new_n522_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n720_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n719_), .A2(KEYINPUT51), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n724_), .B(new_n725_), .ZN(G1338gat));
  NAND3_X1  g525(.A1(new_n711_), .A2(new_n523_), .A3(new_n419_), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n646_), .A2(new_n419_), .A3(new_n610_), .A4(new_n685_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(G106gat), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n729_), .A2(KEYINPUT52), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n729_), .A2(KEYINPUT52), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n727_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g532(.A(KEYINPUT55), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n734_), .B1(new_n578_), .B2(new_n559_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n578_), .A2(new_n559_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n577_), .A2(new_n571_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n575_), .B1(new_n529_), .B2(new_n570_), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n737_), .A2(KEYINPUT55), .A3(new_n558_), .A4(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n735_), .A2(new_n736_), .A3(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(new_n584_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n588_), .B1(new_n741_), .B2(KEYINPUT56), .ZN(new_n742_));
  INV_X1    g541(.A(new_n477_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n473_), .B1(new_n743_), .B2(KEYINPUT116), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n744_), .B1(KEYINPUT116), .B2(new_n743_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n481_), .B1(new_n471_), .B2(new_n473_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n482_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT56), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n740_), .A2(new_n748_), .A3(new_n584_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n742_), .A2(new_n747_), .A3(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT58), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n742_), .A2(KEYINPUT58), .A3(new_n747_), .A4(new_n749_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n555_), .A2(new_n752_), .A3(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT57), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n741_), .A2(KEYINPUT56), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n756_), .A2(new_n485_), .A3(new_n587_), .A4(new_n749_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n747_), .B1(new_n585_), .B2(new_n588_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n755_), .B1(new_n759_), .B2(new_n551_), .ZN(new_n760_));
  AOI211_X1 g559(.A(KEYINPUT57), .B(new_n617_), .C1(new_n757_), .C2(new_n758_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n754_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT117), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n754_), .B(KEYINPUT117), .C1(new_n760_), .C2(new_n761_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n764_), .A2(new_n610_), .A3(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n484_), .A2(new_n653_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n767_), .B1(new_n589_), .B2(new_n592_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n554_), .B1(new_n768_), .B2(KEYINPUT115), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(KEYINPUT115), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(KEYINPUT54), .B1(new_n769_), .B2(new_n771_), .ZN(new_n772_));
  OR2_X1    g571(.A1(new_n768_), .A2(KEYINPUT115), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT54), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n773_), .A2(new_n774_), .A3(new_n554_), .A4(new_n770_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n772_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n766_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT118), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NOR3_X1   g579(.A1(new_n454_), .A2(new_n272_), .A3(new_n455_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n766_), .A2(KEYINPUT118), .A3(new_n777_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n780_), .A2(new_n781_), .A3(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n784_), .A2(new_n263_), .A3(new_n485_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n776_), .B1(new_n610_), .B2(new_n762_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT59), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n781_), .A2(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(KEYINPUT119), .B1(new_n786_), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT119), .ZN(new_n790_));
  INV_X1    g589(.A(new_n788_), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n762_), .A2(new_n610_), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n790_), .B(new_n791_), .C1(new_n792_), .C2(new_n776_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n789_), .A2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n794_), .B1(new_n783_), .B2(KEYINPUT59), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n795_), .A2(new_n485_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n785_), .B1(new_n796_), .B2(new_n263_), .ZN(G1340gat));
  AOI21_X1  g596(.A(new_n261_), .B1(new_n795_), .B2(new_n594_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n261_), .B1(new_n593_), .B2(KEYINPUT60), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n799_), .B1(KEYINPUT60), .B2(new_n261_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n783_), .A2(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(KEYINPUT120), .B1(new_n798_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT120), .ZN(new_n803_));
  INV_X1    g602(.A(new_n801_), .ZN(new_n804_));
  AOI211_X1 g603(.A(new_n593_), .B(new_n794_), .C1(new_n783_), .C2(KEYINPUT59), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n803_), .B(new_n804_), .C1(new_n805_), .C2(new_n261_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n802_), .A2(new_n806_), .ZN(G1341gat));
  NAND3_X1  g606(.A1(new_n784_), .A2(new_n258_), .A3(new_n653_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n795_), .A2(new_n653_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n808_), .B1(new_n809_), .B2(new_n258_), .ZN(G1342gat));
  NAND3_X1  g609(.A1(new_n784_), .A2(new_n256_), .A3(new_n617_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n795_), .A2(new_n555_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n811_), .B1(new_n812_), .B2(new_n256_), .ZN(G1343gat));
  AND2_X1   g612(.A1(new_n780_), .A2(new_n782_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n271_), .A2(new_n381_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n627_), .A2(new_n455_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n814_), .A2(new_n815_), .A3(new_n816_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n817_), .A2(new_n484_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(KEYINPUT121), .B(G141gat), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n818_), .B(new_n819_), .ZN(G1344gat));
  NOR2_X1   g619(.A1(new_n817_), .A2(new_n593_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(new_n356_), .ZN(G1345gat));
  NOR2_X1   g621(.A1(new_n817_), .A2(new_n610_), .ZN(new_n823_));
  XOR2_X1   g622(.A(KEYINPUT61), .B(G155gat), .Z(new_n824_));
  XNOR2_X1  g623(.A(new_n823_), .B(new_n824_), .ZN(G1346gat));
  OAI21_X1  g624(.A(G162gat), .B1(new_n817_), .B2(new_n554_), .ZN(new_n826_));
  OR2_X1    g625(.A1(new_n551_), .A2(G162gat), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n826_), .B1(new_n817_), .B2(new_n827_), .ZN(G1347gat));
  NOR2_X1   g627(.A1(new_n456_), .A2(new_n453_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  NOR3_X1   g629(.A1(new_n786_), .A2(new_n419_), .A3(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n220_), .B1(new_n831_), .B2(new_n485_), .ZN(new_n832_));
  XOR2_X1   g631(.A(KEYINPUT122), .B(KEYINPUT62), .Z(new_n833_));
  OR2_X1    g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n831_), .A2(new_n485_), .A3(new_n232_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n832_), .A2(new_n833_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n834_), .A2(new_n835_), .A3(new_n836_), .ZN(G1348gat));
  AOI21_X1  g636(.A(G176gat), .B1(new_n831_), .B2(new_n594_), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n814_), .A2(new_n381_), .ZN(new_n839_));
  NOR3_X1   g638(.A1(new_n830_), .A2(new_n224_), .A3(new_n593_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n838_), .B1(new_n839_), .B2(new_n840_), .ZN(G1349gat));
  NAND3_X1  g640(.A1(new_n839_), .A2(new_n653_), .A3(new_n829_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n610_), .A2(new_n240_), .ZN(new_n843_));
  AOI22_X1  g642(.A1(new_n842_), .A2(new_n207_), .B1(new_n831_), .B2(new_n843_), .ZN(G1350gat));
  AOI21_X1  g643(.A(new_n208_), .B1(new_n831_), .B2(new_n555_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(KEYINPUT123), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n831_), .A2(new_n241_), .A3(new_n617_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(G1351gat));
  NOR2_X1   g647(.A1(new_n453_), .A2(new_n414_), .ZN(new_n849_));
  AND3_X1   g648(.A1(new_n814_), .A2(new_n815_), .A3(new_n849_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n850_), .A2(KEYINPUT124), .A3(G197gat), .A4(new_n485_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT124), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n814_), .A2(new_n485_), .A3(new_n815_), .A4(new_n849_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n853_), .B2(new_n288_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n288_), .ZN(new_n855_));
  AND3_X1   g654(.A1(new_n851_), .A2(new_n854_), .A3(new_n855_), .ZN(G1352gat));
  NAND4_X1  g655(.A1(new_n814_), .A2(new_n594_), .A3(new_n815_), .A4(new_n849_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT125), .ZN(new_n858_));
  OR3_X1    g657(.A1(new_n857_), .A2(new_n858_), .A3(new_n293_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(G204gat), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n858_), .B1(new_n857_), .B2(new_n293_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n859_), .A2(new_n860_), .A3(new_n861_), .ZN(G1353gat));
  XOR2_X1   g661(.A(KEYINPUT63), .B(G211gat), .Z(new_n863_));
  NAND3_X1  g662(.A1(new_n850_), .A2(new_n653_), .A3(new_n863_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n814_), .A2(new_n815_), .A3(new_n849_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(new_n866_), .B2(new_n610_), .ZN(new_n867_));
  AND2_X1   g666(.A1(new_n864_), .A2(new_n867_), .ZN(G1354gat));
  XOR2_X1   g667(.A(KEYINPUT126), .B(G218gat), .Z(new_n869_));
  NOR3_X1   g668(.A1(new_n866_), .A2(new_n554_), .A3(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n850_), .A2(new_n617_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n870_), .B1(new_n871_), .B2(new_n869_), .ZN(G1355gat));
endmodule


