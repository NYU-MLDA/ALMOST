//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1 0 0 1 1 0 1 0 1 0 1 0 0 1 1 1 1 0 0 0 1 0 0 1 1 0 1 0 0 0 0 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 0 0 1 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n589_, new_n590_, new_n591_, new_n592_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n673_, new_n674_,
    new_n675_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n825_, new_n826_, new_n827_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n873_, new_n874_, new_n875_, new_n876_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n883_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_;
  NAND2_X1  g000(.A1(G232gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT34), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(KEYINPUT70), .B(KEYINPUT35), .Z(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT73), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n207_), .B1(new_n204_), .B2(new_n205_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G99gat), .A2(G106gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT6), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT7), .ZN(new_n211_));
  INV_X1    g010(.A(G99gat), .ZN(new_n212_));
  INV_X1    g011(.A(G106gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n210_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT8), .ZN(new_n217_));
  XOR2_X1   g016(.A(G85gat), .B(G92gat), .Z(new_n218_));
  NAND3_X1  g017(.A1(new_n216_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n220_));
  INV_X1    g019(.A(new_n215_), .ZN(new_n221_));
  NOR3_X1   g020(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n220_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n214_), .A2(KEYINPUT65), .A3(new_n215_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n223_), .A2(new_n210_), .A3(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n225_), .A2(KEYINPUT66), .A3(new_n218_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT8), .ZN(new_n227_));
  AOI21_X1  g026(.A(KEYINPUT66), .B1(new_n225_), .B2(new_n218_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n219_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n218_), .A2(KEYINPUT9), .ZN(new_n230_));
  XOR2_X1   g029(.A(KEYINPUT10), .B(G99gat), .Z(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(new_n213_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT64), .B(G92gat), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT9), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n233_), .A2(new_n234_), .A3(G85gat), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n230_), .A2(new_n232_), .A3(new_n210_), .A4(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n229_), .A2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G29gat), .B(G36gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT71), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G43gat), .B(G50gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n208_), .B1(new_n237_), .B2(new_n241_), .ZN(new_n242_));
  AND2_X1   g041(.A1(new_n239_), .A2(new_n240_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n239_), .A2(new_n240_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  XOR2_X1   g044(.A(KEYINPUT72), .B(KEYINPUT15), .Z(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n246_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n241_), .A2(new_n248_), .ZN(new_n249_));
  AOI22_X1  g048(.A1(new_n247_), .A2(new_n249_), .B1(new_n229_), .B2(new_n236_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n206_), .B1(new_n242_), .B2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n247_), .A2(new_n249_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(new_n237_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n236_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n225_), .A2(new_n218_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT66), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n257_), .A2(KEYINPUT8), .A3(new_n226_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n254_), .B1(new_n258_), .B2(new_n219_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(new_n245_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n206_), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n253_), .A2(new_n260_), .A3(new_n261_), .A4(new_n208_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n251_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT75), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G190gat), .B(G218gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G134gat), .B(G162gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  XOR2_X1   g066(.A(new_n267_), .B(KEYINPUT36), .Z(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT74), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n263_), .A2(new_n264_), .A3(new_n269_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n267_), .A2(KEYINPUT36), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n251_), .A2(new_n262_), .A3(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n264_), .B1(new_n263_), .B2(new_n269_), .ZN(new_n274_));
  OAI21_X1  g073(.A(KEYINPUT37), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT76), .ZN(new_n276_));
  AND3_X1   g075(.A1(new_n251_), .A2(new_n262_), .A3(new_n271_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n268_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n278_), .B1(new_n251_), .B2(new_n262_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT37), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n276_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n275_), .A2(new_n282_), .ZN(new_n283_));
  OAI211_X1 g082(.A(new_n276_), .B(KEYINPUT37), .C1(new_n273_), .C2(new_n274_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G71gat), .B(G78gat), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT67), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G57gat), .B(G64gat), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n286_), .B(new_n287_), .C1(KEYINPUT11), .C2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(G64gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(G57gat), .ZN(new_n291_));
  INV_X1    g090(.A(G57gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(G64gat), .ZN(new_n293_));
  AOI21_X1  g092(.A(KEYINPUT11), .B1(new_n291_), .B2(new_n293_), .ZN(new_n294_));
  OAI21_X1  g093(.A(KEYINPUT67), .B1(new_n294_), .B2(new_n285_), .ZN(new_n295_));
  AND2_X1   g094(.A1(new_n288_), .A2(KEYINPUT11), .ZN(new_n296_));
  AND3_X1   g095(.A1(new_n289_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n296_), .B1(new_n289_), .B2(new_n295_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G231gat), .A2(G233gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G1gat), .B(G8gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT77), .ZN(new_n303_));
  INV_X1    g102(.A(G15gat), .ZN(new_n304_));
  INV_X1    g103(.A(G22gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G15gat), .A2(G22gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G1gat), .A2(G8gat), .ZN(new_n308_));
  AOI22_X1  g107(.A1(new_n306_), .A2(new_n307_), .B1(KEYINPUT14), .B2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n303_), .B(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n301_), .B(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(G183gat), .B(G211gat), .Z(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT79), .ZN(new_n314_));
  XOR2_X1   g113(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G127gat), .B(G155gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT17), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  AND2_X1   g119(.A1(new_n318_), .A2(new_n319_), .ZN(new_n321_));
  OR3_X1    g120(.A1(new_n312_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n312_), .A2(new_n320_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n283_), .A2(new_n284_), .A3(new_n325_), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n326_), .B(KEYINPUT80), .Z(new_n327_));
  XNOR2_X1  g126(.A(G120gat), .B(G148gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT5), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G176gat), .B(G204gat), .ZN(new_n330_));
  XOR2_X1   g129(.A(new_n329_), .B(new_n330_), .Z(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n299_), .ZN(new_n333_));
  OAI21_X1  g132(.A(KEYINPUT68), .B1(new_n237_), .B2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n237_), .A2(new_n333_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT68), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n259_), .A2(new_n336_), .A3(new_n299_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n334_), .A2(new_n335_), .A3(new_n337_), .ZN(new_n338_));
  AND2_X1   g137(.A1(G230gat), .A2(G233gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n339_), .B1(new_n259_), .B2(new_n299_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT12), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n342_), .B1(new_n237_), .B2(new_n333_), .ZN(new_n343_));
  AOI211_X1 g142(.A(KEYINPUT12), .B(new_n299_), .C1(new_n229_), .C2(new_n236_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n341_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n332_), .B1(new_n340_), .B2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n340_), .A2(new_n345_), .A3(new_n332_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT69), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT13), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n347_), .A2(new_n348_), .A3(new_n350_), .ZN(new_n351_));
  XOR2_X1   g150(.A(KEYINPUT69), .B(KEYINPUT13), .Z(new_n352_));
  AND3_X1   g151(.A1(new_n340_), .A2(new_n345_), .A3(new_n332_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n352_), .B1(new_n353_), .B2(new_n346_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n351_), .A2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n327_), .A2(KEYINPUT81), .A3(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n252_), .A2(new_n310_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n311_), .A2(new_n245_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G229gat), .A2(G233gat), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n357_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n241_), .A2(new_n310_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n358_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n359_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n360_), .A2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G113gat), .B(G141gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT82), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G169gat), .B(G197gat), .ZN(new_n368_));
  XOR2_X1   g167(.A(new_n367_), .B(new_n368_), .Z(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n365_), .B(new_n370_), .ZN(new_n371_));
  XOR2_X1   g170(.A(G197gat), .B(G204gat), .Z(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(KEYINPUT21), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G211gat), .B(G218gat), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(KEYINPUT91), .ZN(new_n376_));
  OR2_X1    g175(.A1(new_n372_), .A2(KEYINPUT21), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n377_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(G169gat), .ZN(new_n382_));
  INV_X1    g181(.A(G176gat), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n381_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT83), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n381_), .B(KEYINPUT83), .C1(new_n382_), .C2(new_n383_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT25), .B(G183gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT26), .B(G190gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NOR3_X1   g189(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G183gat), .A2(G190gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(KEYINPUT23), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT23), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n394_), .A2(G183gat), .A3(G190gat), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n391_), .B1(new_n393_), .B2(new_n395_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n386_), .A2(new_n387_), .A3(new_n390_), .A4(new_n396_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(G183gat), .A2(G190gat), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n398_), .B1(new_n394_), .B2(new_n392_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n399_), .B1(new_n394_), .B2(new_n392_), .ZN(new_n400_));
  OAI21_X1  g199(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n401_));
  OR3_X1    g200(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n400_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n397_), .A2(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(KEYINPUT20), .B1(new_n379_), .B2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT92), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  AND2_X1   g206(.A1(new_n390_), .A2(new_n384_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT93), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n396_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n403_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n379_), .A2(new_n412_), .ZN(new_n413_));
  OAI211_X1 g212(.A(KEYINPUT92), .B(KEYINPUT20), .C1(new_n379_), .C2(new_n404_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n407_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G226gat), .A2(G233gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT19), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n415_), .A2(new_n417_), .ZN(new_n418_));
  OR2_X1    g217(.A1(new_n379_), .A2(new_n412_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n417_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n379_), .A2(new_n404_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n419_), .A2(KEYINPUT20), .A3(new_n420_), .A4(new_n421_), .ZN(new_n422_));
  XOR2_X1   g221(.A(G8gat), .B(G36gat), .Z(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G64gat), .B(G92gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n425_), .B(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT32), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n418_), .A2(new_n422_), .A3(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n415_), .A2(new_n417_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n419_), .A2(KEYINPUT20), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT97), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n419_), .A2(KEYINPUT97), .A3(KEYINPUT20), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n433_), .A2(new_n421_), .A3(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n430_), .B1(new_n417_), .B2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n429_), .B1(new_n436_), .B2(new_n428_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G225gat), .A2(G233gat), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT4), .ZN(new_n440_));
  XOR2_X1   g239(.A(G155gat), .B(G162gat), .Z(new_n441_));
  AOI21_X1  g240(.A(KEYINPUT89), .B1(G141gat), .B2(G148gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(KEYINPUT2), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT88), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n444_), .B(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n443_), .A2(new_n446_), .ZN(new_n447_));
  NOR3_X1   g246(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n448_));
  XOR2_X1   g247(.A(new_n448_), .B(KEYINPUT87), .Z(new_n449_));
  OAI21_X1  g248(.A(new_n441_), .B1(new_n447_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT95), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT1), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n441_), .A2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n454_));
  INV_X1    g253(.A(G141gat), .ZN(new_n455_));
  INV_X1    g254(.A(G148gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G141gat), .A2(G148gat), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n453_), .A2(new_n454_), .A3(new_n457_), .A4(new_n458_), .ZN(new_n459_));
  AND3_X1   g258(.A1(new_n450_), .A2(new_n451_), .A3(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G127gat), .B(G134gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G113gat), .B(G120gat), .ZN(new_n462_));
  XOR2_X1   g261(.A(new_n461_), .B(new_n462_), .Z(new_n463_));
  OR2_X1    g262(.A1(new_n460_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n460_), .A2(new_n463_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n440_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  AND2_X1   g265(.A1(new_n450_), .A2(new_n459_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n463_), .ZN(new_n468_));
  NOR3_X1   g267(.A1(new_n467_), .A2(KEYINPUT4), .A3(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n439_), .B1(new_n466_), .B2(new_n469_), .ZN(new_n470_));
  AND2_X1   g269(.A1(new_n464_), .A2(new_n465_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(new_n438_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G1gat), .B(G29gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(G85gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT0), .B(G57gat), .ZN(new_n476_));
  XOR2_X1   g275(.A(new_n475_), .B(new_n476_), .Z(new_n477_));
  NAND2_X1  g276(.A1(new_n473_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n477_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n470_), .A2(new_n472_), .A3(new_n479_), .ZN(new_n480_));
  AND2_X1   g279(.A1(new_n478_), .A2(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(KEYINPUT98), .B1(new_n437_), .B2(new_n481_), .ZN(new_n482_));
  AOI22_X1  g281(.A1(new_n431_), .A2(new_n432_), .B1(new_n379_), .B2(new_n404_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n420_), .B1(new_n483_), .B2(new_n434_), .ZN(new_n484_));
  OAI211_X1 g283(.A(KEYINPUT32), .B(new_n427_), .C1(new_n484_), .C2(new_n430_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n478_), .A2(new_n480_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT98), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n485_), .A2(new_n486_), .A3(new_n487_), .A4(new_n429_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n418_), .A2(new_n427_), .A3(new_n422_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n427_), .B1(new_n418_), .B2(new_n422_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT33), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n478_), .A2(KEYINPUT96), .A3(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(KEYINPUT96), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n473_), .A2(new_n477_), .A3(new_n495_), .ZN(new_n496_));
  OR3_X1    g295(.A1(new_n466_), .A2(new_n439_), .A3(new_n469_), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n497_), .B(new_n479_), .C1(new_n438_), .C2(new_n471_), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n492_), .A2(new_n494_), .A3(new_n496_), .A4(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n482_), .A2(new_n488_), .A3(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G71gat), .B(G99gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(G43gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n404_), .B(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT84), .B(KEYINPUT31), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(KEYINPUT85), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n503_), .B(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G227gat), .A2(G233gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(new_n304_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT30), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(new_n463_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n506_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n506_), .A2(new_n510_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT86), .ZN(new_n514_));
  NOR3_X1   g313(.A1(new_n512_), .A2(new_n513_), .A3(new_n514_), .ZN(new_n515_));
  OR2_X1    g314(.A1(new_n506_), .A2(new_n510_), .ZN(new_n516_));
  AOI21_X1  g315(.A(KEYINPUT86), .B1(new_n516_), .B2(new_n511_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G22gat), .B(G50gat), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT29), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n379_), .B1(new_n521_), .B2(new_n467_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(G78gat), .ZN(new_n523_));
  INV_X1    g322(.A(G78gat), .ZN(new_n524_));
  OAI211_X1 g323(.A(new_n379_), .B(new_n524_), .C1(new_n521_), .C2(new_n467_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n523_), .A2(G106gat), .A3(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(G106gat), .B1(new_n523_), .B2(new_n525_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n520_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n528_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n520_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n530_), .A2(new_n526_), .A3(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n467_), .A2(new_n521_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT28), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G228gat), .A2(G233gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT90), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n534_), .B(new_n536_), .ZN(new_n537_));
  AND3_X1   g336(.A1(new_n529_), .A2(new_n532_), .A3(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n537_), .B1(new_n529_), .B2(new_n532_), .ZN(new_n539_));
  NOR3_X1   g338(.A1(new_n519_), .A2(new_n538_), .A3(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n500_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n489_), .A2(KEYINPUT100), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT100), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n418_), .A2(new_n543_), .A3(new_n427_), .A4(new_n422_), .ZN(new_n544_));
  OAI211_X1 g343(.A(new_n542_), .B(new_n544_), .C1(new_n436_), .C2(new_n427_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(KEYINPUT27), .ZN(new_n546_));
  OR3_X1    g345(.A1(new_n490_), .A2(new_n491_), .A3(KEYINPUT27), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n486_), .B(KEYINPUT99), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n518_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n529_), .A2(new_n532_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n537_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n529_), .A2(new_n532_), .A3(new_n537_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n512_), .A2(new_n513_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n553_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n550_), .A2(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n548_), .A2(new_n549_), .A3(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n371_), .B1(new_n541_), .B2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n356_), .A2(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(KEYINPUT81), .B1(new_n327_), .B2(new_n355_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  OR2_X1    g361(.A1(new_n562_), .A2(KEYINPUT101), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(KEYINPUT101), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n549_), .A2(G1gat), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n563_), .A2(new_n564_), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT38), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n563_), .A2(KEYINPUT38), .A3(new_n564_), .A4(new_n565_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n280_), .B1(new_n541_), .B2(new_n558_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n365_), .B(new_n369_), .ZN(new_n571_));
  AND4_X1   g370(.A1(new_n325_), .A2(new_n570_), .A3(new_n355_), .A4(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n549_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(G1gat), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n575_), .B(KEYINPUT102), .Z(new_n576_));
  NAND3_X1  g375(.A1(new_n568_), .A2(new_n569_), .A3(new_n576_), .ZN(G1324gat));
  NOR2_X1   g376(.A1(new_n548_), .A2(G8gat), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n563_), .A2(new_n564_), .A3(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n548_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n572_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(G8gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT39), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n579_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT40), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n579_), .A2(new_n583_), .A3(KEYINPUT40), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(G1325gat));
  AOI21_X1  g387(.A(new_n304_), .B1(new_n572_), .B2(new_n519_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT41), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n563_), .A2(new_n564_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n519_), .A2(new_n304_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n590_), .B1(new_n591_), .B2(new_n592_), .ZN(G1326gat));
  NOR2_X1   g392(.A1(new_n538_), .A2(new_n539_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(new_n305_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT103), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n563_), .A2(new_n564_), .A3(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n305_), .B1(new_n572_), .B2(new_n595_), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n599_), .B(KEYINPUT42), .Z(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(KEYINPUT104), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT104), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n598_), .A2(new_n600_), .A3(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(G1327gat));
  INV_X1    g404(.A(new_n280_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n325_), .A2(new_n606_), .ZN(new_n607_));
  AND3_X1   g406(.A1(new_n559_), .A2(new_n355_), .A3(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(G29gat), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n608_), .A2(new_n609_), .A3(new_n573_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n355_), .ZN(new_n611_));
  NOR3_X1   g410(.A1(new_n611_), .A2(new_n325_), .A3(new_n371_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n541_), .A2(new_n558_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT43), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n283_), .A2(new_n284_), .ZN(new_n615_));
  AND3_X1   g414(.A1(new_n613_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n614_), .B1(new_n613_), .B2(new_n615_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n612_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT44), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  OAI211_X1 g419(.A(KEYINPUT44), .B(new_n612_), .C1(new_n616_), .C2(new_n617_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n620_), .A2(new_n573_), .A3(new_n621_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n622_), .A2(KEYINPUT105), .ZN(new_n623_));
  OAI21_X1  g422(.A(G29gat), .B1(new_n622_), .B2(KEYINPUT105), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n610_), .B1(new_n623_), .B2(new_n624_), .ZN(G1328gat));
  INV_X1    g424(.A(G36gat), .ZN(new_n626_));
  OR2_X1    g425(.A1(new_n548_), .A2(KEYINPUT106), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n548_), .A2(KEYINPUT106), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n608_), .A2(new_n626_), .A3(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT45), .ZN(new_n631_));
  AND3_X1   g430(.A1(new_n620_), .A2(new_n580_), .A3(new_n621_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n631_), .B1(new_n632_), .B2(new_n626_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT46), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(G1329gat));
  AND2_X1   g434(.A1(new_n555_), .A2(G43gat), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n620_), .A2(new_n621_), .A3(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(KEYINPUT107), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT107), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n620_), .A2(new_n639_), .A3(new_n621_), .A4(new_n636_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n638_), .A2(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(G43gat), .B1(new_n608_), .B2(new_n519_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT108), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(KEYINPUT47), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT47), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n641_), .A2(new_n646_), .A3(new_n643_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(G1330gat));
  INV_X1    g447(.A(G50gat), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n608_), .A2(new_n649_), .A3(new_n595_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n620_), .A2(new_n595_), .A3(new_n621_), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n651_), .A2(KEYINPUT109), .A3(G50gat), .ZN(new_n652_));
  AOI21_X1  g451(.A(KEYINPUT109), .B1(new_n651_), .B2(G50gat), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n650_), .B1(new_n652_), .B2(new_n653_), .ZN(G1331gat));
  NOR2_X1   g453(.A1(new_n355_), .A2(new_n571_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n656_), .B1(new_n541_), .B2(new_n558_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n327_), .A2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n658_), .A2(new_n292_), .A3(new_n573_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n570_), .A2(new_n325_), .A3(new_n655_), .ZN(new_n660_));
  OAI21_X1  g459(.A(G57gat), .B1(new_n660_), .B2(new_n549_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n659_), .A2(new_n661_), .ZN(G1332gat));
  INV_X1    g461(.A(new_n629_), .ZN(new_n663_));
  OAI21_X1  g462(.A(G64gat), .B1(new_n660_), .B2(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT48), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n658_), .A2(new_n290_), .A3(new_n629_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(G1333gat));
  OAI21_X1  g466(.A(G71gat), .B1(new_n660_), .B2(new_n518_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT49), .ZN(new_n669_));
  INV_X1    g468(.A(G71gat), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n658_), .A2(new_n670_), .A3(new_n519_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(G1334gat));
  OAI21_X1  g471(.A(G78gat), .B1(new_n660_), .B2(new_n594_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT50), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n658_), .A2(new_n524_), .A3(new_n595_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(G1335gat));
  NAND2_X1  g475(.A1(new_n657_), .A2(new_n607_), .ZN(new_n677_));
  XOR2_X1   g476(.A(new_n677_), .B(KEYINPUT110), .Z(new_n678_));
  AOI21_X1  g477(.A(G85gat), .B1(new_n678_), .B2(new_n573_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT111), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n616_), .A2(new_n617_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n656_), .A2(new_n325_), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n573_), .A2(G85gat), .ZN(new_n684_));
  XOR2_X1   g483(.A(new_n684_), .B(KEYINPUT112), .Z(new_n685_));
  AOI21_X1  g484(.A(new_n680_), .B1(new_n683_), .B2(new_n685_), .ZN(G1336gat));
  AOI21_X1  g485(.A(G92gat), .B1(new_n678_), .B2(new_n580_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n629_), .A2(new_n233_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(new_n683_), .B2(new_n688_), .ZN(G1337gat));
  NAND2_X1  g488(.A1(new_n683_), .A2(new_n519_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(G99gat), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT113), .ZN(new_n692_));
  OR2_X1    g491(.A1(new_n692_), .A2(KEYINPUT51), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n555_), .A2(new_n231_), .ZN(new_n694_));
  AOI22_X1  g493(.A1(new_n678_), .A2(new_n694_), .B1(new_n692_), .B2(KEYINPUT51), .ZN(new_n695_));
  AND3_X1   g494(.A1(new_n691_), .A2(new_n693_), .A3(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n693_), .B1(new_n691_), .B2(new_n695_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n696_), .A2(new_n697_), .ZN(G1338gat));
  NAND3_X1  g497(.A1(new_n678_), .A2(new_n213_), .A3(new_n595_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n681_), .A2(new_n595_), .A3(new_n682_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT52), .ZN(new_n701_));
  AND3_X1   g500(.A1(new_n700_), .A2(new_n701_), .A3(G106gat), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n701_), .B1(new_n700_), .B2(G106gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n699_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(KEYINPUT53), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT53), .ZN(new_n706_));
  OAI211_X1 g505(.A(new_n706_), .B(new_n699_), .C1(new_n702_), .C2(new_n703_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n707_), .ZN(G1339gat));
  INV_X1    g507(.A(new_n556_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n573_), .A2(new_n548_), .A3(new_n709_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n371_), .A2(new_n353_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n343_), .A2(new_n344_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n334_), .A2(new_n337_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n339_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT55), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n345_), .A2(new_n715_), .ZN(new_n716_));
  OAI211_X1 g515(.A(KEYINPUT55), .B(new_n341_), .C1(new_n343_), .C2(new_n344_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n714_), .A2(new_n716_), .A3(new_n717_), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n718_), .A2(KEYINPUT56), .A3(new_n331_), .ZN(new_n719_));
  AOI21_X1  g518(.A(KEYINPUT56), .B1(new_n718_), .B2(new_n331_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n711_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(KEYINPUT114), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT114), .ZN(new_n723_));
  OAI211_X1 g522(.A(new_n723_), .B(new_n711_), .C1(new_n719_), .C2(new_n720_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n365_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n357_), .A2(new_n358_), .A3(new_n363_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n370_), .B1(new_n362_), .B2(new_n359_), .ZN(new_n727_));
  AOI22_X1  g526(.A1(new_n725_), .A2(new_n370_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n728_), .B1(new_n353_), .B2(new_n346_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT115), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  OAI211_X1 g530(.A(new_n728_), .B(KEYINPUT115), .C1(new_n353_), .C2(new_n346_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n722_), .A2(new_n724_), .A3(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(new_n606_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT57), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n280_), .A2(new_n736_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT58), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n728_), .A2(new_n348_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n740_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n741_));
  AOI22_X1  g540(.A1(new_n739_), .A2(new_n741_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n741_), .A2(new_n739_), .ZN(new_n743_));
  AOI22_X1  g542(.A1(new_n734_), .A2(new_n738_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n325_), .B1(new_n737_), .B2(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n571_), .B1(new_n351_), .B2(new_n354_), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n283_), .A2(new_n746_), .A3(new_n284_), .A4(new_n325_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT54), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n747_), .B(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(KEYINPUT116), .B1(new_n745_), .B2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n571_), .A2(new_n348_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n718_), .A2(new_n331_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT56), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n718_), .A2(KEYINPUT56), .A3(new_n331_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n751_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n733_), .B1(new_n756_), .B2(new_n723_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n724_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n738_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n742_), .A2(new_n743_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(KEYINPUT57), .B1(new_n734_), .B2(new_n606_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n324_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT116), .ZN(new_n764_));
  INV_X1    g563(.A(new_n749_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n763_), .A2(new_n764_), .A3(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n710_), .B1(new_n750_), .B2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(G113gat), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n767_), .A2(new_n768_), .A3(new_n571_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n763_), .A2(new_n765_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n710_), .A2(KEYINPUT59), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n770_), .A2(KEYINPUT117), .A3(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT117), .ZN(new_n773_));
  AOI22_X1  g572(.A1(new_n721_), .A2(KEYINPUT114), .B1(new_n731_), .B2(new_n732_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n280_), .B1(new_n774_), .B2(new_n724_), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n759_), .B(new_n760_), .C1(new_n775_), .C2(KEYINPUT57), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n749_), .B1(new_n776_), .B2(new_n324_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n771_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n773_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n772_), .A2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT59), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n780_), .B(new_n571_), .C1(new_n767_), .C2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n769_), .B1(new_n783_), .B2(new_n768_), .ZN(G1340gat));
  NAND2_X1  g583(.A1(new_n780_), .A2(new_n611_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n750_), .A2(new_n766_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n710_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n781_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(KEYINPUT118), .B1(new_n785_), .B2(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n355_), .B1(new_n772_), .B2(new_n779_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT118), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n790_), .B(new_n791_), .C1(new_n781_), .C2(new_n767_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n789_), .A2(G120gat), .A3(new_n792_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n355_), .A2(KEYINPUT60), .ZN(new_n794_));
  MUX2_X1   g593(.A(new_n794_), .B(KEYINPUT60), .S(G120gat), .Z(new_n795_));
  NAND2_X1  g594(.A1(new_n767_), .A2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n793_), .A2(new_n796_), .ZN(G1341gat));
  NAND2_X1  g596(.A1(new_n767_), .A2(new_n325_), .ZN(new_n798_));
  INV_X1    g597(.A(G127gat), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n324_), .A2(new_n799_), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n780_), .B(new_n801_), .C1(new_n767_), .C2(new_n781_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT119), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n800_), .A2(new_n802_), .A3(KEYINPUT119), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(G1342gat));
  NAND2_X1  g606(.A1(new_n767_), .A2(new_n280_), .ZN(new_n808_));
  INV_X1    g607(.A(G134gat), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n809_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n780_), .B(new_n811_), .C1(new_n767_), .C2(new_n781_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT120), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT120), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n810_), .A2(new_n812_), .A3(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n814_), .A2(new_n816_), .ZN(G1343gat));
  NOR3_X1   g616(.A1(new_n629_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n818_));
  AND3_X1   g617(.A1(new_n786_), .A2(KEYINPUT121), .A3(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(KEYINPUT121), .B1(new_n786_), .B2(new_n818_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n571_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(G141gat), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n455_), .B(new_n571_), .C1(new_n819_), .C2(new_n820_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(G1344gat));
  OAI21_X1  g623(.A(new_n611_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(G148gat), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n456_), .B(new_n611_), .C1(new_n819_), .C2(new_n820_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(G1345gat));
  OAI21_X1  g627(.A(new_n325_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(KEYINPUT61), .B(G155gat), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n830_), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n325_), .B(new_n832_), .C1(new_n819_), .C2(new_n820_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(G1346gat));
  OR2_X1    g633(.A1(new_n819_), .A2(new_n820_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n615_), .A2(G162gat), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n836_), .B(KEYINPUT122), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n280_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n838_));
  INV_X1    g637(.A(G162gat), .ZN(new_n839_));
  AOI22_X1  g638(.A1(new_n835_), .A2(new_n837_), .B1(new_n838_), .B2(new_n839_), .ZN(G1347gat));
  NAND3_X1  g639(.A1(new_n629_), .A2(new_n549_), .A3(new_n519_), .ZN(new_n841_));
  NOR3_X1   g640(.A1(new_n777_), .A2(new_n595_), .A3(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n571_), .ZN(new_n843_));
  OAI21_X1  g642(.A(KEYINPUT62), .B1(new_n843_), .B2(KEYINPUT22), .ZN(new_n844_));
  OAI21_X1  g643(.A(G169gat), .B1(new_n843_), .B2(KEYINPUT62), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n846_), .B1(new_n382_), .B2(new_n844_), .ZN(G1348gat));
  INV_X1    g646(.A(KEYINPUT124), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n841_), .A2(new_n383_), .A3(new_n355_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  AOI211_X1 g649(.A(KEYINPUT116), .B(new_n749_), .C1(new_n776_), .C2(new_n324_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n764_), .B1(new_n763_), .B2(new_n765_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n594_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(KEYINPUT123), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT123), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n786_), .A2(new_n855_), .A3(new_n594_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n850_), .B1(new_n854_), .B2(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(G176gat), .B1(new_n842_), .B2(new_n611_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n848_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n855_), .B1(new_n786_), .B2(new_n594_), .ZN(new_n860_));
  AOI211_X1 g659(.A(KEYINPUT123), .B(new_n595_), .C1(new_n750_), .C2(new_n766_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n849_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n858_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n862_), .A2(KEYINPUT124), .A3(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n859_), .A2(new_n864_), .ZN(G1349gat));
  NOR2_X1   g664(.A1(new_n841_), .A2(new_n595_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n770_), .A2(new_n866_), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n867_), .A2(new_n324_), .A3(new_n388_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n841_), .A2(new_n324_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n869_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n870_));
  INV_X1    g669(.A(G183gat), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n868_), .B1(new_n870_), .B2(new_n871_), .ZN(G1350gat));
  NAND2_X1  g671(.A1(new_n842_), .A2(new_n615_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(G190gat), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n842_), .A2(new_n280_), .A3(new_n389_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(KEYINPUT125), .ZN(G1351gat));
  NOR2_X1   g676(.A1(new_n573_), .A2(new_n550_), .ZN(new_n878_));
  XOR2_X1   g677(.A(new_n878_), .B(KEYINPUT126), .Z(new_n879_));
  AOI211_X1 g678(.A(new_n663_), .B(new_n879_), .C1(new_n750_), .C2(new_n766_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n571_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n611_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g683(.A1(new_n880_), .A2(new_n325_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(KEYINPUT63), .B(G211gat), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n887_), .B1(new_n885_), .B2(new_n888_), .ZN(G1354gat));
  NAND2_X1  g688(.A1(new_n880_), .A2(new_n280_), .ZN(new_n890_));
  XOR2_X1   g689(.A(KEYINPUT127), .B(G218gat), .Z(new_n891_));
  AOI21_X1  g690(.A(new_n891_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n892_));
  AOI22_X1  g691(.A1(new_n890_), .A2(new_n891_), .B1(new_n880_), .B2(new_n892_), .ZN(G1355gat));
endmodule


