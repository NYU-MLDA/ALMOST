//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 1 1 0 0 0 1 0 1 0 1 0 0 0 0 0 1 1 1 1 0 1 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 0 0 0 1 0 0 1 1 1 1 0 1 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n595_, new_n596_, new_n597_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n655_, new_n656_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n842_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n848_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n863_, new_n864_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n886_, new_n888_,
    new_n889_, new_n891_, new_n892_, new_n893_, new_n894_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_,
    new_n905_;
  XNOR2_X1  g000(.A(KEYINPUT25), .B(G183gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT26), .B(G190gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NOR2_X1   g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n206_), .A2(KEYINPUT24), .A3(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n204_), .A2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT82), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n206_), .A2(KEYINPUT24), .ZN(new_n211_));
  INV_X1    g010(.A(G183gat), .ZN(new_n212_));
  INV_X1    g011(.A(G190gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT23), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  XOR2_X1   g013(.A(new_n214_), .B(KEYINPUT83), .Z(new_n215_));
  INV_X1    g014(.A(KEYINPUT23), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n216_), .A2(G183gat), .A3(G190gat), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n211_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(G176gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT22), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT84), .B1(new_n220_), .B2(G169gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT22), .B(G169gat), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n219_), .B(new_n221_), .C1(new_n222_), .C2(KEYINPUT84), .ZN(new_n223_));
  INV_X1    g022(.A(new_n207_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n214_), .A2(new_n217_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n212_), .A2(new_n213_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n224_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  AOI22_X1  g026(.A1(new_n210_), .A2(new_n218_), .B1(new_n223_), .B2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G71gat), .B(G99gat), .ZN(new_n229_));
  INV_X1    g028(.A(G43gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n229_), .B(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n228_), .B(new_n231_), .ZN(new_n232_));
  XOR2_X1   g031(.A(G127gat), .B(G134gat), .Z(new_n233_));
  XOR2_X1   g032(.A(G113gat), .B(G120gat), .Z(new_n234_));
  XOR2_X1   g033(.A(new_n233_), .B(new_n234_), .Z(new_n235_));
  XNOR2_X1  g034(.A(new_n232_), .B(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G227gat), .A2(G233gat), .ZN(new_n237_));
  INV_X1    g036(.A(G15gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT30), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(KEYINPUT31), .ZN(new_n241_));
  XOR2_X1   g040(.A(new_n236_), .B(new_n241_), .Z(new_n242_));
  XOR2_X1   g041(.A(G155gat), .B(G162gat), .Z(new_n243_));
  INV_X1    g042(.A(G141gat), .ZN(new_n244_));
  INV_X1    g043(.A(G148gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT3), .ZN(new_n247_));
  OR3_X1    g046(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G141gat), .A2(G148gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT85), .ZN(new_n250_));
  OAI211_X1 g049(.A(new_n247_), .B(new_n248_), .C1(KEYINPUT2), .C2(new_n250_), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n250_), .A2(KEYINPUT2), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n243_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT1), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n243_), .A2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n255_), .A2(new_n249_), .A3(new_n246_), .A4(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n253_), .A2(new_n257_), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n258_), .A2(KEYINPUT29), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT28), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G22gat), .B(G50gat), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n260_), .B(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT86), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G211gat), .B(G218gat), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  XOR2_X1   g065(.A(G197gat), .B(G204gat), .Z(new_n267_));
  OR2_X1    g066(.A1(new_n267_), .A2(KEYINPUT21), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(KEYINPUT21), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n266_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n265_), .B1(new_n267_), .B2(KEYINPUT21), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n273_), .B1(KEYINPUT29), .B2(new_n258_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G228gat), .A2(G233gat), .ZN(new_n275_));
  INV_X1    g074(.A(G78gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(G106gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n274_), .B(new_n279_), .ZN(new_n280_));
  OR2_X1    g079(.A1(new_n264_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n260_), .B(new_n261_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT86), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n264_), .A2(new_n284_), .A3(new_n280_), .ZN(new_n285_));
  AND2_X1   g084(.A1(new_n281_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT4), .ZN(new_n287_));
  AND3_X1   g086(.A1(new_n253_), .A2(new_n257_), .A3(KEYINPUT95), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n288_), .A2(new_n235_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n288_), .A2(new_n235_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n287_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G225gat), .A2(G233gat), .ZN(new_n293_));
  AND3_X1   g092(.A1(new_n258_), .A2(new_n287_), .A3(new_n235_), .ZN(new_n294_));
  NOR3_X1   g093(.A1(new_n292_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n290_), .A2(new_n291_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n297_), .A2(KEYINPUT97), .A3(new_n293_), .ZN(new_n298_));
  XOR2_X1   g097(.A(G1gat), .B(G29gat), .Z(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT96), .B(G85gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT0), .B(G57gat), .ZN(new_n302_));
  XOR2_X1   g101(.A(new_n301_), .B(new_n302_), .Z(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n291_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n293_), .B1(new_n305_), .B2(new_n289_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT97), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n296_), .A2(new_n298_), .A3(new_n304_), .A4(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n298_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n303_), .B1(new_n310_), .B2(new_n295_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n309_), .A2(KEYINPUT99), .A3(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT20), .ZN(new_n313_));
  INV_X1    g112(.A(new_n228_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n313_), .B1(new_n314_), .B2(new_n272_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT88), .B(KEYINPUT24), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n225_), .B1(new_n316_), .B2(new_n206_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT90), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(new_n207_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT89), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n206_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n204_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n318_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n215_), .A2(new_n217_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(new_n226_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n224_), .B1(new_n222_), .B2(new_n219_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(new_n273_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n315_), .B1(new_n325_), .B2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G226gat), .A2(G233gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n331_), .A2(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n313_), .B1(new_n228_), .B2(new_n273_), .ZN(new_n336_));
  OAI21_X1  g135(.A(KEYINPUT91), .B1(new_n318_), .B2(new_n324_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT90), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n317_), .B(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT91), .ZN(new_n340_));
  INV_X1    g139(.A(new_n323_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(new_n321_), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n339_), .A2(new_n340_), .A3(new_n342_), .A4(new_n204_), .ZN(new_n343_));
  AOI22_X1  g142(.A1(new_n337_), .A2(new_n343_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n336_), .B1(new_n344_), .B2(new_n273_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n335_), .B1(new_n334_), .B2(new_n345_), .ZN(new_n346_));
  XOR2_X1   g145(.A(G8gat), .B(G36gat), .Z(new_n347_));
  XNOR2_X1  g146(.A(G64gat), .B(G92gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  AND2_X1   g150(.A1(new_n351_), .A2(KEYINPUT32), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n346_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT99), .ZN(new_n354_));
  OAI211_X1 g153(.A(new_n354_), .B(new_n303_), .C1(new_n310_), .C2(new_n295_), .ZN(new_n355_));
  AND3_X1   g154(.A1(new_n312_), .A2(new_n353_), .A3(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n334_), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n337_), .A2(new_n343_), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n315_), .B(new_n357_), .C1(new_n358_), .C2(new_n330_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n345_), .A2(KEYINPUT92), .A3(new_n334_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(KEYINPUT92), .B1(new_n345_), .B2(new_n334_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n359_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  OR2_X1    g162(.A1(new_n363_), .A2(new_n352_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n286_), .B1(new_n356_), .B2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n351_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n363_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT94), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n351_), .B(new_n359_), .C1(new_n361_), .C2(new_n362_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n367_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n363_), .A2(KEYINPUT94), .A3(new_n366_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  OR2_X1    g171(.A1(new_n309_), .A2(KEYINPUT33), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n309_), .A2(KEYINPUT33), .ZN(new_n374_));
  INV_X1    g173(.A(new_n293_), .ZN(new_n375_));
  OR3_X1    g174(.A1(new_n292_), .A2(new_n375_), .A3(new_n294_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n304_), .B1(new_n297_), .B2(new_n375_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT98), .ZN(new_n378_));
  AOI22_X1  g177(.A1(new_n373_), .A2(new_n374_), .B1(new_n376_), .B2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n372_), .A2(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n242_), .B1(new_n365_), .B2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT27), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n370_), .A2(new_n382_), .A3(new_n371_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n312_), .A2(new_n355_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n346_), .A2(new_n366_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n385_), .A2(new_n369_), .A3(KEYINPUT27), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n383_), .A2(new_n384_), .A3(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(new_n286_), .ZN(new_n388_));
  AND3_X1   g187(.A1(new_n381_), .A2(new_n388_), .A3(KEYINPUT100), .ZN(new_n389_));
  AOI21_X1  g188(.A(KEYINPUT100), .B1(new_n381_), .B2(new_n388_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n242_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n286_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  OAI22_X1  g192(.A1(new_n389_), .A2(new_n390_), .B1(new_n387_), .B2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G99gat), .A2(G106gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(KEYINPUT6), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT6), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n397_), .A2(G99gat), .A3(G106gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n396_), .A2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT10), .B(G99gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G85gat), .A2(G92gat), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT9), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n401_), .A2(KEYINPUT64), .A3(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(G85gat), .ZN(new_n404_));
  INV_X1    g203(.A(G92gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n403_), .B(new_n406_), .C1(new_n402_), .C2(new_n401_), .ZN(new_n407_));
  AOI21_X1  g206(.A(KEYINPUT64), .B1(new_n401_), .B2(new_n402_), .ZN(new_n408_));
  OAI221_X1 g207(.A(new_n399_), .B1(G106gat), .B2(new_n400_), .C1(new_n407_), .C2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT65), .ZN(new_n410_));
  OAI22_X1  g209(.A1(new_n410_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT7), .ZN(new_n412_));
  INV_X1    g211(.A(G99gat), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n412_), .A2(new_n413_), .A3(new_n278_), .A4(KEYINPUT65), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n410_), .A2(KEYINPUT7), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n399_), .A2(new_n411_), .A3(new_n414_), .A4(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT8), .ZN(new_n417_));
  AND3_X1   g216(.A1(new_n406_), .A2(KEYINPUT66), .A3(new_n401_), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n416_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n417_), .B1(new_n416_), .B2(new_n418_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n409_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT67), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT67), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n423_), .B(new_n409_), .C1(new_n419_), .C2(new_n420_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G71gat), .B(G78gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G57gat), .B(G64gat), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n426_), .B1(KEYINPUT11), .B2(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n428_), .B1(KEYINPUT11), .B2(new_n427_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n427_), .A2(new_n426_), .A3(KEYINPUT11), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n425_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n431_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n422_), .A2(new_n433_), .A3(new_n424_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n432_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(G230gat), .A2(G233gat), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT12), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n434_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT70), .ZN(new_n441_));
  INV_X1    g240(.A(new_n409_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT68), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n443_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n414_), .A2(new_n411_), .A3(new_n415_), .ZN(new_n445_));
  AND2_X1   g244(.A1(new_n396_), .A2(new_n398_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n418_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT8), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n416_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n448_), .A2(KEYINPUT68), .A3(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n442_), .B1(new_n444_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT69), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n429_), .A2(new_n452_), .A3(new_n430_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n452_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n455_));
  OAI21_X1  g254(.A(KEYINPUT12), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n441_), .B1(new_n451_), .B2(new_n456_), .ZN(new_n457_));
  NOR3_X1   g256(.A1(new_n419_), .A2(new_n420_), .A3(new_n443_), .ZN(new_n458_));
  AOI21_X1  g257(.A(KEYINPUT68), .B1(new_n448_), .B2(new_n449_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n409_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n431_), .A2(KEYINPUT69), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n439_), .B1(new_n461_), .B2(new_n453_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n460_), .A2(KEYINPUT70), .A3(new_n462_), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n440_), .A2(new_n457_), .A3(new_n432_), .A4(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n438_), .B1(new_n464_), .B2(new_n437_), .ZN(new_n465_));
  XOR2_X1   g264(.A(G120gat), .B(G148gat), .Z(new_n466_));
  XNOR2_X1  g265(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n466_), .B(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G176gat), .B(G204gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n468_), .B(new_n469_), .ZN(new_n470_));
  OR2_X1    g269(.A1(new_n465_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n465_), .A2(new_n470_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n471_), .A2(KEYINPUT72), .A3(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(KEYINPUT72), .B1(new_n471_), .B2(new_n472_), .ZN(new_n475_));
  OR2_X1    g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT13), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n474_), .A2(new_n475_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT13), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G29gat), .B(G36gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT74), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G43gat), .B(G50gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT74), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n482_), .B(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n484_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n485_), .A2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G15gat), .B(G22gat), .ZN(new_n491_));
  INV_X1    g290(.A(G1gat), .ZN(new_n492_));
  INV_X1    g291(.A(G8gat), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT14), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n491_), .A2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G1gat), .B(G8gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n490_), .B(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n498_), .A2(G229gat), .A3(G233gat), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT80), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n490_), .A2(new_n497_), .ZN(new_n502_));
  XOR2_X1   g301(.A(new_n490_), .B(KEYINPUT15), .Z(new_n503_));
  AOI21_X1  g302(.A(new_n502_), .B1(new_n503_), .B2(new_n497_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G229gat), .A2(G233gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n501_), .A2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G113gat), .B(G141gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G169gat), .B(G197gat), .ZN(new_n509_));
  XOR2_X1   g308(.A(new_n508_), .B(new_n509_), .Z(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n507_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT81), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n501_), .A2(new_n506_), .A3(new_n510_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n512_), .A2(new_n513_), .A3(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n507_), .A2(KEYINPUT81), .A3(new_n511_), .ZN(new_n516_));
  AND2_X1   g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n481_), .A2(new_n518_), .ZN(new_n519_));
  AND2_X1   g318(.A1(new_n394_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n503_), .A2(new_n460_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n425_), .A2(new_n485_), .A3(new_n489_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G232gat), .A2(G233gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT34), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n524_), .A2(KEYINPUT35), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(KEYINPUT35), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT73), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT75), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n525_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n521_), .A2(new_n522_), .A3(new_n529_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n527_), .A2(new_n528_), .ZN(new_n531_));
  XOR2_X1   g330(.A(new_n530_), .B(new_n531_), .Z(new_n532_));
  INV_X1    g331(.A(KEYINPUT76), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(G190gat), .B(G218gat), .Z(new_n535_));
  XNOR2_X1  g334(.A(G134gat), .B(G162gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT36), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n532_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n537_), .A2(new_n538_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n534_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n541_), .ZN(new_n543_));
  OAI211_X1 g342(.A(new_n532_), .B(new_n533_), .C1(new_n543_), .C2(new_n539_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT37), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n542_), .A2(KEYINPUT37), .A3(new_n544_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  XOR2_X1   g349(.A(G127gat), .B(G155gat), .Z(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT16), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G183gat), .B(G211gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(new_n554_), .B(KEYINPUT78), .Z(new_n555_));
  INV_X1    g354(.A(KEYINPUT17), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n555_), .A2(new_n556_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G231gat), .A2(G233gat), .ZN(new_n559_));
  XOR2_X1   g358(.A(new_n497_), .B(new_n559_), .Z(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(new_n431_), .ZN(new_n561_));
  NOR3_X1   g360(.A1(new_n557_), .A2(new_n558_), .A3(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT79), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n454_), .A2(new_n455_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n565_), .A2(new_n560_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n565_), .A2(new_n560_), .ZN(new_n567_));
  XOR2_X1   g366(.A(KEYINPUT77), .B(KEYINPUT17), .Z(new_n568_));
  NOR4_X1   g367(.A1(new_n566_), .A2(new_n567_), .A3(new_n554_), .A4(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n563_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n550_), .A2(new_n571_), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n520_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n384_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n573_), .A2(new_n492_), .A3(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT38), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT101), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n545_), .A2(new_n571_), .ZN(new_n579_));
  AND2_X1   g378(.A1(new_n520_), .A2(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n492_), .B1(new_n580_), .B2(new_n574_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n581_), .B1(new_n576_), .B2(new_n575_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n578_), .A2(new_n582_), .ZN(G1324gat));
  AND2_X1   g382(.A1(new_n383_), .A2(new_n386_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n520_), .A2(new_n585_), .A3(new_n579_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(G8gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT39), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n573_), .A2(new_n493_), .A3(new_n585_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n588_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n590_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n592_), .A2(new_n593_), .ZN(G1325gat));
  AOI21_X1  g393(.A(new_n238_), .B1(new_n580_), .B2(new_n242_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT41), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n573_), .A2(new_n238_), .A3(new_n242_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(G1326gat));
  INV_X1    g397(.A(G22gat), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n599_), .B1(new_n580_), .B2(new_n286_), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n600_), .B(KEYINPUT42), .Z(new_n601_));
  NAND3_X1  g400(.A1(new_n573_), .A2(new_n599_), .A3(new_n286_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(G1327gat));
  NOR3_X1   g402(.A1(new_n481_), .A2(new_n570_), .A3(new_n518_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT43), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n394_), .A2(new_n605_), .A3(new_n550_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n605_), .B1(new_n394_), .B2(new_n550_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n604_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT44), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n394_), .A2(new_n550_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(KEYINPUT43), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(new_n606_), .ZN(new_n614_));
  AOI21_X1  g413(.A(KEYINPUT44), .B1(new_n614_), .B2(new_n604_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n611_), .A2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n616_), .A2(G29gat), .A3(new_n574_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n545_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n618_), .A2(new_n570_), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n520_), .A2(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(G29gat), .B1(new_n620_), .B2(new_n574_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n617_), .A2(KEYINPUT103), .A3(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT103), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n609_), .A2(new_n610_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n614_), .A2(KEYINPUT44), .A3(new_n604_), .ZN(new_n626_));
  AND4_X1   g425(.A1(G29gat), .A2(new_n625_), .A3(new_n574_), .A4(new_n626_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n624_), .B1(new_n627_), .B2(new_n621_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n623_), .A2(new_n628_), .ZN(G1328gat));
  NAND3_X1  g428(.A1(new_n625_), .A2(new_n626_), .A3(new_n585_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(G36gat), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT46), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n632_), .A2(KEYINPUT105), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n584_), .A2(G36gat), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n394_), .A2(new_n519_), .A3(new_n619_), .A4(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(KEYINPUT104), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n635_), .A2(KEYINPUT104), .ZN(new_n638_));
  OAI21_X1  g437(.A(KEYINPUT45), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n638_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT45), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n640_), .A2(new_n641_), .A3(new_n636_), .ZN(new_n642_));
  AOI22_X1  g441(.A1(new_n639_), .A2(new_n642_), .B1(KEYINPUT105), .B2(new_n632_), .ZN(new_n643_));
  AND3_X1   g442(.A1(new_n631_), .A2(new_n633_), .A3(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n633_), .B1(new_n631_), .B2(new_n643_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n644_), .A2(new_n645_), .ZN(G1329gat));
  NOR4_X1   g445(.A1(new_n611_), .A2(new_n615_), .A3(new_n230_), .A4(new_n391_), .ZN(new_n647_));
  AOI21_X1  g446(.A(G43gat), .B1(new_n620_), .B2(new_n242_), .ZN(new_n648_));
  OAI21_X1  g447(.A(KEYINPUT47), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n616_), .A2(G43gat), .A3(new_n242_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT47), .ZN(new_n651_));
  INV_X1    g450(.A(new_n648_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n650_), .A2(new_n651_), .A3(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n649_), .A2(new_n653_), .ZN(G1330gat));
  AOI21_X1  g453(.A(G50gat), .B1(new_n620_), .B2(new_n286_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n286_), .A2(G50gat), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n655_), .B1(new_n616_), .B2(new_n656_), .ZN(G1331gat));
  INV_X1    g456(.A(KEYINPUT107), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n394_), .A2(new_n518_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n481_), .A2(new_n579_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n658_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n660_), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n394_), .A2(KEYINPUT107), .A3(new_n518_), .A4(new_n662_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n664_), .A2(G57gat), .A3(new_n574_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT108), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n665_), .A2(new_n666_), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n659_), .A2(KEYINPUT106), .ZN(new_n669_));
  INV_X1    g468(.A(new_n481_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n670_), .B1(new_n659_), .B2(KEYINPUT106), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n669_), .A2(new_n572_), .A3(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(G57gat), .B1(new_n672_), .B2(new_n574_), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n667_), .A2(new_n668_), .A3(new_n673_), .ZN(G1332gat));
  INV_X1    g473(.A(G64gat), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n672_), .A2(new_n675_), .A3(new_n585_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT48), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n664_), .A2(new_n585_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n677_), .B1(new_n678_), .B2(G64gat), .ZN(new_n679_));
  AOI211_X1 g478(.A(KEYINPUT48), .B(new_n675_), .C1(new_n664_), .C2(new_n585_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n676_), .B1(new_n679_), .B2(new_n680_), .ZN(G1333gat));
  INV_X1    g480(.A(G71gat), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n672_), .A2(new_n682_), .A3(new_n242_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n661_), .A2(new_n242_), .A3(new_n663_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT49), .ZN(new_n685_));
  AND3_X1   g484(.A1(new_n684_), .A2(new_n685_), .A3(G71gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n685_), .B1(new_n684_), .B2(G71gat), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n683_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT109), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n688_), .B(new_n689_), .ZN(G1334gat));
  NAND3_X1  g489(.A1(new_n672_), .A2(new_n276_), .A3(new_n286_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n661_), .A2(new_n286_), .A3(new_n663_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n692_), .A2(G78gat), .A3(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n692_), .B2(G78gat), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n691_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT111), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n696_), .B(new_n697_), .ZN(G1335gat));
  NOR3_X1   g497(.A1(new_n670_), .A2(new_n570_), .A3(new_n517_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT113), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n701_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n613_), .A2(KEYINPUT113), .A3(new_n606_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n700_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n404_), .B1(new_n704_), .B2(new_n574_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n384_), .A2(G85gat), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n669_), .A2(new_n619_), .A3(new_n671_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT112), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NAND4_X1  g510(.A1(new_n669_), .A2(new_n671_), .A3(KEYINPUT112), .A4(new_n619_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n708_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n706_), .A2(new_n714_), .A3(KEYINPUT114), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT114), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n716_), .B1(new_n705_), .B2(new_n713_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(G1336gat));
  INV_X1    g517(.A(new_n704_), .ZN(new_n719_));
  OAI21_X1  g518(.A(G92gat), .B1(new_n719_), .B2(new_n584_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n711_), .A2(new_n712_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n721_), .A2(new_n405_), .A3(new_n585_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(G1337gat));
  AOI21_X1  g522(.A(new_n413_), .B1(new_n704_), .B2(new_n242_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n391_), .A2(new_n400_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n727_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT51), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n725_), .A2(new_n729_), .A3(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(KEYINPUT51), .B1(new_n724_), .B2(new_n728_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(G1338gat));
  NAND2_X1  g532(.A1(new_n699_), .A2(new_n286_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n734_), .B1(new_n613_), .B2(new_n606_), .ZN(new_n735_));
  OR3_X1    g534(.A1(new_n735_), .A2(KEYINPUT52), .A3(new_n278_), .ZN(new_n736_));
  OAI21_X1  g535(.A(KEYINPUT52), .B1(new_n735_), .B2(new_n278_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n286_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n739_), .A2(G106gat), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n741_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n742_));
  OAI21_X1  g541(.A(KEYINPUT53), .B1(new_n738_), .B2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n742_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT53), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n736_), .A2(new_n737_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n744_), .A2(new_n745_), .A3(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n743_), .A2(new_n747_), .ZN(G1339gat));
  AOI211_X1 g547(.A(new_n571_), .B(new_n517_), .C1(new_n547_), .C2(new_n548_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(new_n670_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT54), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT54), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n749_), .A2(new_n752_), .A3(new_n670_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n751_), .A2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT57), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT115), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n464_), .A2(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n433_), .B1(new_n422_), .B2(new_n424_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n759_), .B1(new_n439_), .B2(new_n434_), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n760_), .A2(KEYINPUT115), .A3(new_n457_), .A4(new_n463_), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n758_), .A2(new_n761_), .A3(KEYINPUT116), .A4(new_n437_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT55), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n763_), .B1(new_n464_), .B2(new_n437_), .ZN(new_n764_));
  OR3_X1    g563(.A1(new_n464_), .A2(new_n763_), .A3(new_n437_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n762_), .A2(new_n764_), .A3(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n436_), .B1(new_n464_), .B2(new_n757_), .ZN(new_n767_));
  AOI21_X1  g566(.A(KEYINPUT116), .B1(new_n767_), .B2(new_n761_), .ZN(new_n768_));
  OAI211_X1 g567(.A(KEYINPUT56), .B(new_n470_), .C1(new_n766_), .C2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT118), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n470_), .B1(new_n766_), .B2(new_n768_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT56), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT117), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n772_), .A2(new_n775_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n775_), .A2(new_n770_), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n470_), .B(new_n777_), .C1(new_n766_), .C2(new_n768_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n771_), .A2(new_n776_), .A3(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT119), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n517_), .A2(new_n471_), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n779_), .A2(new_n780_), .A3(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n780_), .B1(new_n779_), .B2(new_n781_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n510_), .B1(new_n498_), .B2(new_n505_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n504_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n784_), .B1(new_n785_), .B2(new_n505_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n514_), .A2(new_n786_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n479_), .A2(new_n787_), .ZN(new_n788_));
  NOR3_X1   g587(.A1(new_n782_), .A2(new_n783_), .A3(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n756_), .B1(new_n789_), .B2(new_n545_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n788_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n517_), .A2(new_n471_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n778_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n758_), .A2(new_n761_), .A3(new_n437_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT116), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n796_), .A2(new_n762_), .A3(new_n764_), .A4(new_n765_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n774_), .B1(new_n797_), .B2(new_n470_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n793_), .A2(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n792_), .B1(new_n799_), .B2(new_n771_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n791_), .B1(new_n800_), .B2(new_n780_), .ZN(new_n801_));
  OAI211_X1 g600(.A(KEYINPUT57), .B(new_n618_), .C1(new_n801_), .C2(new_n782_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n772_), .A2(new_n773_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n769_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n787_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n804_), .A2(new_n471_), .A3(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT58), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n550_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n806_), .A2(new_n807_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n790_), .A2(new_n802_), .A3(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n755_), .B1(new_n813_), .B2(new_n571_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n585_), .A2(new_n384_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n392_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n814_), .A2(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(G113gat), .B1(new_n817_), .B2(new_n517_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT59), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n819_), .B1(new_n814_), .B2(new_n816_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n816_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n618_), .B1(new_n801_), .B2(new_n782_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n811_), .B1(new_n822_), .B2(new_n756_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n570_), .B1(new_n823_), .B2(new_n802_), .ZN(new_n824_));
  OAI211_X1 g623(.A(KEYINPUT59), .B(new_n821_), .C1(new_n824_), .C2(new_n755_), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n820_), .A2(new_n825_), .A3(KEYINPUT120), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT120), .B1(new_n820_), .B2(new_n825_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n517_), .A2(G113gat), .ZN(new_n829_));
  XOR2_X1   g628(.A(new_n829_), .B(KEYINPUT121), .Z(new_n830_));
  AOI21_X1  g629(.A(new_n818_), .B1(new_n828_), .B2(new_n830_), .ZN(G1340gat));
  OR2_X1    g630(.A1(new_n670_), .A2(KEYINPUT60), .ZN(new_n832_));
  INV_X1    g631(.A(G120gat), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n817_), .B(new_n834_), .C1(KEYINPUT60), .C2(new_n833_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n670_), .B1(new_n820_), .B2(new_n825_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n835_), .B1(new_n836_), .B2(new_n833_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(KEYINPUT122), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT122), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n839_), .B(new_n835_), .C1(new_n836_), .C2(new_n833_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n840_), .ZN(G1341gat));
  INV_X1    g640(.A(G127gat), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n817_), .A2(new_n842_), .A3(new_n570_), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n826_), .A2(new_n827_), .A3(new_n571_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n843_), .B1(new_n844_), .B2(new_n842_), .ZN(G1342gat));
  INV_X1    g644(.A(G134gat), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n817_), .A2(new_n846_), .A3(new_n545_), .ZN(new_n847_));
  NOR3_X1   g646(.A1(new_n826_), .A2(new_n827_), .A3(new_n549_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n847_), .B1(new_n848_), .B2(new_n846_), .ZN(G1343gat));
  NAND2_X1  g648(.A1(new_n813_), .A2(new_n571_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n754_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT124), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n739_), .A2(new_n242_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n815_), .A2(new_n853_), .ZN(new_n854_));
  XOR2_X1   g653(.A(new_n854_), .B(KEYINPUT123), .Z(new_n855_));
  NAND3_X1  g654(.A1(new_n851_), .A2(new_n852_), .A3(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n852_), .B1(new_n851_), .B2(new_n855_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(G141gat), .B1(new_n859_), .B2(new_n518_), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n244_), .B(new_n517_), .C1(new_n857_), .C2(new_n858_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(G1344gat));
  OAI21_X1  g661(.A(G148gat), .B1(new_n859_), .B2(new_n670_), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n245_), .B(new_n481_), .C1(new_n857_), .C2(new_n858_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(G1345gat));
  XNOR2_X1  g664(.A(KEYINPUT61), .B(G155gat), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n866_), .B1(new_n859_), .B2(new_n571_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n866_), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n570_), .B(new_n868_), .C1(new_n857_), .C2(new_n858_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n867_), .A2(new_n869_), .ZN(G1346gat));
  INV_X1    g669(.A(new_n858_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n549_), .B1(new_n871_), .B2(new_n856_), .ZN(new_n872_));
  INV_X1    g671(.A(G162gat), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n545_), .A2(new_n873_), .ZN(new_n874_));
  OAI22_X1  g673(.A1(new_n872_), .A2(new_n873_), .B1(new_n859_), .B2(new_n874_), .ZN(G1347gat));
  NOR3_X1   g674(.A1(new_n584_), .A2(new_n393_), .A3(new_n574_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n851_), .A2(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(G169gat), .B1(new_n877_), .B2(new_n518_), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n878_), .A2(KEYINPUT62), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n878_), .A2(KEYINPUT62), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n517_), .A2(new_n222_), .ZN(new_n881_));
  XOR2_X1   g680(.A(new_n881_), .B(KEYINPUT125), .Z(new_n882_));
  OAI22_X1  g681(.A1(new_n879_), .A2(new_n880_), .B1(new_n877_), .B2(new_n882_), .ZN(G1348gat));
  NOR2_X1   g682(.A1(new_n877_), .A2(new_n670_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(new_n219_), .ZN(G1349gat));
  NOR2_X1   g684(.A1(new_n877_), .A2(new_n571_), .ZN(new_n886_));
  MUX2_X1   g685(.A(G183gat), .B(new_n202_), .S(new_n886_), .Z(G1350gat));
  OAI21_X1  g686(.A(G190gat), .B1(new_n877_), .B2(new_n549_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n545_), .A2(new_n203_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n877_), .B2(new_n889_), .ZN(G1351gat));
  NAND2_X1  g689(.A1(new_n853_), .A2(new_n384_), .ZN(new_n891_));
  XOR2_X1   g690(.A(new_n891_), .B(KEYINPUT126), .Z(new_n892_));
  NOR3_X1   g691(.A1(new_n814_), .A2(new_n584_), .A3(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(new_n517_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g694(.A1(new_n893_), .A2(new_n481_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g696(.A1(new_n893_), .A2(new_n570_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n899_));
  AND2_X1   g698(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n898_), .A2(new_n899_), .A3(new_n900_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n901_), .B1(new_n898_), .B2(new_n899_), .ZN(G1354gat));
  NAND2_X1  g701(.A1(new_n893_), .A2(new_n545_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(KEYINPUT127), .B(G218gat), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n549_), .A2(new_n904_), .ZN(new_n905_));
  AOI22_X1  g704(.A1(new_n903_), .A2(new_n904_), .B1(new_n893_), .B2(new_n905_), .ZN(G1355gat));
endmodule


