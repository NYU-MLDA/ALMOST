//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 1 0 1 0 0 1 1 1 0 0 0 0 1 1 1 1 0 0 0 1 0 0 1 1 0 1 0 0 0 1 0 0 1 1 0 0 1 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n807_, new_n808_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n943_, new_n944_, new_n946_, new_n947_,
    new_n948_, new_n950_, new_n952_, new_n953_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n959_, new_n960_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n971_, new_n972_, new_n973_, new_n975_, new_n977_, new_n978_,
    new_n980_, new_n981_, new_n982_, new_n983_, new_n985_, new_n986_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n993_, new_n994_;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G85gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT0), .B(G57gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT3), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G141gat), .A2(G148gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT2), .ZN(new_n210_));
  AOI22_X1  g009(.A1(new_n207_), .A2(new_n208_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(new_n209_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT2), .ZN(new_n213_));
  AND2_X1   g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n215_), .B(KEYINPUT90), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(G155gat), .A2(G162gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT89), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n218_), .B(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n217_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  XOR2_X1   g021(.A(new_n221_), .B(KEYINPUT1), .Z(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(new_n220_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n207_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(new_n225_), .A3(new_n209_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n222_), .A2(new_n226_), .ZN(new_n227_));
  XOR2_X1   g026(.A(G127gat), .B(G134gat), .Z(new_n228_));
  XOR2_X1   g027(.A(G113gat), .B(G120gat), .Z(new_n229_));
  XOR2_X1   g028(.A(new_n228_), .B(new_n229_), .Z(new_n230_));
  NAND2_X1  g029(.A1(new_n227_), .A2(new_n230_), .ZN(new_n231_));
  OR2_X1    g030(.A1(new_n231_), .A2(KEYINPUT4), .ZN(new_n232_));
  INV_X1    g031(.A(new_n230_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n233_), .A2(new_n222_), .A3(new_n226_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n231_), .A2(KEYINPUT4), .A3(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n232_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G225gat), .A2(G233gat), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n236_), .A2(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n238_), .B1(new_n231_), .B2(new_n234_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n206_), .B1(new_n239_), .B2(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n237_), .B1(new_n232_), .B2(new_n235_), .ZN(new_n243_));
  NOR3_X1   g042(.A1(new_n243_), .A2(new_n205_), .A3(new_n240_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G227gat), .A2(G233gat), .ZN(new_n247_));
  INV_X1    g046(.A(G15gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(G43gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G71gat), .B(G99gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n250_), .B(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(G183gat), .ZN(new_n254_));
  INV_X1    g053(.A(G190gat), .ZN(new_n255_));
  OAI21_X1  g054(.A(KEYINPUT23), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT84), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT23), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n258_), .A2(G183gat), .A3(G190gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G169gat), .A2(G176gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT24), .ZN(new_n262_));
  OR2_X1    g061(.A1(G169gat), .A2(G176gat), .ZN(new_n263_));
  MUX2_X1   g062(.A(KEYINPUT24), .B(new_n262_), .S(new_n263_), .Z(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT81), .B(KEYINPUT25), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(G183gat), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT82), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  OR3_X1    g067(.A1(new_n255_), .A2(KEYINPUT83), .A3(KEYINPUT26), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT26), .B1(new_n255_), .B2(KEYINPUT83), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT80), .B(G183gat), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT25), .ZN(new_n272_));
  OAI211_X1 g071(.A(new_n269_), .B(new_n270_), .C1(new_n271_), .C2(new_n272_), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n260_), .B(new_n264_), .C1(new_n268_), .C2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n256_), .A2(new_n259_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n275_), .B1(G190gat), .B2(new_n271_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT86), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  OAI211_X1 g077(.A(new_n275_), .B(KEYINPUT86), .C1(G190gat), .C2(new_n271_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT22), .B(G169gat), .ZN(new_n280_));
  INV_X1    g079(.A(G176gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(new_n261_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n283_), .A2(KEYINPUT85), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT85), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n285_), .B1(new_n282_), .B2(new_n261_), .ZN(new_n286_));
  OAI211_X1 g085(.A(new_n278_), .B(new_n279_), .C1(new_n284_), .C2(new_n286_), .ZN(new_n287_));
  AND3_X1   g086(.A1(new_n274_), .A2(KEYINPUT30), .A3(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(KEYINPUT30), .B1(new_n274_), .B2(new_n287_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n253_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n274_), .A2(new_n287_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT30), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n274_), .A2(KEYINPUT30), .A3(new_n287_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n293_), .A2(new_n294_), .A3(new_n252_), .ZN(new_n295_));
  AOI21_X1  g094(.A(KEYINPUT87), .B1(new_n290_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT88), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n297_), .B1(new_n290_), .B2(new_n295_), .ZN(new_n298_));
  XOR2_X1   g097(.A(new_n230_), .B(KEYINPUT31), .Z(new_n299_));
  OAI22_X1  g098(.A1(KEYINPUT88), .A2(new_n296_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n290_), .A2(new_n295_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT87), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n299_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n303_), .A2(new_n297_), .A3(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n300_), .A2(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G78gat), .B(G106gat), .ZN(new_n307_));
  INV_X1    g106(.A(G233gat), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n308_), .B1(KEYINPUT92), .B2(G228gat), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n309_), .B1(KEYINPUT92), .B2(G228gat), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  XOR2_X1   g110(.A(G197gat), .B(G204gat), .Z(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT21), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G197gat), .B(G204gat), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT21), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G211gat), .B(G218gat), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n313_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  OR3_X1    g117(.A1(new_n314_), .A2(new_n317_), .A3(new_n315_), .ZN(new_n319_));
  AND2_X1   g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT93), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n311_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n227_), .A2(KEYINPUT29), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n318_), .A2(new_n319_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n322_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT29), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n326_), .B1(new_n222_), .B2(new_n226_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n310_), .B1(new_n324_), .B2(KEYINPUT93), .ZN(new_n328_));
  NOR3_X1   g127(.A1(new_n327_), .A2(new_n328_), .A3(new_n320_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n307_), .B1(new_n325_), .B2(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n323_), .A2(new_n322_), .A3(new_n324_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n328_), .B1(new_n327_), .B2(new_n320_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n307_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n331_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n330_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT91), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n222_), .A2(new_n226_), .A3(new_n326_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT28), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT28), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n222_), .A2(new_n226_), .A3(new_n339_), .A4(new_n326_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G22gat), .B(G50gat), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n338_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n341_), .B1(new_n338_), .B2(new_n340_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n336_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n344_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n346_), .A2(KEYINPUT91), .A3(new_n342_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n335_), .A2(new_n345_), .A3(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n334_), .A2(KEYINPUT94), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n343_), .A2(new_n344_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT94), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n331_), .A2(new_n332_), .A3(new_n351_), .A4(new_n333_), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n349_), .A2(new_n350_), .A3(new_n352_), .A4(new_n330_), .ZN(new_n353_));
  AND2_X1   g152(.A1(new_n348_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n306_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n348_), .A2(new_n353_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n356_), .A2(new_n300_), .A3(new_n305_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n246_), .B1(new_n355_), .B2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G226gat), .A2(G233gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT19), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT25), .B(G183gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT26), .B(G190gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n264_), .A2(new_n275_), .A3(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n283_), .B(KEYINPUT95), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n254_), .A2(new_n255_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n260_), .A2(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n365_), .B1(new_n366_), .B2(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(KEYINPUT20), .B1(new_n369_), .B2(new_n320_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n274_), .A2(new_n320_), .A3(new_n287_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n360_), .B1(new_n370_), .B2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n291_), .A2(new_n324_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n360_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT95), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n283_), .B(new_n376_), .ZN(new_n377_));
  AOI22_X1  g176(.A1(new_n257_), .A2(new_n259_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n320_), .B(new_n364_), .C1(new_n377_), .C2(new_n378_), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n374_), .A2(KEYINPUT20), .A3(new_n375_), .A4(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n373_), .A2(new_n380_), .ZN(new_n381_));
  XOR2_X1   g180(.A(G8gat), .B(G36gat), .Z(new_n382_));
  XNOR2_X1  g181(.A(G64gat), .B(G92gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n381_), .A2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n373_), .A2(new_n386_), .A3(new_n380_), .ZN(new_n389_));
  AOI21_X1  g188(.A(KEYINPUT27), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(KEYINPUT27), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT98), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n379_), .A2(new_n392_), .A3(KEYINPUT20), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(new_n374_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n392_), .B1(new_n379_), .B2(KEYINPUT20), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n360_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n364_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(new_n324_), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n398_), .A2(KEYINPUT20), .A3(new_n375_), .A4(new_n371_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n386_), .B1(new_n396_), .B2(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n391_), .B1(new_n400_), .B2(KEYINPUT99), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT99), .ZN(new_n402_));
  INV_X1    g201(.A(new_n399_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n395_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n404_), .A2(new_n374_), .A3(new_n393_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n403_), .B1(new_n405_), .B2(new_n360_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n402_), .B1(new_n406_), .B2(new_n386_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n390_), .B1(new_n401_), .B2(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n205_), .B1(new_n243_), .B2(new_n240_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT33), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n231_), .A2(new_n238_), .A3(new_n234_), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n412_), .A2(new_n206_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n413_), .B1(new_n236_), .B2(new_n238_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT97), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n413_), .B(KEYINPUT97), .C1(new_n236_), .C2(new_n238_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n416_), .A2(new_n388_), .A3(new_n389_), .A4(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT32), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n387_), .A2(new_n419_), .ZN(new_n420_));
  OAI22_X1  g219(.A1(new_n242_), .A2(new_n244_), .B1(new_n381_), .B2(new_n420_), .ZN(new_n421_));
  NOR3_X1   g220(.A1(new_n406_), .A2(new_n419_), .A3(new_n387_), .ZN(new_n422_));
  OAI22_X1  g221(.A1(new_n411_), .A2(new_n418_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n306_), .A2(new_n356_), .ZN(new_n424_));
  AOI22_X1  g223(.A1(new_n358_), .A2(new_n408_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G229gat), .A2(G233gat), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G1gat), .B(G8gat), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G15gat), .B(G22gat), .ZN(new_n430_));
  INV_X1    g229(.A(G1gat), .ZN(new_n431_));
  INV_X1    g230(.A(G8gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(KEYINPUT76), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT76), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(G8gat), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n431_), .B1(new_n433_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT14), .ZN(new_n437_));
  OAI211_X1 g236(.A(KEYINPUT77), .B(new_n430_), .C1(new_n436_), .C2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(KEYINPUT76), .B(G8gat), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT14), .B1(new_n440_), .B2(new_n431_), .ZN(new_n441_));
  AOI21_X1  g240(.A(KEYINPUT77), .B1(new_n441_), .B2(new_n430_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n429_), .B1(new_n439_), .B2(new_n442_), .ZN(new_n443_));
  XOR2_X1   g242(.A(G43gat), .B(G50gat), .Z(new_n444_));
  INV_X1    g243(.A(G36gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(G29gat), .ZN(new_n446_));
  INV_X1    g245(.A(G29gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(G36gat), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n446_), .A2(new_n448_), .A3(KEYINPUT71), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(KEYINPUT71), .B1(new_n446_), .B2(new_n448_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n444_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n446_), .A2(new_n448_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT71), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G43gat), .B(G50gat), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(new_n449_), .A3(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n452_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT77), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n433_), .A2(new_n435_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n437_), .B1(new_n460_), .B2(G1gat), .ZN(new_n461_));
  INV_X1    g260(.A(new_n430_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n459_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n463_), .A2(new_n438_), .A3(new_n428_), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n443_), .A2(new_n458_), .A3(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n458_), .B1(new_n443_), .B2(new_n464_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n427_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT15), .ZN(new_n468_));
  NOR3_X1   g267(.A1(new_n450_), .A2(new_n451_), .A3(new_n444_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n456_), .B1(new_n455_), .B2(new_n449_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n468_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n452_), .A2(new_n457_), .A3(KEYINPUT15), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n473_), .A2(new_n464_), .A3(new_n443_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n458_), .ZN(new_n475_));
  NOR3_X1   g274(.A1(new_n439_), .A2(new_n442_), .A3(new_n429_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n428_), .B1(new_n463_), .B2(new_n438_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n475_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n474_), .A2(new_n478_), .A3(new_n426_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n467_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT79), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G113gat), .B(G141gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G169gat), .B(G197gat), .ZN(new_n483_));
  XOR2_X1   g282(.A(new_n482_), .B(new_n483_), .Z(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n480_), .A2(new_n481_), .A3(new_n485_), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n467_), .B(new_n479_), .C1(KEYINPUT79), .C2(new_n484_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n425_), .A2(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(G120gat), .B(G148gat), .Z(new_n491_));
  XNOR2_X1  g290(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G176gat), .B(G204gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  OR2_X1    g295(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n497_), .A2(KEYINPUT64), .A3(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT64), .ZN(new_n500_));
  AND2_X1   g299(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n501_));
  NOR2_X1   g300(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n500_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(G106gat), .B1(new_n499_), .B2(new_n503_), .ZN(new_n504_));
  AND3_X1   g303(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n505_));
  AOI21_X1  g304(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(G85gat), .ZN(new_n508_));
  INV_X1    g307(.A(G92gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G85gat), .A2(G92gat), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n510_), .A2(KEYINPUT9), .A3(new_n511_), .ZN(new_n512_));
  OR2_X1    g311(.A1(new_n511_), .A2(KEYINPUT9), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n507_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n514_));
  OR2_X1    g313(.A1(new_n504_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT8), .ZN(new_n516_));
  AND2_X1   g315(.A1(new_n510_), .A2(new_n511_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G99gat), .A2(G106gat), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT6), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n521_));
  NOR3_X1   g320(.A1(KEYINPUT65), .A2(G99gat), .A3(G106gat), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT7), .ZN(new_n523_));
  OAI211_X1 g322(.A(new_n520_), .B(new_n521_), .C1(new_n522_), .C2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT65), .ZN(new_n525_));
  INV_X1    g324(.A(G99gat), .ZN(new_n526_));
  INV_X1    g325(.A(G106gat), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n525_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n528_), .A2(KEYINPUT7), .ZN(new_n529_));
  OAI211_X1 g328(.A(new_n516_), .B(new_n517_), .C1(new_n524_), .C2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n528_), .A2(KEYINPUT7), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n522_), .A2(new_n523_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n532_), .A2(new_n507_), .A3(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n516_), .B1(new_n534_), .B2(new_n517_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n515_), .B1(new_n531_), .B2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G57gat), .B(G64gat), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT11), .ZN(new_n538_));
  XOR2_X1   g337(.A(G71gat), .B(G78gat), .Z(new_n539_));
  NOR2_X1   g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n538_), .A2(new_n539_), .ZN(new_n541_));
  OR2_X1    g340(.A1(new_n537_), .A2(KEYINPUT11), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n540_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n536_), .A2(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n504_), .A2(new_n514_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n517_), .B1(new_n524_), .B2(new_n529_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT8), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n545_), .B1(new_n547_), .B2(new_n530_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n543_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n544_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G230gat), .A2(G233gat), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n551_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(KEYINPUT66), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT66), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n551_), .A2(new_n556_), .A3(new_n553_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n553_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT67), .ZN(new_n560_));
  AOI21_X1  g359(.A(KEYINPUT12), .B1(new_n544_), .B2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT12), .ZN(new_n562_));
  AOI211_X1 g361(.A(KEYINPUT67), .B(new_n562_), .C1(new_n536_), .C2(new_n543_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n559_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n496_), .B1(new_n558_), .B2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n557_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n556_), .B1(new_n551_), .B2(new_n553_), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n564_), .B(new_n496_), .C1(new_n567_), .C2(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n566_), .A2(KEYINPUT13), .A3(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT13), .ZN(new_n571_));
  INV_X1    g370(.A(new_n569_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n571_), .B1(new_n572_), .B2(new_n565_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n570_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n575_), .A2(KEYINPUT69), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(KEYINPUT69), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G190gat), .B(G218gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G134gat), .B(G162gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n581_), .B(KEYINPUT36), .Z(new_n582_));
  XNOR2_X1  g381(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n583_));
  AND2_X1   g382(.A1(G232gat), .A2(G233gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  OAI22_X1  g384(.A1(new_n536_), .A2(new_n458_), .B1(KEYINPUT35), .B2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n547_), .A2(new_n530_), .ZN(new_n587_));
  AOI22_X1  g386(.A1(new_n587_), .A2(new_n515_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n585_), .A2(KEYINPUT35), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NOR3_X1   g389(.A1(new_n586_), .A2(new_n588_), .A3(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n585_), .A2(KEYINPUT35), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n592_), .B1(new_n548_), .B2(new_n475_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n473_), .A2(new_n536_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n589_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n582_), .B1(new_n591_), .B2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(KEYINPUT74), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n590_), .B1(new_n586_), .B2(new_n588_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n593_), .A2(new_n589_), .A3(new_n594_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT74), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n600_), .A2(new_n601_), .A3(new_n582_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n597_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT37), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n581_), .A2(KEYINPUT36), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n598_), .A2(new_n605_), .A3(new_n599_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(KEYINPUT72), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT72), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n598_), .A2(new_n608_), .A3(new_n605_), .A4(new_n599_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n607_), .A2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n603_), .A2(new_n604_), .A3(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(KEYINPUT75), .ZN(new_n612_));
  AOI22_X1  g411(.A1(new_n597_), .A2(new_n602_), .B1(new_n607_), .B2(new_n609_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT75), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n613_), .A2(new_n614_), .A3(new_n604_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n582_), .B(KEYINPUT73), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n600_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n610_), .A2(new_n617_), .ZN(new_n618_));
  AOI22_X1  g417(.A1(new_n612_), .A2(new_n615_), .B1(KEYINPUT37), .B2(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n476_), .A2(new_n477_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G127gat), .B(G155gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT16), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G183gat), .B(G211gat), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT16), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n622_), .B(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n624_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n625_), .A2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT17), .ZN(new_n631_));
  NAND2_X1  g430(.A1(G231gat), .A2(G233gat), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n631_), .A2(KEYINPUT78), .A3(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n632_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT17), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n635_), .B1(new_n625_), .B2(new_n629_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT78), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n634_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n633_), .A2(new_n543_), .A3(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n543_), .B1(new_n633_), .B2(new_n638_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n621_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n632_), .B1(new_n631_), .B2(KEYINPUT78), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n636_), .A2(new_n637_), .A3(new_n634_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n549_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n645_), .A2(new_n620_), .A3(new_n639_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n625_), .A2(new_n629_), .A3(new_n635_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n642_), .A2(new_n646_), .A3(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n619_), .A2(new_n649_), .ZN(new_n650_));
  AND3_X1   g449(.A1(new_n490_), .A2(new_n578_), .A3(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n651_), .A2(new_n431_), .A3(new_n246_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT38), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT102), .Z(new_n655_));
  NOR2_X1   g454(.A1(new_n652_), .A2(new_n653_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT100), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n425_), .A2(new_n613_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n575_), .A2(new_n488_), .A3(new_n648_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT101), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n659_), .A2(new_n660_), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n658_), .A2(new_n661_), .A3(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(G1gat), .B1(new_n664_), .B2(new_n245_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n655_), .A2(new_n657_), .A3(new_n665_), .ZN(G1324gat));
  INV_X1    g465(.A(new_n408_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n651_), .A2(new_n667_), .A3(new_n440_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT39), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n663_), .A2(new_n667_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n669_), .B1(new_n670_), .B2(G8gat), .ZN(new_n671_));
  AOI211_X1 g470(.A(KEYINPUT39), .B(new_n432_), .C1(new_n663_), .C2(new_n667_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n668_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT40), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n673_), .B(new_n674_), .ZN(G1325gat));
  NAND3_X1  g474(.A1(new_n651_), .A2(new_n248_), .A3(new_n306_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n663_), .A2(new_n306_), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n677_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n678_));
  AOI21_X1  g477(.A(KEYINPUT41), .B1(new_n677_), .B2(G15gat), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n676_), .B1(new_n678_), .B2(new_n679_), .ZN(G1326gat));
  INV_X1    g479(.A(G22gat), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n651_), .A2(new_n681_), .A3(new_n356_), .ZN(new_n682_));
  OAI21_X1  g481(.A(G22gat), .B1(new_n664_), .B2(new_n354_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n683_), .A2(KEYINPUT42), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n683_), .A2(KEYINPUT42), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n682_), .B1(new_n684_), .B2(new_n685_), .ZN(G1327gat));
  INV_X1    g485(.A(KEYINPUT104), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n618_), .A2(KEYINPUT37), .ZN(new_n688_));
  AND4_X1   g487(.A1(new_n614_), .A2(new_n603_), .A3(new_n604_), .A4(new_n610_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n614_), .B1(new_n613_), .B2(new_n604_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n688_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(KEYINPUT43), .B1(new_n425_), .B2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n357_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n356_), .B1(new_n300_), .B2(new_n305_), .ZN(new_n694_));
  OAI211_X1 g493(.A(new_n408_), .B(new_n245_), .C1(new_n693_), .C2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n423_), .A2(new_n424_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT43), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n697_), .A2(new_n698_), .A3(new_n619_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n692_), .A2(new_n699_), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n574_), .A2(new_n489_), .A3(new_n648_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n687_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n701_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n705_), .B1(new_n692_), .B2(new_n699_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n706_), .A2(KEYINPUT104), .A3(KEYINPUT44), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n704_), .A2(new_n707_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(KEYINPUT103), .B(KEYINPUT44), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  AOI211_X1 g509(.A(new_n447_), .B(new_n245_), .C1(new_n702_), .C2(new_n710_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n708_), .A2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n613_), .A2(new_n649_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n574_), .A2(new_n713_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n490_), .A2(new_n714_), .ZN(new_n715_));
  AOI21_X1  g514(.A(G29gat), .B1(new_n715_), .B2(new_n246_), .ZN(new_n716_));
  OAI21_X1  g515(.A(KEYINPUT105), .B1(new_n712_), .B2(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n716_), .B1(new_n708_), .B2(new_n711_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT105), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n717_), .A2(new_n720_), .ZN(G1328gat));
  INV_X1    g520(.A(KEYINPUT107), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n722_), .A2(KEYINPUT46), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n667_), .B1(new_n706_), .B2(new_n709_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n445_), .B1(new_n708_), .B2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT45), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n408_), .A2(G36gat), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n490_), .A2(new_n714_), .A3(new_n728_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n729_), .A2(KEYINPUT106), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n729_), .A2(KEYINPUT106), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n727_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  OR2_X1    g531(.A1(new_n729_), .A2(KEYINPUT106), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n729_), .A2(KEYINPUT106), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n733_), .A2(KEYINPUT45), .A3(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n732_), .A2(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n723_), .B1(new_n726_), .B2(new_n736_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n732_), .A2(new_n735_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n723_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n724_), .B1(new_n704_), .B2(new_n707_), .ZN(new_n740_));
  OAI211_X1 g539(.A(new_n738_), .B(new_n739_), .C1(new_n445_), .C2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n737_), .A2(new_n741_), .ZN(G1329gat));
  XNOR2_X1  g541(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n702_), .A2(new_n710_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n745_), .A2(G43gat), .A3(new_n306_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n746_), .B1(new_n704_), .B2(new_n707_), .ZN(new_n747_));
  AOI21_X1  g546(.A(G43gat), .B1(new_n715_), .B2(new_n306_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n744_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n745_), .A2(G43gat), .A3(new_n306_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n748_), .B1(new_n750_), .B2(new_n708_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(new_n743_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n749_), .A2(new_n752_), .ZN(G1330gat));
  INV_X1    g552(.A(G50gat), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n715_), .A2(new_n754_), .A3(new_n356_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n356_), .B1(new_n706_), .B2(new_n709_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n756_), .B1(new_n704_), .B2(new_n707_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(KEYINPUT109), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(G50gat), .B1(new_n757_), .B2(KEYINPUT109), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n755_), .B1(new_n759_), .B2(new_n760_), .ZN(G1331gat));
  INV_X1    g560(.A(new_n578_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n649_), .A2(new_n488_), .ZN(new_n763_));
  AND3_X1   g562(.A1(new_n762_), .A2(new_n658_), .A3(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n764_), .A2(G57gat), .A3(new_n246_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT111), .ZN(new_n766_));
  OR3_X1    g565(.A1(new_n425_), .A2(KEYINPUT110), .A3(new_n488_), .ZN(new_n767_));
  OAI21_X1  g566(.A(KEYINPUT110), .B1(new_n425_), .B2(new_n488_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n769_), .A2(new_n574_), .A3(new_n650_), .ZN(new_n770_));
  AOI21_X1  g569(.A(G57gat), .B1(new_n770_), .B2(new_n246_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n766_), .A2(new_n771_), .ZN(G1332gat));
  INV_X1    g571(.A(G64gat), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n770_), .A2(new_n773_), .A3(new_n667_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n764_), .A2(new_n667_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(G64gat), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n776_), .A2(KEYINPUT48), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n776_), .A2(KEYINPUT48), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n774_), .B1(new_n777_), .B2(new_n778_), .ZN(G1333gat));
  INV_X1    g578(.A(G71gat), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n770_), .A2(new_n780_), .A3(new_n306_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n764_), .A2(new_n306_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(G71gat), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n783_), .A2(KEYINPUT49), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n783_), .A2(KEYINPUT49), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n781_), .B1(new_n784_), .B2(new_n785_), .ZN(G1334gat));
  INV_X1    g585(.A(G78gat), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n770_), .A2(new_n787_), .A3(new_n356_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n764_), .A2(new_n356_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n790_));
  AND3_X1   g589(.A1(new_n789_), .A2(G78gat), .A3(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n789_), .B2(G78gat), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n788_), .B1(new_n791_), .B2(new_n792_), .ZN(G1335gat));
  NAND4_X1  g592(.A1(new_n577_), .A2(new_n576_), .A3(new_n613_), .A4(new_n649_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n769_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT113), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n769_), .A2(KEYINPUT113), .A3(new_n795_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n800_), .A2(new_n508_), .A3(new_n246_), .ZN(new_n801_));
  NOR3_X1   g600(.A1(new_n575_), .A2(new_n488_), .A3(new_n648_), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n700_), .A2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(G85gat), .B1(new_n804_), .B2(new_n245_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n801_), .A2(new_n805_), .ZN(G1336gat));
  NAND3_X1  g605(.A1(new_n800_), .A2(new_n509_), .A3(new_n667_), .ZN(new_n807_));
  OAI21_X1  g606(.A(G92gat), .B1(new_n804_), .B2(new_n408_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(G1337gat));
  NAND2_X1  g608(.A1(new_n499_), .A2(new_n503_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n306_), .A2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n811_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n526_), .B1(new_n803_), .B2(new_n306_), .ZN(new_n813_));
  OR3_X1    g612(.A1(new_n812_), .A2(KEYINPUT51), .A3(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(KEYINPUT51), .B1(new_n812_), .B2(new_n813_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(G1338gat));
  NOR3_X1   g615(.A1(new_n425_), .A2(KEYINPUT43), .A3(new_n691_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n698_), .B1(new_n697_), .B2(new_n619_), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n356_), .B(new_n802_), .C1(new_n817_), .C2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT114), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT114), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n700_), .A2(new_n821_), .A3(new_n356_), .A4(new_n802_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n527_), .B1(KEYINPUT115), .B2(KEYINPUT52), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n820_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(KEYINPUT115), .A2(KEYINPUT52), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT113), .B1(new_n769_), .B2(new_n795_), .ZN(new_n827_));
  AOI211_X1 g626(.A(new_n797_), .B(new_n794_), .C1(new_n767_), .C2(new_n768_), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n527_), .B(new_n356_), .C1(new_n827_), .C2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n825_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n820_), .A2(new_n822_), .A3(new_n823_), .A4(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n826_), .A2(new_n829_), .A3(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT53), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT53), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n826_), .A2(new_n829_), .A3(new_n834_), .A4(new_n831_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n835_), .ZN(G1339gat));
  INV_X1    g635(.A(G113gat), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n489_), .A2(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n426_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n474_), .A2(new_n478_), .A3(new_n427_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n484_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n485_), .B1(new_n467_), .B2(new_n479_), .ZN(new_n842_));
  OAI21_X1  g641(.A(KEYINPUT118), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n839_), .A2(new_n840_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n485_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n480_), .A2(new_n484_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT118), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n845_), .A2(new_n846_), .A3(new_n847_), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n843_), .B(new_n848_), .C1(new_n572_), .C2(new_n565_), .ZN(new_n849_));
  OAI211_X1 g648(.A(KEYINPUT55), .B(new_n559_), .C1(new_n561_), .C2(new_n563_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT116), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT55), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n564_), .A2(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n550_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n553_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n560_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n562_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n544_), .A2(new_n560_), .A3(KEYINPUT12), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n860_), .A2(KEYINPUT116), .A3(KEYINPUT55), .A4(new_n559_), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n852_), .A2(new_n854_), .A3(new_n856_), .A4(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT117), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n863_), .A2(KEYINPUT56), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n862_), .A2(new_n495_), .A3(new_n864_), .ZN(new_n865_));
  AND2_X1   g664(.A1(new_n488_), .A2(new_n569_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n864_), .B1(new_n862_), .B2(new_n495_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n849_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n613_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT57), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n869_), .A2(KEYINPUT57), .A3(new_n870_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n862_), .A2(new_n495_), .ZN(new_n875_));
  XOR2_X1   g674(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(KEYINPUT119), .A2(KEYINPUT56), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n862_), .A2(new_n495_), .A3(new_n878_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n848_), .A2(new_n843_), .A3(new_n569_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n877_), .A2(new_n879_), .A3(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT58), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n880_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n885_), .A2(KEYINPUT58), .A3(new_n879_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n884_), .A2(new_n619_), .A3(new_n886_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n873_), .A2(new_n874_), .A3(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(new_n649_), .ZN(new_n889_));
  AND3_X1   g688(.A1(new_n570_), .A2(new_n763_), .A3(new_n573_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT54), .ZN(new_n891_));
  AND3_X1   g690(.A1(new_n691_), .A2(new_n890_), .A3(new_n891_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n891_), .B1(new_n691_), .B2(new_n890_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n889_), .A2(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n408_), .A2(new_n246_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(new_n694_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  AOI21_X1  g699(.A(KEYINPUT59), .B1(new_n896_), .B2(new_n900_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n894_), .B1(new_n888_), .B2(new_n649_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT59), .ZN(new_n903_));
  NOR3_X1   g702(.A1(new_n902_), .A2(new_n903_), .A3(new_n899_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n838_), .B1(new_n901_), .B2(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n899_), .B1(new_n889_), .B2(new_n895_), .ZN(new_n906_));
  AOI211_X1 g705(.A(KEYINPUT120), .B(G113gat), .C1(new_n906_), .C2(new_n488_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT120), .ZN(new_n908_));
  AOI21_X1  g707(.A(KEYINPUT58), .B1(new_n885_), .B2(new_n879_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n909_), .A2(new_n691_), .ZN(new_n910_));
  AOI22_X1  g709(.A1(new_n910_), .A2(new_n886_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n648_), .B1(new_n911_), .B2(new_n874_), .ZN(new_n912_));
  OAI211_X1 g711(.A(new_n488_), .B(new_n900_), .C1(new_n912_), .C2(new_n894_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n908_), .B1(new_n913_), .B2(new_n837_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n905_), .B1(new_n907_), .B2(new_n914_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(KEYINPUT121), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT121), .ZN(new_n917_));
  OAI211_X1 g716(.A(new_n905_), .B(new_n917_), .C1(new_n907_), .C2(new_n914_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n916_), .A2(new_n918_), .ZN(G1340gat));
  INV_X1    g718(.A(G120gat), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n896_), .A2(KEYINPUT59), .A3(new_n900_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n903_), .B1(new_n902_), .B2(new_n899_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n920_), .B1(new_n923_), .B2(new_n762_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n906_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n920_), .B1(new_n575_), .B2(KEYINPUT60), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n926_), .B1(KEYINPUT60), .B2(new_n920_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n925_), .A2(new_n927_), .ZN(new_n928_));
  OAI21_X1  g727(.A(KEYINPUT122), .B1(new_n924_), .B2(new_n928_), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT122), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n578_), .B1(new_n921_), .B2(new_n922_), .ZN(new_n931_));
  OAI221_X1 g730(.A(new_n930_), .B1(new_n925_), .B2(new_n927_), .C1(new_n931_), .C2(new_n920_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n929_), .A2(new_n932_), .ZN(G1341gat));
  NAND2_X1  g732(.A1(new_n648_), .A2(G127gat), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n934_), .B(KEYINPUT123), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n935_), .B1(new_n921_), .B2(new_n922_), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT124), .ZN(new_n937_));
  AOI21_X1  g736(.A(G127gat), .B1(new_n906_), .B2(new_n648_), .ZN(new_n938_));
  OR3_X1    g737(.A1(new_n936_), .A2(new_n937_), .A3(new_n938_), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n937_), .B1(new_n936_), .B2(new_n938_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n939_), .A2(new_n940_), .ZN(G1342gat));
  AOI21_X1  g740(.A(G134gat), .B1(new_n906_), .B2(new_n613_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n619_), .A2(G134gat), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n943_), .B(KEYINPUT125), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n942_), .B1(new_n923_), .B2(new_n944_), .ZN(G1343gat));
  NOR2_X1   g744(.A1(new_n902_), .A2(new_n357_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n946_), .A2(new_n898_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n947_), .A2(new_n489_), .ZN(new_n948_));
  XOR2_X1   g747(.A(new_n948_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g748(.A1(new_n947_), .A2(new_n578_), .ZN(new_n950_));
  XOR2_X1   g749(.A(new_n950_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g750(.A1(new_n947_), .A2(new_n649_), .ZN(new_n952_));
  XNOR2_X1  g751(.A(KEYINPUT61), .B(G155gat), .ZN(new_n953_));
  XOR2_X1   g752(.A(new_n952_), .B(new_n953_), .Z(G1346gat));
  INV_X1    g753(.A(G162gat), .ZN(new_n955_));
  NOR3_X1   g754(.A1(new_n947_), .A2(new_n955_), .A3(new_n691_), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n955_), .B1(new_n947_), .B2(new_n870_), .ZN(new_n957_));
  INV_X1    g756(.A(KEYINPUT126), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n957_), .A2(new_n958_), .ZN(new_n959_));
  OAI211_X1 g758(.A(KEYINPUT126), .B(new_n955_), .C1(new_n947_), .C2(new_n870_), .ZN(new_n960_));
  AOI21_X1  g759(.A(new_n956_), .B1(new_n959_), .B2(new_n960_), .ZN(G1347gat));
  NOR3_X1   g760(.A1(new_n408_), .A2(new_n355_), .A3(new_n246_), .ZN(new_n962_));
  AND2_X1   g761(.A1(new_n896_), .A2(new_n962_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n963_), .A2(new_n488_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n964_), .A2(G169gat), .ZN(new_n965_));
  INV_X1    g764(.A(KEYINPUT62), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n965_), .A2(new_n966_), .ZN(new_n967_));
  NAND3_X1  g766(.A1(new_n964_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n968_));
  INV_X1    g767(.A(new_n280_), .ZN(new_n969_));
  OAI211_X1 g768(.A(new_n967_), .B(new_n968_), .C1(new_n969_), .C2(new_n964_), .ZN(G1348gat));
  NAND3_X1  g769(.A1(new_n963_), .A2(new_n281_), .A3(new_n574_), .ZN(new_n971_));
  NAND2_X1  g770(.A1(new_n896_), .A2(new_n962_), .ZN(new_n972_));
  OAI21_X1  g771(.A(G176gat), .B1(new_n972_), .B2(new_n578_), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n971_), .A2(new_n973_), .ZN(G1349gat));
  NOR2_X1   g773(.A1(new_n972_), .A2(new_n649_), .ZN(new_n975_));
  MUX2_X1   g774(.A(new_n271_), .B(new_n361_), .S(new_n975_), .Z(G1350gat));
  NAND3_X1  g775(.A1(new_n963_), .A2(new_n362_), .A3(new_n613_), .ZN(new_n977_));
  OAI21_X1  g776(.A(G190gat), .B1(new_n972_), .B2(new_n691_), .ZN(new_n978_));
  NAND2_X1  g777(.A1(new_n977_), .A2(new_n978_), .ZN(G1351gat));
  NOR2_X1   g778(.A1(new_n408_), .A2(new_n246_), .ZN(new_n980_));
  NAND2_X1  g779(.A1(new_n946_), .A2(new_n980_), .ZN(new_n981_));
  INV_X1    g780(.A(new_n981_), .ZN(new_n982_));
  NAND2_X1  g781(.A1(new_n982_), .A2(new_n488_), .ZN(new_n983_));
  XNOR2_X1  g782(.A(new_n983_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g783(.A1(new_n981_), .A2(new_n578_), .ZN(new_n985_));
  XNOR2_X1  g784(.A(KEYINPUT127), .B(G204gat), .ZN(new_n986_));
  XNOR2_X1  g785(.A(new_n985_), .B(new_n986_), .ZN(G1353gat));
  NOR2_X1   g786(.A1(new_n981_), .A2(new_n649_), .ZN(new_n988_));
  NOR2_X1   g787(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n989_));
  AND2_X1   g788(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n990_));
  OAI21_X1  g789(.A(new_n988_), .B1(new_n989_), .B2(new_n990_), .ZN(new_n991_));
  OAI21_X1  g790(.A(new_n991_), .B1(new_n988_), .B2(new_n989_), .ZN(G1354gat));
  OR3_X1    g791(.A1(new_n981_), .A2(G218gat), .A3(new_n870_), .ZN(new_n993_));
  OAI21_X1  g792(.A(G218gat), .B1(new_n981_), .B2(new_n691_), .ZN(new_n994_));
  NAND2_X1  g793(.A1(new_n993_), .A2(new_n994_), .ZN(G1355gat));
endmodule


