//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 1 1 1 0 0 0 0 0 0 1 1 1 0 1 1 0 0 0 0 1 0 1 0 0 1 0 0 1 1 0 0 0 0 1 1 1 0 0 0 0 1 0 0 1 0 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n745_, new_n746_, new_n747_,
    new_n749_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n766_, new_n767_, new_n768_, new_n770_,
    new_n771_, new_n772_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n794_, new_n795_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n900_,
    new_n902_, new_n903_, new_n905_, new_n906_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_, new_n920_, new_n921_, new_n923_,
    new_n925_, new_n926_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n933_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_, new_n943_;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(new_n202_), .B(G15gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(G43gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G71gat), .B(G99gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT84), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT23), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  OR2_X1    g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT22), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(G169gat), .ZN(new_n217_));
  INV_X1    g016(.A(G176gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(KEYINPUT82), .A2(G169gat), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(KEYINPUT82), .A2(G169gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT22), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n219_), .B1(new_n223_), .B2(KEYINPUT83), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT83), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n225_), .B(KEYINPUT22), .C1(new_n221_), .C2(new_n222_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n215_), .B1(new_n224_), .B2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT25), .B(G183gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT26), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(G190gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT81), .ZN(new_n231_));
  INV_X1    g030(.A(G190gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n231_), .A2(new_n232_), .A3(KEYINPUT26), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT81), .B1(new_n229_), .B2(G190gat), .ZN(new_n234_));
  AND4_X1   g033(.A1(new_n228_), .A2(new_n230_), .A3(new_n233_), .A4(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n212_), .ZN(new_n236_));
  AOI21_X1  g035(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(G169gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(new_n218_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n240_), .A2(KEYINPUT24), .A3(new_n214_), .ZN(new_n241_));
  OR3_X1    g040(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n238_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n235_), .A2(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n207_), .B1(new_n227_), .B2(new_n244_), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n213_), .A2(new_n214_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n219_), .ZN(new_n247_));
  OR2_X1    g046(.A1(KEYINPUT82), .A2(G169gat), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n216_), .B1(new_n248_), .B2(new_n220_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n247_), .B1(new_n249_), .B2(new_n225_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n226_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n246_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  AND2_X1   g051(.A1(new_n241_), .A2(new_n242_), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n228_), .A2(new_n230_), .A3(new_n233_), .A4(new_n234_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n253_), .A2(new_n238_), .A3(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n252_), .A2(KEYINPUT84), .A3(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n245_), .A2(new_n256_), .A3(KEYINPUT30), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(KEYINPUT30), .B1(new_n245_), .B2(new_n256_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n206_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n259_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n206_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n261_), .A2(new_n262_), .A3(new_n257_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n205_), .B1(new_n260_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G127gat), .B(G134gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G113gat), .B(G120gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT31), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(KEYINPUT85), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(KEYINPUT86), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n260_), .A2(new_n263_), .A3(new_n205_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n265_), .A2(new_n272_), .A3(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT86), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n272_), .B1(new_n275_), .B2(new_n269_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n273_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n276_), .B1(new_n277_), .B2(new_n264_), .ZN(new_n278_));
  AND2_X1   g077(.A1(new_n274_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G225gat), .A2(G233gat), .ZN(new_n280_));
  INV_X1    g079(.A(G155gat), .ZN(new_n281_));
  INV_X1    g080(.A(G162gat), .ZN(new_n282_));
  OAI21_X1  g081(.A(KEYINPUT1), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT1), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n284_), .A2(G155gat), .A3(G162gat), .ZN(new_n285_));
  OAI21_X1  g084(.A(KEYINPUT87), .B1(G155gat), .B2(G162gat), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  NOR3_X1   g086(.A1(KEYINPUT87), .A2(G155gat), .A3(G162gat), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n283_), .B(new_n285_), .C1(new_n287_), .C2(new_n288_), .ZN(new_n289_));
  XOR2_X1   g088(.A(G141gat), .B(G148gat), .Z(new_n290_));
  NOR2_X1   g089(.A1(G141gat), .A2(G148gat), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT3), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G141gat), .A2(G148gat), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT2), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n298_));
  NAND4_X1  g097(.A1(new_n293_), .A2(new_n296_), .A3(new_n297_), .A4(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT87), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n300_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n301_));
  AOI22_X1  g100(.A1(new_n301_), .A2(new_n286_), .B1(G155gat), .B2(G162gat), .ZN(new_n302_));
  AOI22_X1  g101(.A1(new_n289_), .A2(new_n290_), .B1(new_n299_), .B2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(new_n268_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n289_), .A2(new_n290_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n299_), .A2(new_n302_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  XOR2_X1   g106(.A(new_n266_), .B(new_n267_), .Z(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  OAI211_X1 g108(.A(KEYINPUT4), .B(new_n304_), .C1(new_n309_), .C2(KEYINPUT94), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT94), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT4), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n307_), .A2(new_n308_), .A3(new_n311_), .A4(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n280_), .B1(new_n310_), .B2(new_n313_), .ZN(new_n314_));
  AND2_X1   g113(.A1(new_n309_), .A2(new_n304_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n280_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  XOR2_X1   g116(.A(G1gat), .B(G29gat), .Z(new_n318_));
  XNOR2_X1  g117(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G57gat), .B(G85gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  OR3_X1    g121(.A1(new_n314_), .A2(new_n317_), .A3(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n322_), .B1(new_n314_), .B2(new_n317_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT89), .B(G106gat), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  OR2_X1    g126(.A1(G197gat), .A2(G204gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G197gat), .A2(G204gat), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n328_), .A2(KEYINPUT21), .A3(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(G218gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(G211gat), .ZN(new_n333_));
  INV_X1    g132(.A(G211gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(G218gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT88), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT88), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n333_), .A2(new_n335_), .A3(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n331_), .A2(new_n337_), .A3(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G197gat), .B(G204gat), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT21), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  AND3_X1   g142(.A1(new_n333_), .A2(new_n335_), .A3(new_n338_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n338_), .B1(new_n333_), .B2(new_n335_), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n343_), .B(new_n330_), .C1(new_n344_), .C2(new_n345_), .ZN(new_n346_));
  AOI22_X1  g145(.A1(new_n307_), .A2(KEYINPUT29), .B1(new_n340_), .B2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT28), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT29), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n348_), .B1(new_n303_), .B2(new_n349_), .ZN(new_n350_));
  AND4_X1   g149(.A1(new_n348_), .A2(new_n305_), .A3(new_n349_), .A4(new_n306_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n347_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n346_), .A2(new_n340_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n353_), .B1(new_n303_), .B2(new_n349_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n305_), .A2(new_n349_), .A3(new_n306_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT28), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n303_), .A2(new_n348_), .A3(new_n349_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n354_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G22gat), .B(G50gat), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n352_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n359_), .B1(new_n352_), .B2(new_n358_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G228gat), .A2(G233gat), .ZN(new_n363_));
  XOR2_X1   g162(.A(new_n363_), .B(G78gat), .Z(new_n364_));
  NOR3_X1   g163(.A1(new_n361_), .A2(new_n362_), .A3(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n364_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n352_), .A2(new_n358_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n359_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n366_), .B1(new_n369_), .B2(new_n360_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n327_), .B1(new_n365_), .B2(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n364_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n369_), .A2(new_n360_), .A3(new_n366_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n372_), .A2(new_n373_), .A3(new_n326_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n325_), .B1(new_n371_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT27), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT26), .B(G190gat), .ZN(new_n377_));
  AOI211_X1 g176(.A(new_n237_), .B(new_n236_), .C1(new_n228_), .C2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(new_n253_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n239_), .A2(KEYINPUT22), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n217_), .A2(new_n380_), .A3(new_n218_), .ZN(new_n381_));
  AND3_X1   g180(.A1(new_n381_), .A2(KEYINPUT90), .A3(new_n214_), .ZN(new_n382_));
  AOI21_X1  g181(.A(KEYINPUT90), .B1(new_n381_), .B2(new_n214_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n213_), .B(KEYINPUT91), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT92), .ZN(new_n386_));
  NOR3_X1   g185(.A1(new_n384_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n381_), .A2(new_n214_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT90), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n381_), .A2(KEYINPUT90), .A3(new_n214_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT91), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n213_), .B(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(KEYINPUT92), .B1(new_n392_), .B2(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n379_), .B1(new_n387_), .B2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(new_n353_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G226gat), .A2(G233gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT19), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n353_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n245_), .A2(new_n256_), .A3(new_n401_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n397_), .A2(KEYINPUT20), .A3(new_n400_), .A4(new_n402_), .ZN(new_n403_));
  NOR3_X1   g202(.A1(new_n227_), .A2(new_n244_), .A3(new_n207_), .ZN(new_n404_));
  AOI21_X1  g203(.A(KEYINPUT84), .B1(new_n252_), .B2(new_n255_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n353_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n401_), .B(new_n379_), .C1(new_n384_), .C2(new_n385_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n406_), .A2(KEYINPUT20), .A3(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(new_n399_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n403_), .A2(new_n409_), .ZN(new_n410_));
  XOR2_X1   g209(.A(G8gat), .B(G36gat), .Z(new_n411_));
  XNOR2_X1  g210(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G64gat), .B(G92gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n376_), .B1(new_n410_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT97), .ZN(new_n417_));
  INV_X1    g216(.A(new_n379_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n386_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n392_), .A2(new_n394_), .A3(KEYINPUT92), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n418_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  OAI211_X1 g220(.A(KEYINPUT20), .B(new_n402_), .C1(new_n421_), .C2(new_n401_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n399_), .B1(new_n421_), .B2(new_n401_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT20), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n245_), .A2(new_n256_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n424_), .B1(new_n425_), .B2(new_n353_), .ZN(new_n426_));
  AOI22_X1  g225(.A1(new_n422_), .A2(new_n399_), .B1(new_n423_), .B2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n415_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n417_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n422_), .A2(new_n399_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n423_), .A2(new_n426_), .ZN(new_n431_));
  AND4_X1   g230(.A1(new_n417_), .A2(new_n430_), .A3(new_n428_), .A4(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n416_), .B1(new_n429_), .B2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n430_), .A2(new_n431_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(new_n415_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n427_), .A2(new_n428_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(KEYINPUT98), .B1(new_n437_), .B2(new_n376_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT98), .ZN(new_n439_));
  AOI211_X1 g238(.A(new_n439_), .B(KEYINPUT27), .C1(new_n435_), .C2(new_n436_), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n375_), .B(new_n433_), .C1(new_n438_), .C2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n410_), .A2(KEYINPUT32), .A3(new_n428_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT32), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n427_), .B1(new_n443_), .B2(new_n415_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n442_), .A2(new_n325_), .A3(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT33), .ZN(new_n446_));
  OR3_X1    g245(.A1(new_n324_), .A2(KEYINPUT96), .A3(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n310_), .A2(new_n280_), .A3(new_n313_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n322_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n449_));
  AOI22_X1  g248(.A1(new_n324_), .A2(new_n446_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(KEYINPUT96), .B1(new_n324_), .B2(new_n446_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n447_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n445_), .B1(new_n452_), .B2(new_n437_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n371_), .A2(new_n374_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n279_), .B1(new_n441_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n325_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n274_), .A2(new_n278_), .A3(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n459_), .A2(new_n454_), .ZN(new_n460_));
  AND3_X1   g259(.A1(new_n430_), .A2(new_n428_), .A3(new_n431_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n428_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n376_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n439_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n437_), .A2(KEYINPUT98), .A3(new_n376_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  AND3_X1   g265(.A1(new_n460_), .A2(new_n466_), .A3(new_n433_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n457_), .A2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G29gat), .B(G36gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n469_), .B(KEYINPUT71), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G43gat), .B(G50gat), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n470_), .B(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT15), .ZN(new_n474_));
  NOR2_X1   g273(.A1(G85gat), .A2(G92gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G85gat), .A2(G92gat), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n475_), .B1(new_n477_), .B2(KEYINPUT9), .ZN(new_n478_));
  NOR3_X1   g277(.A1(new_n477_), .A2(KEYINPUT65), .A3(KEYINPUT9), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT65), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT9), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n480_), .B1(new_n476_), .B2(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n478_), .B1(new_n479_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G99gat), .A2(G106gat), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT6), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(KEYINPUT10), .B(G99gat), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT64), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n488_), .B(new_n489_), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n483_), .B(new_n487_), .C1(new_n490_), .C2(G106gat), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n477_), .A2(new_n475_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(G99gat), .A2(G106gat), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT7), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n492_), .B1(new_n495_), .B2(new_n486_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(KEYINPUT8), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT8), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n498_), .B(new_n492_), .C1(new_n495_), .C2(new_n486_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n497_), .A2(KEYINPUT67), .A3(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(KEYINPUT67), .B1(new_n497_), .B2(new_n499_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n491_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n474_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n497_), .A2(new_n499_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(new_n491_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n470_), .B(new_n471_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT35), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G232gat), .A2(G233gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(KEYINPUT34), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n508_), .B1(new_n509_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n504_), .A2(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n512_), .A2(new_n509_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n504_), .B(new_n513_), .C1(new_n509_), .C2(new_n512_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n516_), .A2(KEYINPUT72), .A3(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G190gat), .B(G218gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G134gat), .B(G162gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n521_), .A2(KEYINPUT36), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n518_), .A2(new_n523_), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n516_), .A2(KEYINPUT72), .A3(new_n517_), .A4(new_n522_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n516_), .A2(new_n517_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n527_), .A2(KEYINPUT36), .A3(new_n521_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n526_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G230gat), .A2(G233gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G57gat), .B(G64gat), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT11), .ZN(new_n532_));
  XOR2_X1   g331(.A(G71gat), .B(G78gat), .Z(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n531_), .A2(KEYINPUT11), .ZN(new_n535_));
  OR2_X1    g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n532_), .A2(new_n533_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n506_), .A2(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n538_), .A2(new_n505_), .A3(new_n491_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n530_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT66), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT68), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n544_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n537_), .B(new_n544_), .C1(new_n535_), .C2(new_n534_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n545_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT69), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n503_), .A2(new_n548_), .A3(new_n549_), .A4(KEYINPUT12), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT67), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n505_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n490_), .ZN(new_n553_));
  INV_X1    g352(.A(G106gat), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n486_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  AOI22_X1  g354(.A1(new_n552_), .A2(new_n500_), .B1(new_n483_), .B2(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(KEYINPUT12), .B1(new_n545_), .B2(new_n547_), .ZN(new_n557_));
  OAI21_X1  g356(.A(KEYINPUT69), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n538_), .B1(new_n505_), .B2(new_n491_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n541_), .B1(new_n559_), .B2(KEYINPUT12), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n550_), .A2(new_n558_), .A3(new_n561_), .A4(new_n530_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n543_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G120gat), .B(G148gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT5), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G176gat), .B(G204gat), .ZN(new_n566_));
  XOR2_X1   g365(.A(new_n565_), .B(new_n566_), .Z(new_n567_));
  XOR2_X1   g366(.A(new_n567_), .B(KEYINPUT70), .Z(new_n568_));
  NAND2_X1  g367(.A1(new_n563_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n567_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n543_), .A2(new_n562_), .A3(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  OR2_X1    g371(.A1(new_n572_), .A2(KEYINPUT13), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(KEYINPUT13), .ZN(new_n574_));
  AND2_X1   g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  XOR2_X1   g374(.A(G1gat), .B(G8gat), .Z(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT75), .ZN(new_n578_));
  XOR2_X1   g377(.A(KEYINPUT74), .B(G15gat), .Z(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(G22gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(KEYINPUT74), .B(G15gat), .ZN(new_n581_));
  INV_X1    g380(.A(G22gat), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n580_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT14), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n585_), .B1(G1gat), .B2(G8gat), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n578_), .B1(new_n584_), .B2(new_n587_), .ZN(new_n588_));
  AOI211_X1 g387(.A(KEYINPUT75), .B(new_n586_), .C1(new_n580_), .C2(new_n583_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n577_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n579_), .A2(G22gat), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n581_), .A2(new_n582_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n587_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(KEYINPUT75), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n584_), .A2(new_n578_), .A3(new_n587_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n594_), .A2(new_n576_), .A3(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n590_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(new_n473_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n590_), .A2(new_n596_), .A3(new_n507_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n598_), .A2(KEYINPUT76), .A3(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G229gat), .A2(G233gat), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n597_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT76), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n603_), .A2(new_n604_), .A3(new_n507_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n600_), .A2(new_n602_), .A3(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n474_), .A2(new_n603_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n607_), .A2(new_n601_), .A3(new_n598_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G113gat), .B(G141gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G169gat), .B(G197gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(KEYINPUT77), .B(KEYINPUT78), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n612_), .B(new_n613_), .Z(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n609_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(KEYINPUT80), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n606_), .A2(new_n608_), .A3(new_n614_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT79), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT80), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n609_), .A2(new_n621_), .A3(new_n615_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n617_), .A2(new_n620_), .A3(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n618_), .A2(new_n619_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n621_), .B1(new_n609_), .B2(new_n615_), .ZN(new_n625_));
  AOI211_X1 g424(.A(KEYINPUT80), .B(new_n614_), .C1(new_n606_), .C2(new_n608_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n624_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n623_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT17), .ZN(new_n630_));
  NAND2_X1  g429(.A1(G231gat), .A2(G233gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n597_), .B(new_n631_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n632_), .A2(new_n548_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n632_), .A2(new_n548_), .ZN(new_n634_));
  XOR2_X1   g433(.A(G127gat), .B(G155gat), .Z(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT16), .ZN(new_n636_));
  XNOR2_X1  g435(.A(G183gat), .B(G211gat), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  OR4_X1    g437(.A1(new_n630_), .A2(new_n633_), .A3(new_n634_), .A4(new_n638_), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n632_), .A2(new_n538_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n632_), .A2(new_n538_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n638_), .B(KEYINPUT17), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n640_), .A2(new_n641_), .A3(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n639_), .A2(new_n643_), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n575_), .A2(new_n629_), .A3(new_n644_), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n645_), .A2(KEYINPUT100), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(KEYINPUT100), .ZN(new_n647_));
  AOI211_X1 g446(.A(new_n468_), .B(new_n529_), .C1(new_n646_), .C2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT101), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n648_), .B(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(G1gat), .B1(new_n651_), .B2(new_n458_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n468_), .A2(new_n629_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(KEYINPUT73), .B(KEYINPUT37), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n529_), .A2(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n526_), .A2(new_n528_), .A3(new_n654_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NOR3_X1   g457(.A1(new_n575_), .A2(new_n658_), .A3(new_n644_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n653_), .A2(new_n659_), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n660_), .A2(G1gat), .A3(new_n458_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n661_), .B(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n652_), .A2(new_n663_), .ZN(G1324gat));
  AOI21_X1  g463(.A(new_n529_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n466_), .A2(new_n433_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n460_), .A2(new_n466_), .A3(new_n433_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n375_), .A2(new_n433_), .ZN(new_n668_));
  AOI22_X1  g467(.A1(new_n668_), .A2(new_n466_), .B1(new_n455_), .B2(new_n453_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n667_), .B1(new_n669_), .B2(new_n279_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n665_), .A2(new_n666_), .A3(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(KEYINPUT102), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT102), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n648_), .A2(new_n673_), .A3(new_n666_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n672_), .A2(new_n674_), .A3(G8gat), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT103), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n676_), .A2(KEYINPUT39), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(KEYINPUT103), .B(KEYINPUT39), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n672_), .A2(new_n674_), .A3(G8gat), .A4(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n666_), .ZN(new_n681_));
  OR3_X1    g480(.A1(new_n660_), .A2(G8gat), .A3(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n678_), .A2(new_n680_), .A3(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT40), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n678_), .A2(KEYINPUT40), .A3(new_n680_), .A4(new_n682_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(G1325gat));
  INV_X1    g486(.A(new_n279_), .ZN(new_n688_));
  OR3_X1    g487(.A1(new_n660_), .A2(G15gat), .A3(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n650_), .A2(new_n279_), .ZN(new_n690_));
  AND3_X1   g489(.A1(new_n690_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n691_));
  AOI21_X1  g490(.A(KEYINPUT41), .B1(new_n690_), .B2(G15gat), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n689_), .B1(new_n691_), .B2(new_n692_), .ZN(G1326gat));
  INV_X1    g492(.A(KEYINPUT42), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n650_), .A2(new_n454_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n695_), .B2(G22gat), .ZN(new_n696_));
  AOI211_X1 g495(.A(KEYINPUT42), .B(new_n582_), .C1(new_n650_), .C2(new_n454_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n454_), .A2(new_n582_), .ZN(new_n698_));
  OAI22_X1  g497(.A1(new_n696_), .A2(new_n697_), .B1(new_n660_), .B2(new_n698_), .ZN(G1327gat));
  INV_X1    g498(.A(new_n644_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n529_), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n575_), .A2(new_n700_), .A3(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n653_), .A2(new_n702_), .ZN(new_n703_));
  OR3_X1    g502(.A1(new_n703_), .A2(G29gat), .A3(new_n458_), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n575_), .A2(new_n629_), .A3(new_n700_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT43), .ZN(new_n706_));
  OAI211_X1 g505(.A(new_n658_), .B(new_n706_), .C1(new_n457_), .C2(new_n467_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n706_), .B1(new_n670_), .B2(new_n658_), .ZN(new_n709_));
  OAI211_X1 g508(.A(KEYINPUT104), .B(new_n705_), .C1(new_n708_), .C2(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n705_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT104), .ZN(new_n712_));
  AOI21_X1  g511(.A(KEYINPUT44), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  OAI211_X1 g512(.A(KEYINPUT44), .B(new_n705_), .C1(new_n708_), .C2(new_n709_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT105), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n656_), .A2(new_n657_), .ZN(new_n717_));
  OAI21_X1  g516(.A(KEYINPUT43), .B1(new_n468_), .B2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(new_n707_), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n719_), .A2(KEYINPUT105), .A3(KEYINPUT44), .A4(new_n705_), .ZN(new_n720_));
  AOI22_X1  g519(.A1(new_n710_), .A2(new_n713_), .B1(new_n716_), .B2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT106), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n721_), .A2(new_n722_), .A3(new_n325_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(G29gat), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n722_), .B1(new_n721_), .B2(new_n325_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n704_), .B1(new_n724_), .B2(new_n725_), .ZN(G1328gat));
  NOR3_X1   g525(.A1(new_n703_), .A2(G36gat), .A3(new_n681_), .ZN(new_n727_));
  XOR2_X1   g526(.A(new_n727_), .B(KEYINPUT45), .Z(new_n728_));
  XNOR2_X1  g527(.A(KEYINPUT108), .B(KEYINPUT46), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n716_), .A2(new_n720_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n711_), .A2(new_n712_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT44), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n731_), .A2(new_n732_), .A3(new_n710_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT107), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n730_), .A2(new_n733_), .A3(new_n734_), .A4(new_n666_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(G36gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n734_), .B1(new_n721_), .B2(new_n666_), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n728_), .B(new_n729_), .C1(new_n736_), .C2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n730_), .A2(new_n733_), .A3(new_n666_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT107), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n741_), .A2(G36gat), .A3(new_n735_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n729_), .B1(new_n742_), .B2(new_n728_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n739_), .A2(new_n743_), .ZN(G1329gat));
  NAND3_X1  g543(.A1(new_n721_), .A2(G43gat), .A3(new_n279_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n703_), .A2(new_n688_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n745_), .B1(G43gat), .B2(new_n746_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g547(.A(new_n703_), .ZN(new_n749_));
  AOI21_X1  g548(.A(G50gat), .B1(new_n749_), .B2(new_n454_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n454_), .A2(G50gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(new_n721_), .B2(new_n751_), .ZN(G1331gat));
  NOR2_X1   g551(.A1(new_n468_), .A2(new_n628_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n753_), .A2(new_n700_), .A3(new_n575_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n754_), .A2(new_n658_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  OR3_X1    g555(.A1(new_n756_), .A2(G57gat), .A3(new_n458_), .ZN(new_n757_));
  OR2_X1    g556(.A1(new_n754_), .A2(new_n529_), .ZN(new_n758_));
  OAI21_X1  g557(.A(G57gat), .B1(new_n758_), .B2(new_n458_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(G1332gat));
  OAI21_X1  g559(.A(G64gat), .B1(new_n758_), .B2(new_n681_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT48), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n681_), .A2(G64gat), .ZN(new_n763_));
  XOR2_X1   g562(.A(new_n763_), .B(KEYINPUT109), .Z(new_n764_));
  OAI21_X1  g563(.A(new_n762_), .B1(new_n756_), .B2(new_n764_), .ZN(G1333gat));
  OAI21_X1  g564(.A(G71gat), .B1(new_n758_), .B2(new_n688_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT49), .ZN(new_n767_));
  OR2_X1    g566(.A1(new_n688_), .A2(G71gat), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n767_), .B1(new_n756_), .B2(new_n768_), .ZN(G1334gat));
  OAI21_X1  g568(.A(G78gat), .B1(new_n758_), .B2(new_n455_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT50), .ZN(new_n771_));
  OR2_X1    g570(.A1(new_n455_), .A2(G78gat), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n771_), .B1(new_n756_), .B2(new_n772_), .ZN(G1335gat));
  NAND2_X1  g572(.A1(new_n573_), .A2(new_n574_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n774_), .A2(new_n700_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n753_), .A2(new_n529_), .A3(new_n775_), .ZN(new_n776_));
  XOR2_X1   g575(.A(new_n776_), .B(KEYINPUT110), .Z(new_n777_));
  AOI21_X1  g576(.A(G85gat), .B1(new_n777_), .B2(new_n325_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT112), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n629_), .B(new_n775_), .C1(new_n708_), .C2(new_n709_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT111), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n780_), .A2(new_n781_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n779_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n784_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n786_), .A2(KEYINPUT112), .A3(new_n782_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n785_), .A2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n325_), .A2(G85gat), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT113), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n778_), .B1(new_n788_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT114), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n791_), .B(new_n792_), .ZN(G1336gat));
  AOI21_X1  g592(.A(G92gat), .B1(new_n777_), .B2(new_n666_), .ZN(new_n794_));
  AND2_X1   g593(.A1(new_n666_), .A2(G92gat), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n794_), .B1(new_n788_), .B2(new_n795_), .ZN(G1337gat));
  NAND3_X1  g595(.A1(new_n777_), .A2(new_n279_), .A3(new_n553_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n688_), .B1(new_n786_), .B2(new_n782_), .ZN(new_n798_));
  INV_X1    g597(.A(G99gat), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n797_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  XOR2_X1   g599(.A(KEYINPUT115), .B(KEYINPUT51), .Z(new_n801_));
  XNOR2_X1  g600(.A(new_n800_), .B(new_n801_), .ZN(G1338gat));
  NAND3_X1  g601(.A1(new_n777_), .A2(new_n554_), .A3(new_n454_), .ZN(new_n803_));
  OAI21_X1  g602(.A(G106gat), .B1(new_n780_), .B2(new_n455_), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n804_), .A2(KEYINPUT52), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n804_), .A2(KEYINPUT52), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n803_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n807_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n558_), .A2(new_n550_), .A3(new_n561_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n530_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n809_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n562_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n810_), .A2(new_n809_), .A3(new_n811_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n568_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT56), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n503_), .A2(new_n548_), .A3(KEYINPUT12), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n560_), .B1(new_n818_), .B2(KEYINPUT69), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n530_), .B1(new_n819_), .B2(new_n550_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n562_), .B1(new_n820_), .B2(new_n809_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n815_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT56), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n824_), .A3(new_n568_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n601_), .B1(new_n597_), .B2(new_n473_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n614_), .B1(new_n607_), .B2(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n600_), .A2(new_n601_), .A3(new_n605_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT118), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT118), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n827_), .A2(new_n828_), .A3(new_n831_), .ZN(new_n832_));
  AND4_X1   g631(.A1(new_n618_), .A2(new_n830_), .A3(new_n571_), .A4(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n817_), .A2(new_n825_), .A3(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT58), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n817_), .A2(new_n825_), .A3(KEYINPUT58), .A4(new_n833_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n836_), .A2(new_n658_), .A3(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT117), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n823_), .A2(new_n839_), .A3(new_n824_), .A4(new_n568_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n824_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n816_), .A2(new_n841_), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n628_), .A2(new_n840_), .A3(new_n571_), .A4(new_n842_), .ZN(new_n843_));
  AND3_X1   g642(.A1(new_n830_), .A2(new_n618_), .A3(new_n832_), .ZN(new_n844_));
  AND3_X1   g643(.A1(new_n844_), .A2(new_n572_), .A3(KEYINPUT119), .ZN(new_n845_));
  AOI21_X1  g644(.A(KEYINPUT119), .B1(new_n844_), .B2(new_n572_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n529_), .B1(new_n843_), .B2(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n838_), .B1(new_n848_), .B2(KEYINPUT57), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT57), .ZN(new_n850_));
  AOI211_X1 g649(.A(new_n850_), .B(new_n529_), .C1(new_n843_), .C2(new_n847_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n644_), .B1(new_n849_), .B2(new_n851_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n717_), .A2(new_n629_), .A3(new_n700_), .A4(new_n774_), .ZN(new_n853_));
  AND2_X1   g652(.A1(KEYINPUT116), .A2(KEYINPUT54), .ZN(new_n854_));
  NOR2_X1   g653(.A1(KEYINPUT116), .A2(KEYINPUT54), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n853_), .A2(new_n856_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n575_), .A2(new_n644_), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n858_), .A2(new_n629_), .A3(new_n717_), .A4(new_n854_), .ZN(new_n859_));
  AND2_X1   g658(.A1(new_n857_), .A2(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n454_), .B1(new_n852_), .B2(new_n860_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n666_), .A2(new_n458_), .A3(new_n688_), .ZN(new_n862_));
  AND3_X1   g661(.A1(new_n861_), .A2(KEYINPUT120), .A3(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(KEYINPUT120), .B1(new_n861_), .B2(new_n862_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(G113gat), .B1(new_n865_), .B2(new_n628_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n852_), .A2(new_n860_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT121), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n867_), .A2(new_n868_), .A3(new_n455_), .A4(new_n862_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT122), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n861_), .A2(new_n868_), .A3(KEYINPUT59), .A4(new_n862_), .ZN(new_n873_));
  AND3_X1   g672(.A1(new_n871_), .A2(new_n872_), .A3(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n872_), .B1(new_n871_), .B2(new_n873_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  AND2_X1   g675(.A1(new_n628_), .A2(G113gat), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n866_), .B1(new_n876_), .B2(new_n877_), .ZN(G1340gat));
  INV_X1    g677(.A(new_n865_), .ZN(new_n879_));
  INV_X1    g678(.A(G120gat), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n880_), .B1(new_n774_), .B2(KEYINPUT60), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n881_), .B1(KEYINPUT60), .B2(new_n880_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n774_), .B1(new_n871_), .B2(new_n873_), .ZN(new_n883_));
  OAI22_X1  g682(.A1(new_n879_), .A2(new_n882_), .B1(new_n883_), .B2(new_n880_), .ZN(G1341gat));
  AOI21_X1  g683(.A(G127gat), .B1(new_n865_), .B2(new_n700_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT123), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n700_), .A2(new_n886_), .A3(G127gat), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n887_), .B1(new_n886_), .B2(G127gat), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n885_), .B1(new_n876_), .B2(new_n888_), .ZN(G1342gat));
  AOI21_X1  g688(.A(G134gat), .B1(new_n865_), .B2(new_n529_), .ZN(new_n890_));
  AND2_X1   g689(.A1(new_n658_), .A2(G134gat), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n890_), .B1(new_n876_), .B2(new_n891_), .ZN(G1343gat));
  AOI21_X1  g691(.A(new_n279_), .B1(new_n852_), .B2(new_n860_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n681_), .A2(new_n325_), .A3(new_n454_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n893_), .A2(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n628_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g698(.A1(new_n897_), .A2(new_n575_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g700(.A1(new_n896_), .A2(new_n644_), .ZN(new_n902_));
  XOR2_X1   g701(.A(KEYINPUT61), .B(G155gat), .Z(new_n903_));
  XNOR2_X1  g702(.A(new_n902_), .B(new_n903_), .ZN(G1346gat));
  OAI21_X1  g703(.A(G162gat), .B1(new_n896_), .B2(new_n717_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n529_), .A2(new_n282_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n905_), .B1(new_n896_), .B2(new_n906_), .ZN(G1347gat));
  INV_X1    g706(.A(new_n861_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n681_), .A2(new_n459_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(new_n628_), .ZN(new_n910_));
  XOR2_X1   g709(.A(new_n910_), .B(KEYINPUT124), .Z(new_n911_));
  OAI21_X1  g710(.A(G169gat), .B1(new_n908_), .B2(new_n911_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n912_), .B(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n861_), .A2(new_n909_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n628_), .A2(new_n217_), .A3(new_n380_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n914_), .B1(new_n915_), .B2(new_n916_), .ZN(G1348gat));
  AND2_X1   g716(.A1(KEYINPUT126), .A2(G176gat), .ZN(new_n918_));
  NOR2_X1   g717(.A1(KEYINPUT126), .A2(G176gat), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n918_), .A2(new_n919_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n915_), .A2(new_n774_), .ZN(new_n921_));
  MUX2_X1   g720(.A(new_n918_), .B(new_n920_), .S(new_n921_), .Z(G1349gat));
  NOR2_X1   g721(.A1(new_n915_), .A2(new_n644_), .ZN(new_n923_));
  MUX2_X1   g722(.A(G183gat), .B(new_n228_), .S(new_n923_), .Z(G1350gat));
  OAI21_X1  g723(.A(G190gat), .B1(new_n915_), .B2(new_n717_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n529_), .A2(new_n377_), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n925_), .B1(new_n915_), .B2(new_n926_), .ZN(G1351gat));
  AND2_X1   g726(.A1(new_n666_), .A2(new_n375_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n893_), .A2(new_n928_), .ZN(new_n929_));
  INV_X1    g728(.A(new_n929_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n930_), .A2(new_n628_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g731(.A1(new_n930_), .A2(new_n575_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g733(.A1(new_n930_), .A2(new_n700_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n936_));
  AND2_X1   g735(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n937_));
  NOR3_X1   g736(.A1(new_n935_), .A2(new_n936_), .A3(new_n937_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n938_), .B1(new_n935_), .B2(new_n936_), .ZN(G1354gat));
  NOR3_X1   g738(.A1(new_n929_), .A2(new_n332_), .A3(new_n717_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n929_), .A2(new_n701_), .ZN(new_n941_));
  OR2_X1    g740(.A1(new_n941_), .A2(KEYINPUT127), .ZN(new_n942_));
  AOI21_X1  g741(.A(G218gat), .B1(new_n941_), .B2(KEYINPUT127), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n940_), .B1(new_n942_), .B2(new_n943_), .ZN(G1355gat));
endmodule


