//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 1 0 1 1 0 1 1 0 1 0 0 1 0 0 0 0 1 1 1 0 0 1 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 0 1 0 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n782_, new_n783_, new_n784_,
    new_n786_, new_n787_, new_n788_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n889_, new_n891_, new_n892_, new_n893_,
    new_n895_, new_n897_, new_n898_, new_n900_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n916_, new_n917_,
    new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n935_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n943_;
  XNOR2_X1  g000(.A(KEYINPUT25), .B(G183gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT26), .B(G190gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G169gat), .ZN(new_n205_));
  INV_X1    g004(.A(G176gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  OR2_X1    g006(.A1(new_n207_), .A2(KEYINPUT24), .ZN(new_n208_));
  AND2_X1   g007(.A1(new_n204_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT81), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n207_), .A2(KEYINPUT24), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(G183gat), .ZN(new_n216_));
  INV_X1    g015(.A(G190gat), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT23), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT23), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n219_), .A2(G183gat), .A3(G190gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n209_), .A2(new_n215_), .A3(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT22), .B(G169gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(new_n206_), .ZN(new_n224_));
  AND2_X1   g023(.A1(new_n224_), .A2(new_n212_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(G183gat), .A2(G190gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n218_), .A2(KEYINPUT82), .A3(new_n220_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT82), .ZN(new_n228_));
  OAI211_X1 g027(.A(new_n228_), .B(KEYINPUT23), .C1(new_n216_), .C2(new_n217_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n227_), .A2(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n225_), .B1(new_n226_), .B2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n222_), .A2(new_n231_), .ZN(new_n232_));
  XOR2_X1   g031(.A(KEYINPUT83), .B(G15gat), .Z(new_n233_));
  NAND2_X1  g032(.A1(G227gat), .A2(G233gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n232_), .B(new_n235_), .ZN(new_n236_));
  XOR2_X1   g035(.A(G127gat), .B(G134gat), .Z(new_n237_));
  XOR2_X1   g036(.A(G113gat), .B(G120gat), .Z(new_n238_));
  NOR2_X1   g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n237_), .A2(new_n238_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT84), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT85), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n241_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n243_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n240_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n246_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n248_), .A2(new_n239_), .A3(new_n244_), .ZN(new_n249_));
  AND2_X1   g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  XOR2_X1   g049(.A(new_n236_), .B(new_n250_), .Z(new_n251_));
  XNOR2_X1  g050(.A(G71gat), .B(G99gat), .ZN(new_n252_));
  INV_X1    g051(.A(G43gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n252_), .B(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(KEYINPUT30), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT31), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n251_), .B(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(G228gat), .ZN(new_n259_));
  INV_X1    g058(.A(G233gat), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT29), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G155gat), .A2(G162gat), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT86), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(KEYINPUT86), .A2(G155gat), .A3(G162gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(G155gat), .ZN(new_n268_));
  INV_X1    g067(.A(G162gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n267_), .A2(new_n270_), .ZN(new_n271_));
  OAI21_X1  g070(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT88), .ZN(new_n273_));
  NOR3_X1   g072(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n274_));
  INV_X1    g073(.A(G141gat), .ZN(new_n275_));
  INV_X1    g074(.A(G148gat), .ZN(new_n276_));
  OAI21_X1  g075(.A(KEYINPUT2), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT2), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n278_), .A2(G141gat), .A3(G148gat), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n274_), .B1(new_n277_), .B2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n273_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT89), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT89), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n273_), .A2(new_n280_), .A3(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n271_), .B1(new_n282_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  AOI22_X1  g085(.A1(new_n267_), .A2(KEYINPUT1), .B1(new_n268_), .B2(new_n269_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT87), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT1), .ZN(new_n289_));
  AND2_X1   g088(.A1(new_n265_), .A2(new_n266_), .ZN(new_n290_));
  AOI22_X1  g089(.A1(new_n287_), .A2(new_n288_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n270_), .B1(new_n290_), .B2(new_n289_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT87), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  XOR2_X1   g093(.A(G141gat), .B(G148gat), .Z(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n262_), .B1(new_n286_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT93), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G197gat), .B(G204gat), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  XOR2_X1   g101(.A(G211gat), .B(G218gat), .Z(new_n303_));
  NAND3_X1  g102(.A1(new_n302_), .A2(new_n303_), .A3(KEYINPUT21), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n304_), .A2(KEYINPUT92), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(KEYINPUT92), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(G204gat), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n308_), .A2(KEYINPUT91), .A3(G197gat), .ZN(new_n309_));
  OAI211_X1 g108(.A(KEYINPUT21), .B(new_n309_), .C1(new_n302_), .C2(KEYINPUT91), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT21), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n303_), .B1(new_n311_), .B2(new_n301_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n310_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n307_), .A2(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n314_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n261_), .B1(new_n300_), .B2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G78gat), .B(G106gat), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT90), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n297_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n261_), .ZN(new_n322_));
  OAI211_X1 g121(.A(new_n322_), .B(new_n314_), .C1(new_n297_), .C2(new_n319_), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n316_), .B(new_n318_), .C1(new_n321_), .C2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(KEYINPUT94), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n286_), .A2(new_n296_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(new_n262_), .ZN(new_n328_));
  XOR2_X1   g127(.A(G22gat), .B(G50gat), .Z(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT28), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n328_), .B(new_n330_), .ZN(new_n331_));
  AOI22_X1  g130(.A1(new_n305_), .A2(new_n306_), .B1(new_n310_), .B2(new_n312_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n326_), .A2(KEYINPUT29), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n332_), .B1(new_n333_), .B2(KEYINPUT93), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n322_), .B1(new_n334_), .B2(new_n299_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n321_), .A2(new_n323_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n317_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  AOI22_X1  g136(.A1(new_n325_), .A2(new_n331_), .B1(new_n324_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT94), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n337_), .A2(new_n324_), .A3(new_n339_), .A4(new_n331_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n338_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G8gat), .B(G36gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(KEYINPUT18), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G64gat), .B(G92gat), .ZN(new_n345_));
  XOR2_X1   g144(.A(new_n344_), .B(new_n345_), .Z(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT95), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G226gat), .A2(G233gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT19), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n214_), .A2(new_n210_), .ZN(new_n351_));
  AND3_X1   g150(.A1(new_n351_), .A2(new_n208_), .A3(new_n204_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n230_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n221_), .B1(G183gat), .B2(G190gat), .ZN(new_n354_));
  AOI22_X1  g153(.A1(new_n352_), .A2(new_n353_), .B1(new_n225_), .B2(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(KEYINPUT20), .B1(new_n332_), .B2(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n314_), .A2(new_n232_), .ZN(new_n357_));
  OAI211_X1 g156(.A(new_n348_), .B(new_n350_), .C1(new_n356_), .C2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n314_), .A2(new_n232_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n332_), .A2(new_n355_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n350_), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n359_), .A2(new_n360_), .A3(KEYINPUT20), .A4(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n358_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n352_), .A2(new_n353_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n225_), .A2(new_n354_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n314_), .A2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n332_), .A2(new_n231_), .A3(new_n222_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n367_), .A2(new_n368_), .A3(KEYINPUT20), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n348_), .B1(new_n369_), .B2(new_n350_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n347_), .B1(new_n363_), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT96), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n350_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT95), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n374_), .A2(new_n346_), .A3(new_n362_), .A4(new_n358_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n371_), .A2(new_n372_), .A3(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT27), .ZN(new_n377_));
  OAI211_X1 g176(.A(KEYINPUT96), .B(new_n347_), .C1(new_n363_), .C2(new_n370_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n376_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n367_), .A2(new_n368_), .A3(KEYINPUT20), .A4(new_n361_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT99), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  OR2_X1    g181(.A1(new_n380_), .A2(new_n381_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n360_), .A2(KEYINPUT20), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n332_), .B1(new_n231_), .B2(new_n222_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n350_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT98), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  OAI211_X1 g187(.A(KEYINPUT98), .B(new_n350_), .C1(new_n384_), .C2(new_n385_), .ZN(new_n389_));
  AOI22_X1  g188(.A1(new_n382_), .A2(new_n383_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  OAI211_X1 g189(.A(KEYINPUT27), .B(new_n375_), .C1(new_n390_), .C2(new_n346_), .ZN(new_n391_));
  AOI22_X1  g190(.A1(new_n286_), .A2(new_n296_), .B1(new_n247_), .B2(new_n249_), .ZN(new_n392_));
  OR2_X1    g191(.A1(new_n392_), .A2(KEYINPUT4), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n240_), .A2(new_n241_), .ZN(new_n394_));
  AND3_X1   g193(.A1(new_n286_), .A2(new_n296_), .A3(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(KEYINPUT4), .B1(new_n395_), .B2(new_n392_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G225gat), .A2(G233gat), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n393_), .A2(new_n396_), .A3(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G1gat), .B(G29gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n400_), .B(new_n401_), .ZN(new_n402_));
  XOR2_X1   g201(.A(G57gat), .B(G85gat), .Z(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n397_), .B1(new_n395_), .B2(new_n392_), .ZN(new_n405_));
  AND3_X1   g204(.A1(new_n399_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n404_), .B1(new_n399_), .B2(new_n405_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n379_), .A2(new_n391_), .A3(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n258_), .B1(new_n342_), .B2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n337_), .A2(new_n324_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n333_), .A2(KEYINPUT93), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n412_), .A2(new_n299_), .A3(new_n314_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n314_), .A2(new_n322_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n414_), .B1(new_n333_), .B2(KEYINPUT90), .ZN(new_n415_));
  AOI22_X1  g214(.A1(new_n413_), .A2(new_n261_), .B1(new_n320_), .B2(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n339_), .B1(new_n416_), .B2(new_n318_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n331_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n411_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(new_n340_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n398_), .B1(new_n393_), .B2(new_n396_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n286_), .A2(new_n296_), .A3(new_n394_), .ZN(new_n422_));
  OAI211_X1 g221(.A(new_n422_), .B(new_n398_), .C1(new_n327_), .C2(new_n250_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(new_n404_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n421_), .A2(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT33), .B1(new_n407_), .B2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n376_), .A2(new_n378_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT33), .ZN(new_n428_));
  AND2_X1   g227(.A1(new_n399_), .A2(new_n405_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n428_), .B1(new_n429_), .B2(new_n404_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n426_), .A2(new_n427_), .A3(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n346_), .A2(KEYINPUT32), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n374_), .A2(new_n362_), .A3(new_n358_), .A4(new_n432_), .ZN(new_n433_));
  OAI221_X1 g232(.A(new_n433_), .B1(new_n390_), .B2(new_n432_), .C1(new_n406_), .C2(new_n407_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n420_), .A2(new_n431_), .A3(new_n434_), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n379_), .A2(new_n391_), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n420_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n408_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n438_), .A2(new_n257_), .ZN(new_n439_));
  AOI22_X1  g238(.A1(new_n410_), .A2(new_n435_), .B1(new_n437_), .B2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G229gat), .A2(G233gat), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  XOR2_X1   g241(.A(G1gat), .B(G8gat), .Z(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(G1gat), .A2(G8gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT14), .ZN(new_n446_));
  INV_X1    g245(.A(G15gat), .ZN(new_n447_));
  INV_X1    g246(.A(G22gat), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(G15gat), .A2(G22gat), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n446_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n451_), .A2(KEYINPUT77), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n451_), .A2(KEYINPUT77), .ZN(new_n453_));
  NOR3_X1   g252(.A1(new_n452_), .A2(new_n453_), .A3(KEYINPUT78), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT78), .ZN(new_n455_));
  OR2_X1    g254(.A1(new_n451_), .A2(KEYINPUT77), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n451_), .A2(KEYINPUT77), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n455_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n444_), .B1(new_n454_), .B2(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT78), .B1(new_n452_), .B2(new_n453_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n456_), .A2(new_n455_), .A3(new_n457_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n460_), .A2(new_n461_), .A3(new_n443_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n459_), .A2(new_n462_), .ZN(new_n463_));
  XOR2_X1   g262(.A(G43gat), .B(G50gat), .Z(new_n464_));
  XNOR2_X1  g263(.A(G29gat), .B(G36gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n463_), .A2(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n466_), .B1(new_n459_), .B2(new_n462_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n442_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n469_), .ZN(new_n471_));
  XOR2_X1   g270(.A(new_n466_), .B(KEYINPUT15), .Z(new_n472_));
  NAND3_X1  g271(.A1(new_n472_), .A2(new_n462_), .A3(new_n459_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n471_), .A2(new_n441_), .A3(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n470_), .A2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G113gat), .B(G141gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G169gat), .B(G197gat), .ZN(new_n477_));
  XOR2_X1   g276(.A(new_n476_), .B(new_n477_), .Z(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n475_), .B(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT80), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n440_), .A2(new_n481_), .ZN(new_n482_));
  XOR2_X1   g281(.A(G190gat), .B(G218gat), .Z(new_n483_));
  XNOR2_X1  g282(.A(G134gat), .B(G162gat), .ZN(new_n484_));
  OR2_X1    g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n483_), .A2(new_n484_), .ZN(new_n486_));
  AOI21_X1  g285(.A(KEYINPUT36), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  XOR2_X1   g286(.A(new_n487_), .B(KEYINPUT75), .Z(new_n488_));
  NAND2_X1  g287(.A1(G232gat), .A2(G233gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT34), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(KEYINPUT35), .ZN(new_n491_));
  XOR2_X1   g290(.A(new_n491_), .B(KEYINPUT73), .Z(new_n492_));
  NAND2_X1  g291(.A1(G99gat), .A2(G106gat), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT65), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n494_), .A2(KEYINPUT6), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT6), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n496_), .A2(KEYINPUT65), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n493_), .B1(new_n495_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(KEYINPUT65), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n494_), .A2(KEYINPUT6), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n499_), .A2(new_n500_), .A3(G99gat), .A4(G106gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n498_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT66), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n498_), .A2(KEYINPUT66), .A3(new_n501_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(G99gat), .A2(G106gat), .ZN(new_n507_));
  AND2_X1   g306(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n508_));
  NOR2_X1   g307(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n507_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  OAI22_X1  g309(.A1(KEYINPUT67), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n506_), .A2(new_n513_), .ZN(new_n514_));
  XOR2_X1   g313(.A(G85gat), .B(G92gat), .Z(new_n515_));
  INV_X1    g314(.A(KEYINPUT8), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n514_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT68), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n512_), .A2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n510_), .A2(KEYINPUT68), .A3(new_n511_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n521_), .A2(new_n522_), .A3(new_n502_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n523_), .A2(KEYINPUT69), .A3(new_n515_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT8), .ZN(new_n525_));
  AOI21_X1  g324(.A(KEYINPUT69), .B1(new_n523_), .B2(new_n515_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n519_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  AND2_X1   g326(.A1(new_n515_), .A2(KEYINPUT9), .ZN(new_n528_));
  XNOR2_X1  g327(.A(KEYINPUT10), .B(G99gat), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n529_), .A2(G106gat), .ZN(new_n530_));
  INV_X1    g329(.A(G85gat), .ZN(new_n531_));
  INV_X1    g330(.A(G92gat), .ZN(new_n532_));
  NOR3_X1   g331(.A1(new_n531_), .A2(new_n532_), .A3(KEYINPUT9), .ZN(new_n533_));
  NOR3_X1   g332(.A1(new_n528_), .A2(new_n530_), .A3(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n506_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n527_), .A2(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(KEYINPUT74), .B1(new_n536_), .B2(new_n466_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n535_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n523_), .A2(new_n515_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT69), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n541_), .A2(KEYINPUT8), .A3(new_n524_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n538_), .B1(new_n542_), .B2(new_n519_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT74), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n543_), .A2(new_n544_), .A3(new_n467_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n537_), .A2(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n490_), .A2(KEYINPUT35), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n506_), .A2(new_n534_), .A3(KEYINPUT71), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(KEYINPUT71), .B1(new_n506_), .B2(new_n534_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n527_), .A2(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n547_), .B1(new_n552_), .B2(new_n472_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n492_), .B1(new_n546_), .B2(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n544_), .B1(new_n543_), .B2(new_n467_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n517_), .B1(new_n506_), .B2(new_n513_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n515_), .ZN(new_n557_));
  AOI22_X1  g356(.A1(new_n512_), .A2(new_n520_), .B1(new_n498_), .B2(new_n501_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n557_), .B1(new_n558_), .B2(new_n522_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n516_), .B1(new_n559_), .B2(KEYINPUT69), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n556_), .B1(new_n560_), .B2(new_n541_), .ZN(new_n561_));
  NOR4_X1   g360(.A1(new_n561_), .A2(KEYINPUT74), .A3(new_n466_), .A4(new_n538_), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n553_), .B(new_n492_), .C1(new_n555_), .C2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n488_), .B1(new_n554_), .B2(new_n564_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n553_), .B1(new_n555_), .B2(new_n562_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n492_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n485_), .A2(new_n486_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT36), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT76), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n568_), .A2(new_n563_), .A3(new_n571_), .ZN(new_n572_));
  AND3_X1   g371(.A1(new_n565_), .A2(KEYINPUT37), .A3(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n568_), .A2(new_n563_), .A3(new_n570_), .ZN(new_n574_));
  AOI21_X1  g373(.A(KEYINPUT37), .B1(new_n565_), .B2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G57gat), .B(G64gat), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(KEYINPUT11), .ZN(new_n577_));
  XOR2_X1   g376(.A(G71gat), .B(G78gat), .Z(new_n578_));
  OR2_X1    g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n576_), .A2(KEYINPUT11), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n577_), .A2(new_n578_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n579_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G231gat), .A2(G233gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n463_), .B(new_n584_), .ZN(new_n585_));
  XOR2_X1   g384(.A(G127gat), .B(G155gat), .Z(new_n586_));
  XNOR2_X1  g385(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G183gat), .B(G211gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n585_), .A2(KEYINPUT17), .A3(new_n591_), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n590_), .B(KEYINPUT17), .Z(new_n593_));
  OAI21_X1  g392(.A(new_n592_), .B1(new_n585_), .B2(new_n593_), .ZN(new_n594_));
  NOR3_X1   g393(.A1(new_n573_), .A2(new_n575_), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT13), .ZN(new_n597_));
  NAND2_X1  g396(.A1(G230gat), .A2(G233gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT64), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT70), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n527_), .A2(new_n601_), .A3(new_n535_), .A4(new_n582_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n602_), .B1(new_n543_), .B2(new_n582_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n601_), .B1(new_n543_), .B2(new_n582_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n600_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT12), .ZN(new_n606_));
  OR2_X1    g405(.A1(new_n582_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  AOI22_X1  g407(.A1(new_n552_), .A2(new_n608_), .B1(new_n543_), .B2(new_n582_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n606_), .B1(new_n543_), .B2(new_n582_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n609_), .A2(new_n599_), .A3(new_n610_), .ZN(new_n611_));
  XOR2_X1   g410(.A(G120gat), .B(G148gat), .Z(new_n612_));
  XNOR2_X1  g411(.A(G176gat), .B(G204gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n614_), .B(new_n615_), .Z(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  AND3_X1   g416(.A1(new_n605_), .A2(new_n611_), .A3(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n617_), .B1(new_n605_), .B2(new_n611_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n597_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n605_), .A2(new_n611_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(new_n616_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n605_), .A2(new_n611_), .A3(new_n617_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n622_), .A2(KEYINPUT13), .A3(new_n623_), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n620_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n596_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n482_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT100), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n482_), .A2(KEYINPUT100), .A3(new_n627_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(G1gat), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n632_), .A2(KEYINPUT38), .A3(new_n633_), .A4(new_n438_), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n634_), .A2(KEYINPUT101), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n632_), .A2(new_n633_), .A3(new_n438_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n565_), .A2(new_n574_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT103), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n565_), .A2(KEYINPUT103), .A3(new_n574_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n409_), .A2(new_n340_), .A3(new_n419_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n435_), .A2(new_n642_), .A3(new_n257_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n420_), .A2(new_n436_), .A3(new_n439_), .ZN(new_n644_));
  AOI211_X1 g443(.A(new_n594_), .B(new_n641_), .C1(new_n643_), .C2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n625_), .A2(new_n480_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(KEYINPUT102), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n646_), .A2(KEYINPUT102), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n645_), .A2(new_n647_), .A3(new_n648_), .ZN(new_n649_));
  OAI21_X1  g448(.A(G1gat), .B1(new_n649_), .B2(new_n408_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(KEYINPUT38), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n636_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n634_), .A2(KEYINPUT101), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n635_), .A2(new_n652_), .A3(new_n653_), .ZN(G1324gat));
  OAI21_X1  g453(.A(G8gat), .B1(new_n649_), .B2(new_n436_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT39), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n436_), .A2(G8gat), .ZN(new_n657_));
  AOI21_X1  g456(.A(KEYINPUT104), .B1(new_n632_), .B2(new_n657_), .ZN(new_n658_));
  AND4_X1   g457(.A1(KEYINPUT104), .A2(new_n630_), .A3(new_n631_), .A4(new_n657_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n656_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT40), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  OAI211_X1 g461(.A(new_n656_), .B(KEYINPUT40), .C1(new_n658_), .C2(new_n659_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1325gat));
  NAND3_X1  g463(.A1(new_n632_), .A2(new_n447_), .A3(new_n258_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT105), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n665_), .B(new_n666_), .ZN(new_n667_));
  OAI21_X1  g466(.A(G15gat), .B1(new_n649_), .B2(new_n257_), .ZN(new_n668_));
  XOR2_X1   g467(.A(new_n668_), .B(KEYINPUT41), .Z(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(G1326gat));
  OAI21_X1  g469(.A(G22gat), .B1(new_n649_), .B2(new_n420_), .ZN(new_n671_));
  XOR2_X1   g470(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n672_));
  XNOR2_X1  g471(.A(new_n671_), .B(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n342_), .A2(new_n448_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT107), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n632_), .A2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n673_), .A2(new_n676_), .ZN(G1327gat));
  INV_X1    g476(.A(new_n641_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n594_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n678_), .A2(new_n626_), .A3(new_n679_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n482_), .A2(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(G29gat), .B1(new_n681_), .B2(new_n438_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT43), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT37), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n568_), .A2(new_n563_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n685_), .B2(new_n488_), .ZN(new_n686_));
  AOI22_X1  g485(.A1(new_n637_), .A2(new_n684_), .B1(new_n686_), .B2(new_n572_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n687_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n683_), .B1(new_n688_), .B2(KEYINPUT108), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT108), .ZN(new_n690_));
  OAI211_X1 g489(.A(new_n690_), .B(KEYINPUT43), .C1(new_n440_), .C2(new_n687_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n648_), .A2(new_n594_), .A3(new_n647_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n692_), .A2(KEYINPUT44), .A3(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(KEYINPUT109), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n693_), .B1(new_n689_), .B2(new_n691_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT109), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n697_), .A2(new_n698_), .A3(KEYINPUT44), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n696_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n697_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n700_), .A2(new_n703_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n438_), .A2(G29gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n682_), .B1(new_n704_), .B2(new_n705_), .ZN(G1328gat));
  INV_X1    g505(.A(KEYINPUT46), .ZN(new_n707_));
  INV_X1    g506(.A(G36gat), .ZN(new_n708_));
  INV_X1    g507(.A(new_n436_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n709_), .B1(new_n697_), .B2(KEYINPUT44), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n708_), .B1(new_n700_), .B2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT45), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT111), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n436_), .B(KEYINPUT110), .Z(new_n715_));
  NOR2_X1   g514(.A1(new_n715_), .A2(G36gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n714_), .B1(new_n681_), .B2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n482_), .A2(new_n680_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n716_), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n718_), .A2(KEYINPUT111), .A3(new_n719_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n713_), .B1(new_n717_), .B2(new_n720_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n681_), .A2(new_n714_), .A3(new_n716_), .ZN(new_n722_));
  OAI21_X1  g521(.A(KEYINPUT111), .B1(new_n718_), .B2(new_n719_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n722_), .A2(KEYINPUT45), .A3(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n721_), .A2(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n707_), .B1(new_n712_), .B2(new_n725_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n721_), .A2(new_n724_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n710_), .B1(new_n696_), .B2(new_n699_), .ZN(new_n728_));
  OAI211_X1 g527(.A(new_n727_), .B(KEYINPUT46), .C1(new_n708_), .C2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n726_), .A2(new_n729_), .ZN(G1329gat));
  NOR2_X1   g529(.A1(new_n257_), .A2(new_n253_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n695_), .A2(KEYINPUT109), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n698_), .B1(new_n697_), .B2(KEYINPUT44), .ZN(new_n733_));
  OAI211_X1 g532(.A(new_n703_), .B(new_n731_), .C1(new_n732_), .C2(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n253_), .B1(new_n718_), .B2(new_n257_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n734_), .A2(new_n735_), .A3(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n737_), .A2(new_n738_), .ZN(G1330gat));
  AOI21_X1  g538(.A(G50gat), .B1(new_n681_), .B2(new_n342_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n342_), .A2(G50gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n704_), .B2(new_n741_), .ZN(G1331gat));
  AND3_X1   g541(.A1(new_n645_), .A2(new_n481_), .A3(new_n626_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n743_), .A2(G57gat), .A3(new_n438_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT114), .ZN(new_n745_));
  INV_X1    g544(.A(G57gat), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n440_), .A2(new_n480_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n596_), .A2(new_n625_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n408_), .B1(new_n749_), .B2(KEYINPUT113), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n750_), .B1(KEYINPUT113), .B2(new_n749_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n745_), .B1(new_n746_), .B2(new_n751_), .ZN(G1332gat));
  OR3_X1    g551(.A1(new_n749_), .A2(G64gat), .A3(new_n715_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n715_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n743_), .A2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT48), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n755_), .A2(new_n756_), .A3(G64gat), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n755_), .B2(G64gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n753_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT115), .ZN(G1333gat));
  INV_X1    g559(.A(G71gat), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n761_), .B1(new_n743_), .B2(new_n258_), .ZN(new_n762_));
  XOR2_X1   g561(.A(new_n762_), .B(KEYINPUT49), .Z(new_n763_));
  INV_X1    g562(.A(new_n749_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n764_), .A2(new_n761_), .A3(new_n258_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n763_), .A2(new_n765_), .ZN(G1334gat));
  INV_X1    g565(.A(G78gat), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n767_), .B1(new_n743_), .B2(new_n342_), .ZN(new_n768_));
  XOR2_X1   g567(.A(new_n768_), .B(KEYINPUT50), .Z(new_n769_));
  NAND3_X1  g568(.A1(new_n764_), .A2(new_n767_), .A3(new_n342_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(G1335gat));
  NAND4_X1  g570(.A1(new_n747_), .A2(new_n626_), .A3(new_n594_), .A4(new_n641_), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n772_), .A2(G85gat), .A3(new_n408_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n480_), .A2(new_n679_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n626_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT116), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n775_), .B(new_n776_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n692_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(new_n438_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n773_), .B1(new_n779_), .B2(G85gat), .ZN(new_n780_));
  XOR2_X1   g579(.A(new_n780_), .B(KEYINPUT117), .Z(G1336gat));
  OAI21_X1  g580(.A(new_n532_), .B1(new_n772_), .B2(new_n436_), .ZN(new_n782_));
  XOR2_X1   g581(.A(new_n782_), .B(KEYINPUT118), .Z(new_n783_));
  NOR2_X1   g582(.A1(new_n715_), .A2(new_n532_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n783_), .B1(new_n778_), .B2(new_n784_), .ZN(G1337gat));
  NOR3_X1   g584(.A1(new_n772_), .A2(new_n257_), .A3(new_n529_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n778_), .A2(new_n258_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n787_), .B2(G99gat), .ZN(new_n788_));
  XOR2_X1   g587(.A(new_n788_), .B(KEYINPUT51), .Z(G1338gat));
  NOR3_X1   g588(.A1(new_n772_), .A2(G106gat), .A3(new_n420_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n692_), .A2(new_n342_), .A3(new_n777_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(G106gat), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT52), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT52), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n791_), .A2(new_n794_), .A3(G106gat), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n790_), .B1(new_n793_), .B2(new_n795_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(KEYINPUT119), .B(KEYINPUT53), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n797_), .ZN(new_n799_));
  AOI211_X1 g598(.A(new_n790_), .B(new_n799_), .C1(new_n793_), .C2(new_n795_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n798_), .A2(new_n800_), .ZN(G1339gat));
  NAND4_X1  g600(.A1(new_n687_), .A2(new_n625_), .A3(new_n481_), .A4(new_n679_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT120), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n595_), .A2(KEYINPUT120), .A3(new_n481_), .A4(new_n625_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n804_), .A2(KEYINPUT54), .A3(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT54), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n802_), .A2(new_n803_), .A3(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n480_), .A2(new_n623_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n812_));
  INV_X1    g611(.A(new_n550_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n548_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n608_), .B1(new_n561_), .B2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n527_), .A2(new_n535_), .A3(new_n582_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n582_), .B1(new_n527_), .B2(new_n535_), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n815_), .B(new_n816_), .C1(new_n817_), .C2(KEYINPUT12), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n812_), .B1(new_n818_), .B2(new_n600_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n600_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n609_), .A2(KEYINPUT55), .A3(new_n599_), .A4(new_n610_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n819_), .A2(new_n820_), .A3(new_n821_), .ZN(new_n822_));
  AND3_X1   g621(.A1(new_n822_), .A2(KEYINPUT56), .A3(new_n616_), .ZN(new_n823_));
  AOI21_X1  g622(.A(KEYINPUT56), .B1(new_n822_), .B2(new_n616_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n811_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT121), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT121), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n811_), .B(new_n827_), .C1(new_n823_), .C2(new_n824_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n622_), .A2(new_n623_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n475_), .A2(new_n479_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n441_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n479_), .ZN(new_n832_));
  OR2_X1    g631(.A1(new_n832_), .A2(KEYINPUT122), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n469_), .A2(new_n441_), .ZN(new_n834_));
  AOI22_X1  g633(.A1(new_n832_), .A2(KEYINPUT122), .B1(new_n473_), .B2(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n830_), .B1(new_n833_), .B2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n829_), .A2(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n826_), .A2(new_n828_), .A3(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT57), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n641_), .A2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n840_), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n836_), .A2(new_n623_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n842_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT58), .ZN(new_n844_));
  OR2_X1    g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n575_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n686_), .A2(new_n572_), .ZN(new_n847_));
  AOI22_X1  g646(.A1(new_n843_), .A2(new_n844_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n845_), .A2(new_n848_), .ZN(new_n849_));
  AOI22_X1  g648(.A1(new_n825_), .A2(KEYINPUT121), .B1(new_n829_), .B2(new_n836_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n641_), .B1(new_n850_), .B2(new_n828_), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n841_), .B(new_n849_), .C1(new_n851_), .C2(KEYINPUT57), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n809_), .B1(new_n594_), .B2(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n437_), .A2(new_n438_), .A3(new_n258_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(G113gat), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n855_), .A2(new_n856_), .A3(new_n480_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT59), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n858_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n854_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n822_), .A2(new_n616_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT56), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n822_), .A2(KEYINPUT56), .A3(new_n616_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n810_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n837_), .B1(new_n865_), .B2(new_n827_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n828_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n678_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n839_), .ZN(new_n869_));
  AOI22_X1  g668(.A1(new_n838_), .A2(new_n840_), .B1(new_n845_), .B2(new_n848_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n679_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  OAI211_X1 g670(.A(KEYINPUT59), .B(new_n860_), .C1(new_n871_), .C2(new_n809_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n481_), .B1(new_n859_), .B2(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n857_), .B1(new_n873_), .B2(new_n856_), .ZN(G1340gat));
  NOR2_X1   g673(.A1(new_n625_), .A2(KEYINPUT60), .ZN(new_n875_));
  MUX2_X1   g674(.A(new_n875_), .B(KEYINPUT60), .S(G120gat), .Z(new_n876_));
  NAND2_X1  g675(.A1(new_n855_), .A2(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n625_), .B1(new_n859_), .B2(new_n872_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT123), .ZN(new_n879_));
  OAI21_X1  g678(.A(G120gat), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  AOI211_X1 g679(.A(KEYINPUT123), .B(new_n625_), .C1(new_n859_), .C2(new_n872_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n877_), .B1(new_n880_), .B2(new_n881_), .ZN(G1341gat));
  INV_X1    g681(.A(G127gat), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n855_), .A2(new_n883_), .A3(new_n679_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n594_), .B1(new_n859_), .B2(new_n872_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n885_), .B2(new_n883_), .ZN(G1342gat));
  INV_X1    g685(.A(G134gat), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n855_), .A2(new_n887_), .A3(new_n641_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n687_), .B1(new_n859_), .B2(new_n872_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n889_), .B2(new_n887_), .ZN(G1343gat));
  NAND3_X1  g689(.A1(new_n342_), .A2(new_n438_), .A3(new_n257_), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n853_), .A2(new_n754_), .A3(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n480_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n626_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g695(.A1(new_n892_), .A2(new_n679_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(KEYINPUT61), .B(G155gat), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n897_), .B(new_n898_), .ZN(G1346gat));
  NAND3_X1  g698(.A1(new_n892_), .A2(new_n269_), .A3(new_n641_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n687_), .ZN(new_n901_));
  AND2_X1   g700(.A1(new_n892_), .A2(new_n901_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n900_), .B1(new_n902_), .B2(new_n269_), .ZN(G1347gat));
  INV_X1    g702(.A(KEYINPUT62), .ZN(new_n904_));
  INV_X1    g703(.A(new_n853_), .ZN(new_n905_));
  NOR4_X1   g704(.A1(new_n715_), .A2(new_n342_), .A3(new_n438_), .A4(new_n257_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n480_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n907_), .A2(new_n908_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n904_), .B1(new_n909_), .B2(new_n205_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n223_), .ZN(new_n911_));
  OAI211_X1 g710(.A(KEYINPUT62), .B(G169gat), .C1(new_n907_), .C2(new_n908_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n910_), .A2(new_n911_), .A3(new_n912_), .ZN(G1348gat));
  NOR2_X1   g712(.A1(new_n907_), .A2(new_n625_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(new_n206_), .ZN(G1349gat));
  NAND3_X1  g714(.A1(new_n905_), .A2(new_n679_), .A3(new_n906_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n916_), .A2(new_n202_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n917_), .B1(new_n216_), .B2(new_n916_), .ZN(G1350gat));
  NAND4_X1  g717(.A1(new_n905_), .A2(new_n203_), .A3(new_n641_), .A4(new_n906_), .ZN(new_n919_));
  OAI211_X1 g718(.A(new_n901_), .B(new_n906_), .C1(new_n871_), .C2(new_n809_), .ZN(new_n920_));
  AND3_X1   g719(.A1(new_n920_), .A2(KEYINPUT124), .A3(G190gat), .ZN(new_n921_));
  AOI21_X1  g720(.A(KEYINPUT124), .B1(new_n920_), .B2(G190gat), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n919_), .B1(new_n921_), .B2(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(KEYINPUT125), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT125), .ZN(new_n925_));
  OAI211_X1 g724(.A(new_n925_), .B(new_n919_), .C1(new_n921_), .C2(new_n922_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n924_), .A2(new_n926_), .ZN(G1351gat));
  NAND3_X1  g726(.A1(new_n342_), .A2(new_n408_), .A3(new_n257_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n754_), .B1(KEYINPUT126), .B2(new_n928_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n929_), .B1(KEYINPUT126), .B2(new_n928_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n905_), .A2(new_n930_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n931_), .A2(new_n908_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(KEYINPUT127), .B(G197gat), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n932_), .B(new_n933_), .ZN(G1352gat));
  NOR2_X1   g733(.A1(new_n931_), .A2(new_n625_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(new_n308_), .ZN(G1353gat));
  NOR2_X1   g735(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n937_), .B1(new_n931_), .B2(new_n594_), .ZN(new_n938_));
  XOR2_X1   g737(.A(KEYINPUT63), .B(G211gat), .Z(new_n939_));
  NAND4_X1  g738(.A1(new_n905_), .A2(new_n679_), .A3(new_n930_), .A4(new_n939_), .ZN(new_n940_));
  AND2_X1   g739(.A1(new_n938_), .A2(new_n940_), .ZN(G1354gat));
  OAI21_X1  g740(.A(G218gat), .B1(new_n931_), .B2(new_n687_), .ZN(new_n942_));
  OR2_X1    g741(.A1(new_n678_), .A2(G218gat), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n942_), .B1(new_n931_), .B2(new_n943_), .ZN(G1355gat));
endmodule


