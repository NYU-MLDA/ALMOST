//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1 0 1 0 1 0 0 1 1 0 1 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n656_, new_n657_,
    new_n658_, new_n660_, new_n661_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n682_, new_n683_, new_n684_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n694_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n807_,
    new_n808_, new_n809_, new_n811_, new_n812_, new_n813_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n824_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n877_, new_n878_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n892_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_;
  XNOR2_X1  g000(.A(G22gat), .B(G50gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT86), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n206_), .B1(G155gat), .B2(G162gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT87), .ZN(new_n208_));
  AND2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n207_), .A2(new_n208_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G141gat), .A2(G148gat), .ZN(new_n211_));
  XOR2_X1   g010(.A(new_n211_), .B(KEYINPUT2), .Z(new_n212_));
  NOR2_X1   g011(.A1(G141gat), .A2(G148gat), .ZN(new_n213_));
  XOR2_X1   g012(.A(new_n213_), .B(KEYINPUT3), .Z(new_n214_));
  OAI22_X1  g013(.A1(new_n209_), .A2(new_n210_), .B1(new_n212_), .B2(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n216_), .B1(new_n206_), .B2(KEYINPUT1), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n217_), .B1(KEYINPUT1), .B2(new_n206_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n213_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n218_), .A2(new_n211_), .A3(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n215_), .A2(new_n220_), .ZN(new_n221_));
  NOR3_X1   g020(.A1(new_n221_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT28), .B1(new_n221_), .B2(KEYINPUT29), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n203_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n223_), .A2(new_n224_), .A3(new_n203_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G78gat), .B(G106gat), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n226_), .A2(new_n227_), .A3(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n224_), .ZN(new_n231_));
  NOR3_X1   g030(.A1(new_n231_), .A2(new_n222_), .A3(new_n202_), .ZN(new_n232_));
  OAI211_X1 g031(.A(KEYINPUT90), .B(new_n228_), .C1(new_n232_), .C2(new_n225_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n230_), .A2(new_n233_), .ZN(new_n234_));
  XOR2_X1   g033(.A(G197gat), .B(G204gat), .Z(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(KEYINPUT21), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G211gat), .B(G218gat), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT89), .ZN(new_n239_));
  INV_X1    g038(.A(new_n235_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT21), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n240_), .A2(KEYINPUT88), .A3(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(KEYINPUT88), .B1(new_n240_), .B2(new_n241_), .ZN(new_n244_));
  OAI211_X1 g043(.A(new_n236_), .B(new_n237_), .C1(new_n243_), .C2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n239_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n247_), .B1(KEYINPUT29), .B2(new_n221_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G228gat), .A2(G233gat), .ZN(new_n249_));
  XOR2_X1   g048(.A(new_n248_), .B(new_n249_), .Z(new_n250_));
  NAND2_X1  g049(.A1(new_n234_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n250_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n252_), .A2(new_n230_), .A3(new_n233_), .ZN(new_n253_));
  AND2_X1   g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G1gat), .B(G29gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(G85gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT0), .B(G57gat), .ZN(new_n257_));
  XOR2_X1   g056(.A(new_n256_), .B(new_n257_), .Z(new_n258_));
  XNOR2_X1  g057(.A(G127gat), .B(G134gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G113gat), .B(G120gat), .ZN(new_n260_));
  XOR2_X1   g059(.A(new_n259_), .B(new_n260_), .Z(new_n261_));
  OR2_X1    g060(.A1(new_n221_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n221_), .A2(new_n261_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G225gat), .A2(G233gat), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n262_), .A2(KEYINPUT4), .A3(new_n263_), .ZN(new_n269_));
  OR2_X1    g068(.A1(new_n263_), .A2(KEYINPUT4), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n266_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n258_), .B1(new_n268_), .B2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT33), .ZN(new_n273_));
  OR2_X1    g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n273_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G183gat), .A2(G190gat), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT23), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(G183gat), .A2(G190gat), .ZN(new_n279_));
  OR2_X1    g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G169gat), .A2(G176gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT22), .B(G169gat), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  AND2_X1   g082(.A1(new_n283_), .A2(KEYINPUT83), .ZN(new_n284_));
  XNOR2_X1  g083(.A(KEYINPUT84), .B(G176gat), .ZN(new_n285_));
  INV_X1    g084(.A(G169gat), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n286_), .A2(KEYINPUT22), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n285_), .B1(KEYINPUT83), .B2(new_n287_), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n280_), .B(new_n281_), .C1(new_n284_), .C2(new_n288_), .ZN(new_n289_));
  OR2_X1    g088(.A1(G169gat), .A2(G176gat), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n290_), .A2(KEYINPUT24), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n278_), .A2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT25), .B(G183gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT26), .B(G190gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n290_), .A2(KEYINPUT24), .A3(new_n281_), .ZN(new_n296_));
  AND2_X1   g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n292_), .B1(new_n297_), .B2(KEYINPUT82), .ZN(new_n298_));
  AND3_X1   g097(.A1(new_n295_), .A2(KEYINPUT82), .A3(new_n296_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n289_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  OR2_X1    g099(.A1(new_n246_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT20), .ZN(new_n302_));
  INV_X1    g101(.A(new_n285_), .ZN(new_n303_));
  OAI211_X1 g102(.A(new_n280_), .B(new_n281_), .C1(new_n283_), .C2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n297_), .A2(new_n292_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n302_), .B1(new_n246_), .B2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n301_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G226gat), .A2(G233gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT19), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n306_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n302_), .B1(new_n247_), .B2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n310_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n246_), .A2(new_n300_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n313_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n311_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G8gat), .B(G36gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT18), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G64gat), .B(G92gat), .ZN(new_n320_));
  XOR2_X1   g119(.A(new_n319_), .B(new_n320_), .Z(new_n321_));
  XNOR2_X1  g120(.A(new_n317_), .B(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n258_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n269_), .A2(new_n270_), .ZN(new_n324_));
  AND2_X1   g123(.A1(new_n264_), .A2(KEYINPUT91), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n267_), .B1(new_n264_), .B2(KEYINPUT91), .ZN(new_n326_));
  OAI221_X1 g125(.A(new_n323_), .B1(new_n324_), .B2(new_n267_), .C1(new_n325_), .C2(new_n326_), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n274_), .A2(new_n275_), .A3(new_n322_), .A4(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n324_), .A2(new_n267_), .ZN(new_n329_));
  OAI211_X1 g128(.A(new_n329_), .B(new_n323_), .C1(new_n267_), .C2(new_n265_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT92), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n330_), .A2(new_n331_), .A3(new_n272_), .ZN(new_n332_));
  OAI211_X1 g131(.A(KEYINPUT92), .B(new_n258_), .C1(new_n268_), .C2(new_n271_), .ZN(new_n333_));
  AND2_X1   g132(.A1(new_n321_), .A2(KEYINPUT32), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n317_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n313_), .A2(new_n315_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(new_n310_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n337_), .B1(new_n310_), .B2(new_n308_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n335_), .B1(new_n338_), .B2(new_n334_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n332_), .A2(new_n333_), .A3(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n254_), .A2(new_n328_), .A3(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G71gat), .B(G99gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(G43gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n300_), .B(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G227gat), .A2(G233gat), .ZN(new_n345_));
  INV_X1    g144(.A(G15gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT30), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n344_), .B(new_n348_), .ZN(new_n349_));
  OR2_X1    g148(.A1(new_n349_), .A2(KEYINPUT85), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(KEYINPUT85), .ZN(new_n351_));
  XOR2_X1   g150(.A(new_n261_), .B(KEYINPUT31), .Z(new_n352_));
  NAND3_X1  g151(.A1(new_n350_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n352_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n349_), .A2(KEYINPUT85), .A3(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n353_), .A2(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n311_), .A2(new_n321_), .A3(new_n316_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT93), .ZN(new_n358_));
  OR2_X1    g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n321_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n338_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n357_), .A2(new_n358_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n359_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(KEYINPUT27), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT27), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n322_), .A2(new_n365_), .ZN(new_n366_));
  AOI22_X1  g165(.A1(new_n364_), .A2(new_n366_), .B1(new_n333_), .B2(new_n332_), .ZN(new_n367_));
  OAI211_X1 g166(.A(new_n341_), .B(new_n356_), .C1(new_n367_), .C2(new_n254_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n356_), .B1(new_n333_), .B2(new_n332_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n364_), .A2(new_n366_), .ZN(new_n370_));
  AND4_X1   g169(.A1(KEYINPUT94), .A2(new_n369_), .A3(new_n254_), .A4(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n251_), .A2(new_n253_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n372_), .B1(new_n364_), .B2(new_n366_), .ZN(new_n373_));
  AOI21_X1  g172(.A(KEYINPUT94), .B1(new_n373_), .B2(new_n369_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n368_), .B1(new_n371_), .B2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G15gat), .B(G22gat), .ZN(new_n376_));
  INV_X1    g175(.A(G1gat), .ZN(new_n377_));
  INV_X1    g176(.A(G8gat), .ZN(new_n378_));
  OAI21_X1  g177(.A(KEYINPUT14), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n376_), .A2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G1gat), .B(G8gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(G36gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(G29gat), .ZN(new_n384_));
  INV_X1    g183(.A(G29gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(G36gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(G50gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(G43gat), .ZN(new_n389_));
  INV_X1    g188(.A(G43gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(G50gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n387_), .A2(new_n392_), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n384_), .A2(new_n386_), .A3(new_n389_), .A4(new_n391_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  XOR2_X1   g194(.A(new_n382_), .B(new_n395_), .Z(new_n396_));
  NAND3_X1  g195(.A1(new_n396_), .A2(G229gat), .A3(G233gat), .ZN(new_n397_));
  INV_X1    g196(.A(new_n382_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(new_n395_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT69), .B(KEYINPUT15), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n393_), .A2(new_n394_), .A3(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n400_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(new_n382_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G229gat), .A2(G233gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(KEYINPUT80), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n399_), .A2(new_n404_), .A3(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G113gat), .B(G141gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT81), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G169gat), .B(G197gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n397_), .A2(new_n407_), .A3(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n411_), .B1(new_n397_), .B2(new_n407_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  AND2_X1   g215(.A1(new_n375_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT73), .ZN(new_n418_));
  INV_X1    g217(.A(G85gat), .ZN(new_n419_));
  INV_X1    g218(.A(G92gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT65), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT8), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G85gat), .A2(G92gat), .ZN(new_n424_));
  AND3_X1   g223(.A1(new_n421_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G99gat), .A2(G106gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT6), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT6), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n428_), .A2(G99gat), .A3(G106gat), .ZN(new_n429_));
  AND2_X1   g228(.A1(new_n427_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT7), .ZN(new_n431_));
  INV_X1    g230(.A(G99gat), .ZN(new_n432_));
  INV_X1    g231(.A(G106gat), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n431_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n425_), .B1(new_n430_), .B2(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n422_), .A2(KEYINPUT8), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  OAI221_X1 g238(.A(new_n425_), .B1(new_n422_), .B2(KEYINPUT8), .C1(new_n430_), .C2(new_n436_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n427_), .A2(new_n429_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(KEYINPUT10), .B(G99gat), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n442_), .B1(new_n443_), .B2(G106gat), .ZN(new_n444_));
  AND2_X1   g243(.A1(G85gat), .A2(G92gat), .ZN(new_n445_));
  NOR2_X1   g244(.A1(G85gat), .A2(G92gat), .ZN(new_n446_));
  OAI22_X1  g245(.A1(new_n445_), .A2(new_n446_), .B1(KEYINPUT9), .B2(new_n420_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT9), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n421_), .A2(new_n448_), .A3(new_n424_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT64), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n447_), .A2(new_n449_), .A3(KEYINPUT64), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n444_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n403_), .B1(new_n441_), .B2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(KEYINPUT68), .B(KEYINPUT34), .ZN(new_n456_));
  AND2_X1   g255(.A1(G232gat), .A2(G233gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT35), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n458_), .A2(new_n459_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n444_), .ZN(new_n463_));
  AND3_X1   g262(.A1(new_n447_), .A2(new_n449_), .A3(KEYINPUT64), .ZN(new_n464_));
  AOI21_X1  g263(.A(KEYINPUT64), .B1(new_n447_), .B2(new_n449_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n463_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n466_), .A2(new_n395_), .A3(new_n439_), .A4(new_n440_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n455_), .A2(new_n461_), .A3(new_n462_), .A4(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(KEYINPUT72), .ZN(new_n469_));
  AND2_X1   g268(.A1(new_n467_), .A2(new_n462_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT72), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n466_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n460_), .B1(new_n472_), .B2(new_n403_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n470_), .A2(new_n471_), .A3(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n469_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n455_), .A2(KEYINPUT70), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT70), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n472_), .A2(new_n477_), .A3(new_n403_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n476_), .A2(new_n470_), .A3(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(new_n460_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n475_), .A2(new_n480_), .ZN(new_n481_));
  XOR2_X1   g280(.A(G190gat), .B(G218gat), .Z(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT71), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G134gat), .B(G162gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT36), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n418_), .B1(new_n481_), .B2(new_n487_), .ZN(new_n488_));
  AOI22_X1  g287(.A1(new_n469_), .A2(new_n474_), .B1(new_n479_), .B2(new_n460_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n487_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n489_), .A2(KEYINPUT73), .A3(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n488_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n485_), .B(new_n486_), .ZN(new_n493_));
  XOR2_X1   g292(.A(new_n493_), .B(KEYINPUT74), .Z(new_n494_));
  OAI21_X1  g293(.A(new_n492_), .B1(new_n489_), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(KEYINPUT37), .ZN(new_n496_));
  OAI21_X1  g295(.A(KEYINPUT75), .B1(new_n489_), .B2(new_n493_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT75), .ZN(new_n498_));
  INV_X1    g297(.A(new_n493_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n481_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n497_), .A2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(KEYINPUT76), .B(KEYINPUT37), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n492_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n496_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G231gat), .A2(G233gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n382_), .B(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(KEYINPUT66), .B(G71gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(G78gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G57gat), .B(G64gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT11), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n509_), .A2(KEYINPUT11), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n508_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(G78gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n507_), .B(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(new_n510_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n513_), .A2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n506_), .B(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT78), .ZN(new_n519_));
  XOR2_X1   g318(.A(G127gat), .B(G155gat), .Z(new_n520_));
  XNOR2_X1  g319(.A(G183gat), .B(G211gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n525_), .A2(KEYINPUT17), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n519_), .B(new_n526_), .ZN(new_n527_));
  NOR3_X1   g326(.A1(new_n518_), .A2(KEYINPUT17), .A3(new_n525_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n504_), .A2(new_n529_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n441_), .A2(new_n454_), .ZN(new_n531_));
  AND2_X1   g330(.A1(new_n513_), .A2(new_n516_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n472_), .A2(new_n517_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(G230gat), .ZN(new_n536_));
  INV_X1    g335(.A(G233gat), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n535_), .A2(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n538_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT12), .ZN(new_n541_));
  AND3_X1   g340(.A1(new_n472_), .A2(new_n517_), .A3(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n541_), .B1(new_n472_), .B2(new_n517_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n540_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G120gat), .B(G148gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT5), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G176gat), .B(G204gat), .ZN(new_n547_));
  XOR2_X1   g346(.A(new_n546_), .B(new_n547_), .Z(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n539_), .A2(new_n544_), .A3(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n549_), .B1(new_n539_), .B2(new_n544_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n553_), .A2(KEYINPUT13), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(KEYINPUT13), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT67), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(KEYINPUT67), .B1(new_n554_), .B2(new_n555_), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  AND2_X1   g359(.A1(new_n530_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(KEYINPUT79), .ZN(new_n562_));
  OR2_X1    g361(.A1(new_n561_), .A2(KEYINPUT79), .ZN(new_n563_));
  AND3_X1   g362(.A1(new_n417_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n332_), .A2(new_n333_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n564_), .A2(new_n377_), .A3(new_n566_), .ZN(new_n567_));
  OR2_X1    g366(.A1(new_n567_), .A2(KEYINPUT95), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(KEYINPUT95), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT38), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n529_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n560_), .A2(new_n416_), .A3(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(KEYINPUT96), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n498_), .B1(new_n481_), .B2(new_n499_), .ZN(new_n576_));
  AOI211_X1 g375(.A(KEYINPUT75), .B(new_n493_), .C1(new_n475_), .C2(new_n480_), .ZN(new_n577_));
  AOI21_X1  g376(.A(KEYINPUT73), .B1(new_n489_), .B2(new_n490_), .ZN(new_n578_));
  AND4_X1   g377(.A1(KEYINPUT73), .A2(new_n475_), .A3(new_n480_), .A4(new_n490_), .ZN(new_n579_));
  OAI22_X1  g378(.A1(new_n576_), .A2(new_n577_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT97), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n492_), .A2(new_n501_), .A3(KEYINPUT97), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT96), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n560_), .A2(new_n586_), .A3(new_n416_), .A4(new_n573_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n375_), .A2(new_n575_), .A3(new_n585_), .A4(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(G1gat), .B1(new_n588_), .B2(new_n565_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n568_), .A2(KEYINPUT38), .A3(new_n569_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n572_), .A2(new_n589_), .A3(new_n590_), .ZN(G1324gat));
  INV_X1    g390(.A(new_n370_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n564_), .A2(new_n378_), .A3(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(G8gat), .B1(new_n588_), .B2(new_n370_), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n594_), .A2(KEYINPUT39), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n594_), .A2(KEYINPUT39), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n593_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT40), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(G1325gat));
  OAI21_X1  g399(.A(G15gat), .B1(new_n588_), .B2(new_n356_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(KEYINPUT98), .B(KEYINPUT41), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n356_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n564_), .A2(new_n346_), .A3(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n601_), .A2(new_n602_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n603_), .A2(new_n605_), .A3(new_n606_), .ZN(G1326gat));
  NOR2_X1   g406(.A1(new_n254_), .A2(G22gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT101), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n564_), .A2(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(G22gat), .B1(new_n588_), .B2(new_n254_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(KEYINPUT100), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT100), .ZN(new_n613_));
  OAI211_X1 g412(.A(new_n613_), .B(G22gat), .C1(new_n588_), .C2(new_n254_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(KEYINPUT99), .B(KEYINPUT42), .ZN(new_n615_));
  AND3_X1   g414(.A1(new_n612_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n615_), .B1(new_n612_), .B2(new_n614_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n610_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT102), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  OAI211_X1 g419(.A(KEYINPUT102), .B(new_n610_), .C1(new_n616_), .C2(new_n617_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(G1327gat));
  NOR2_X1   g421(.A1(new_n585_), .A2(new_n573_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(new_n560_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n417_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(G29gat), .B1(new_n627_), .B2(new_n566_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT44), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n496_), .A2(new_n503_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT103), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n375_), .A2(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n630_), .A2(KEYINPUT43), .ZN(new_n633_));
  AOI22_X1  g432(.A1(new_n632_), .A2(KEYINPUT43), .B1(new_n375_), .B2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n560_), .A2(new_n416_), .A3(new_n529_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n629_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n635_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n375_), .A2(new_n633_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT43), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n640_), .B1(new_n375_), .B2(new_n631_), .ZN(new_n641_));
  OAI211_X1 g440(.A(KEYINPUT44), .B(new_n637_), .C1(new_n639_), .C2(new_n641_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n636_), .A2(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n565_), .A2(new_n385_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n628_), .B1(new_n643_), .B2(new_n644_), .ZN(G1328gat));
  NAND3_X1  g444(.A1(new_n636_), .A2(new_n592_), .A3(new_n642_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(G36gat), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n417_), .A2(new_n383_), .A3(new_n592_), .A4(new_n625_), .ZN(new_n648_));
  XOR2_X1   g447(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n649_));
  XNOR2_X1  g448(.A(new_n648_), .B(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n647_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT46), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n647_), .A2(KEYINPUT46), .A3(new_n650_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1329gat));
  NAND4_X1  g454(.A1(new_n636_), .A2(G43gat), .A3(new_n604_), .A4(new_n642_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n390_), .B1(new_n626_), .B2(new_n356_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g458(.A(G50gat), .B1(new_n627_), .B2(new_n372_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n254_), .A2(new_n388_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(new_n643_), .B2(new_n661_), .ZN(G1331gat));
  NOR2_X1   g461(.A1(new_n560_), .A2(new_n416_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n375_), .A2(new_n663_), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n664_), .A2(new_n530_), .ZN(new_n665_));
  INV_X1    g464(.A(G57gat), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n665_), .A2(new_n666_), .A3(new_n566_), .ZN(new_n667_));
  AND4_X1   g466(.A1(new_n375_), .A2(new_n573_), .A3(new_n585_), .A4(new_n663_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(G57gat), .B1(new_n669_), .B2(new_n565_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n667_), .A2(new_n670_), .ZN(G1332gat));
  INV_X1    g470(.A(G64gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n672_), .B1(new_n668_), .B2(new_n592_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT48), .Z(new_n674_));
  NAND3_X1  g473(.A1(new_n665_), .A2(new_n672_), .A3(new_n592_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(G1333gat));
  INV_X1    g475(.A(G71gat), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n677_), .B1(new_n668_), .B2(new_n604_), .ZN(new_n678_));
  XOR2_X1   g477(.A(new_n678_), .B(KEYINPUT49), .Z(new_n679_));
  NAND3_X1  g478(.A1(new_n665_), .A2(new_n677_), .A3(new_n604_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(G1334gat));
  AOI21_X1  g480(.A(new_n514_), .B1(new_n668_), .B2(new_n372_), .ZN(new_n682_));
  XOR2_X1   g481(.A(new_n682_), .B(KEYINPUT50), .Z(new_n683_));
  NAND3_X1  g482(.A1(new_n665_), .A2(new_n514_), .A3(new_n372_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(G1335gat));
  AND2_X1   g484(.A1(new_n664_), .A2(new_n623_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n686_), .A2(new_n419_), .A3(new_n566_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n632_), .A2(KEYINPUT43), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(new_n638_), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n560_), .A2(new_n416_), .A3(new_n573_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n691_), .A2(new_n566_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n687_), .B1(new_n692_), .B2(new_n419_), .ZN(G1336gat));
  AOI21_X1  g492(.A(G92gat), .B1(new_n686_), .B2(new_n592_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n370_), .A2(new_n420_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT105), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n694_), .B1(new_n691_), .B2(new_n696_), .ZN(G1337gat));
  AOI21_X1  g496(.A(new_n432_), .B1(new_n691_), .B2(new_n604_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n664_), .A2(new_n623_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n699_), .A2(new_n356_), .A3(new_n443_), .ZN(new_n700_));
  OR3_X1    g499(.A1(new_n698_), .A2(KEYINPUT51), .A3(new_n700_), .ZN(new_n701_));
  OAI21_X1  g500(.A(KEYINPUT51), .B1(new_n698_), .B2(new_n700_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(G1338gat));
  NAND3_X1  g502(.A1(new_n686_), .A2(new_n433_), .A3(new_n372_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n689_), .A2(new_n372_), .A3(new_n690_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT52), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n705_), .A2(new_n706_), .A3(G106gat), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n705_), .B2(G106gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n704_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(KEYINPUT106), .B(KEYINPUT53), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n709_), .A2(new_n711_), .ZN(new_n712_));
  OAI211_X1 g511(.A(new_n704_), .B(new_n710_), .C1(new_n707_), .C2(new_n708_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1339gat));
  INV_X1    g513(.A(KEYINPUT111), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT109), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT55), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n533_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n718_));
  AOI22_X1  g517(.A1(new_n544_), .A2(new_n717_), .B1(new_n718_), .B2(new_n538_), .ZN(new_n719_));
  OAI211_X1 g518(.A(new_n540_), .B(KEYINPUT55), .C1(new_n542_), .C2(new_n543_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n549_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n716_), .B1(new_n721_), .B2(KEYINPUT56), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n544_), .A2(new_n717_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n718_), .A2(new_n538_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n723_), .A2(new_n724_), .A3(new_n720_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n725_), .A2(KEYINPUT56), .A3(new_n548_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT108), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n548_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT56), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n728_), .A2(KEYINPUT109), .A3(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT108), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n725_), .A2(new_n731_), .A3(KEYINPUT56), .A4(new_n548_), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n722_), .A2(new_n727_), .A3(new_n730_), .A4(new_n732_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(KEYINPUT110), .A2(KEYINPUT58), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n411_), .B1(new_n396_), .B2(new_n406_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n406_), .B1(new_n398_), .B2(new_n395_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(new_n404_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n412_), .A2(new_n739_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n551_), .A2(new_n740_), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n733_), .A2(new_n735_), .A3(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n735_), .B1(new_n733_), .B2(new_n741_), .ZN(new_n743_));
  NOR3_X1   g542(.A1(new_n742_), .A2(new_n743_), .A3(new_n630_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT57), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n553_), .A2(new_n740_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n728_), .A2(new_n729_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(new_n726_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n415_), .A2(new_n551_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n746_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n745_), .B1(new_n584_), .B2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n726_), .ZN(new_n752_));
  AOI21_X1  g551(.A(KEYINPUT56), .B1(new_n725_), .B2(new_n548_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n749_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n746_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n756_), .A2(KEYINPUT57), .A3(new_n582_), .A4(new_n583_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n751_), .A2(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n715_), .B1(new_n744_), .B2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n733_), .A2(new_n741_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(new_n734_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n733_), .A2(new_n735_), .A3(new_n741_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n761_), .A2(new_n504_), .A3(new_n762_), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n763_), .A2(KEYINPUT111), .A3(new_n751_), .A4(new_n757_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n759_), .A2(new_n529_), .A3(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT107), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n766_), .B1(new_n573_), .B2(new_n415_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n529_), .A2(KEYINPUT107), .A3(new_n416_), .ZN(new_n768_));
  NOR3_X1   g567(.A1(new_n767_), .A2(new_n556_), .A3(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(new_n630_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT54), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT54), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n769_), .A2(new_n772_), .A3(new_n630_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n765_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT112), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n765_), .A2(KEYINPUT112), .A3(new_n774_), .ZN(new_n778_));
  AND3_X1   g577(.A1(new_n373_), .A2(new_n566_), .A3(new_n604_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n777_), .A2(new_n778_), .A3(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT113), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n780_), .B(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(new_n416_), .ZN(new_n783_));
  INV_X1    g582(.A(G113gat), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n780_), .A2(KEYINPUT59), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n529_), .B1(new_n744_), .B2(new_n758_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n774_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT59), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n787_), .A2(new_n788_), .A3(new_n779_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n785_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n416_), .A2(G113gat), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n792_), .B(KEYINPUT114), .ZN(new_n793_));
  AOI22_X1  g592(.A1(new_n783_), .A2(new_n784_), .B1(new_n791_), .B2(new_n793_), .ZN(G1340gat));
  INV_X1    g593(.A(new_n560_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n785_), .A2(new_n795_), .A3(new_n789_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT116), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n785_), .A2(KEYINPUT116), .A3(new_n795_), .A4(new_n789_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n798_), .A2(G120gat), .A3(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT60), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT115), .B1(new_n801_), .B2(G120gat), .ZN(new_n802_));
  AOI21_X1  g601(.A(G120gat), .B1(new_n795_), .B2(new_n801_), .ZN(new_n803_));
  MUX2_X1   g602(.A(new_n802_), .B(KEYINPUT115), .S(new_n803_), .Z(new_n804_));
  NAND2_X1  g603(.A1(new_n782_), .A2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n800_), .A2(new_n805_), .ZN(G1341gat));
  INV_X1    g605(.A(G127gat), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n782_), .A2(new_n807_), .A3(new_n573_), .ZN(new_n808_));
  OAI21_X1  g607(.A(G127gat), .B1(new_n790_), .B2(new_n529_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(G1342gat));
  INV_X1    g609(.A(G134gat), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n782_), .A2(new_n811_), .A3(new_n584_), .ZN(new_n812_));
  OAI21_X1  g611(.A(G134gat), .B1(new_n790_), .B2(new_n630_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(G1343gat));
  AND3_X1   g613(.A1(new_n765_), .A2(KEYINPUT112), .A3(new_n774_), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT112), .B1(new_n765_), .B2(new_n774_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n254_), .A2(new_n604_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n817_), .A2(new_n566_), .A3(new_n370_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n818_), .B(KEYINPUT117), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  NOR3_X1   g619(.A1(new_n815_), .A2(new_n816_), .A3(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n416_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n822_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n795_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n824_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g624(.A(KEYINPUT61), .B(G155gat), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n815_), .A2(new_n816_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT118), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n828_), .A2(new_n829_), .A3(new_n573_), .A4(new_n819_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n777_), .A2(new_n573_), .A3(new_n778_), .A4(new_n819_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(KEYINPUT118), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT119), .ZN(new_n833_));
  AND3_X1   g632(.A1(new_n830_), .A2(new_n832_), .A3(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n833_), .B1(new_n830_), .B2(new_n832_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n827_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n829_), .B1(new_n821_), .B2(new_n573_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n831_), .A2(KEYINPUT118), .ZN(new_n838_));
  OAI21_X1  g637(.A(KEYINPUT119), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n830_), .A2(new_n832_), .A3(new_n833_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n839_), .A2(new_n826_), .A3(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n836_), .A2(new_n841_), .ZN(G1346gat));
  NAND4_X1  g641(.A1(new_n777_), .A2(new_n584_), .A3(new_n778_), .A4(new_n819_), .ZN(new_n843_));
  INV_X1    g642(.A(G162gat), .ZN(new_n844_));
  AND3_X1   g643(.A1(new_n843_), .A2(KEYINPUT120), .A3(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(KEYINPUT120), .B1(new_n843_), .B2(new_n844_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n821_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n631_), .A2(G162gat), .ZN(new_n848_));
  OAI22_X1  g647(.A1(new_n845_), .A2(new_n846_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(KEYINPUT121), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT121), .ZN(new_n851_));
  OAI221_X1 g650(.A(new_n851_), .B1(new_n847_), .B2(new_n848_), .C1(new_n845_), .C2(new_n846_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n852_), .ZN(G1347gat));
  NAND2_X1  g652(.A1(new_n592_), .A2(new_n369_), .ZN(new_n854_));
  XOR2_X1   g653(.A(new_n854_), .B(KEYINPUT122), .Z(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n254_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n787_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n416_), .ZN(new_n859_));
  AOI21_X1  g658(.A(KEYINPUT123), .B1(new_n859_), .B2(G169gat), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT62), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n859_), .A2(KEYINPUT123), .A3(G169gat), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n860_), .A2(new_n861_), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n864_), .B(new_n865_), .C1(new_n283_), .C2(new_n859_), .ZN(G1348gat));
  AOI21_X1  g665(.A(new_n303_), .B1(new_n858_), .B2(new_n795_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n777_), .A2(new_n778_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n868_), .A2(new_n372_), .ZN(new_n869_));
  AND3_X1   g668(.A1(new_n855_), .A2(G176gat), .A3(new_n795_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n867_), .B1(new_n869_), .B2(new_n870_), .ZN(G1349gat));
  INV_X1    g670(.A(new_n858_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n872_), .A2(new_n293_), .A3(new_n529_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n869_), .A2(new_n573_), .A3(new_n855_), .ZN(new_n874_));
  INV_X1    g673(.A(G183gat), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n873_), .B1(new_n874_), .B2(new_n875_), .ZN(G1350gat));
  OAI21_X1  g675(.A(G190gat), .B1(new_n872_), .B2(new_n630_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n858_), .A2(new_n294_), .A3(new_n584_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(G1351gat));
  NAND3_X1  g678(.A1(new_n817_), .A2(new_n592_), .A3(new_n565_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n777_), .A2(new_n416_), .A3(new_n778_), .A4(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT124), .ZN(new_n883_));
  OR3_X1    g682(.A1(new_n882_), .A2(new_n883_), .A3(KEYINPUT125), .ZN(new_n884_));
  OAI21_X1  g683(.A(KEYINPUT125), .B1(new_n882_), .B2(new_n883_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n882_), .A2(new_n883_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(G197gat), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n888_), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n884_), .A2(G197gat), .A3(new_n885_), .A4(new_n887_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(G1352gat));
  NOR2_X1   g690(.A1(new_n868_), .A2(new_n880_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n795_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g693(.A(KEYINPUT126), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n529_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n892_), .A2(new_n895_), .A3(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n895_), .B1(new_n892_), .B2(new_n896_), .ZN(new_n899_));
  OAI22_X1  g698(.A1(new_n898_), .A2(new_n899_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n900_));
  INV_X1    g699(.A(new_n899_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n901_), .A2(new_n902_), .A3(new_n897_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n900_), .A2(new_n903_), .ZN(G1354gat));
  NOR4_X1   g703(.A1(new_n868_), .A2(G218gat), .A3(new_n585_), .A4(new_n880_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(G218gat), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n868_), .A2(new_n630_), .A3(new_n880_), .ZN(new_n908_));
  OAI211_X1 g707(.A(new_n906_), .B(KEYINPUT127), .C1(new_n907_), .C2(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT127), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n908_), .A2(new_n907_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n911_), .B2(new_n905_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n909_), .A2(new_n912_), .ZN(G1355gat));
endmodule


