//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 0 1 1 1 1 1 1 0 0 0 0 0 0 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 0 0 1 1 1 0 1 0 1 1 1 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n638_, new_n639_, new_n640_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n699_, new_n700_, new_n701_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n828_, new_n829_, new_n831_, new_n832_,
    new_n833_, new_n835_, new_n836_, new_n837_, new_n839_, new_n840_,
    new_n842_, new_n843_, new_n844_, new_n846_, new_n847_, new_n848_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n871_, new_n872_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n889_, new_n890_;
  INV_X1    g000(.A(KEYINPUT97), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT27), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G226gat), .A2(G233gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT19), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT84), .B(G204gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(G197gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT21), .ZN(new_n208_));
  INV_X1    g007(.A(G204gat), .ZN(new_n209_));
  OAI211_X1 g008(.A(new_n207_), .B(new_n208_), .C1(G197gat), .C2(new_n209_), .ZN(new_n210_));
  XOR2_X1   g009(.A(G211gat), .B(G218gat), .Z(new_n211_));
  INV_X1    g010(.A(G197gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n206_), .A2(new_n212_), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n208_), .B1(G197gat), .B2(G204gat), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n211_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n210_), .A2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT85), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n207_), .B1(G197gat), .B2(new_n209_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(KEYINPUT21), .A3(new_n211_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(G183gat), .ZN(new_n221_));
  INV_X1    g020(.A(G190gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT23), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NOR3_X1   g023(.A1(new_n221_), .A2(new_n222_), .A3(KEYINPUT23), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n224_), .B1(new_n226_), .B2(KEYINPUT79), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n227_), .B1(KEYINPUT79), .B2(new_n226_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n221_), .A2(new_n222_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(KEYINPUT22), .B(G169gat), .ZN(new_n231_));
  INV_X1    g030(.A(G176gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G169gat), .A2(G176gat), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n230_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(G169gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(new_n232_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n237_), .A2(KEYINPUT24), .ZN(new_n238_));
  AND3_X1   g037(.A1(new_n237_), .A2(KEYINPUT24), .A3(new_n234_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(KEYINPUT25), .B(G183gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT26), .B(G190gat), .ZN(new_n241_));
  AOI211_X1 g040(.A(new_n238_), .B(new_n239_), .C1(new_n240_), .C2(new_n241_), .ZN(new_n242_));
  OR2_X1    g041(.A1(new_n223_), .A2(KEYINPUT78), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n223_), .A2(KEYINPUT78), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n243_), .A2(new_n226_), .A3(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n242_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n235_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n220_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n245_), .A2(new_n229_), .ZN(new_n249_));
  XOR2_X1   g048(.A(new_n234_), .B(KEYINPUT88), .Z(new_n250_));
  NAND3_X1  g049(.A1(new_n249_), .A2(new_n233_), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n242_), .A2(new_n228_), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n217_), .A2(new_n219_), .A3(new_n251_), .A4(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n248_), .A2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(KEYINPUT94), .B(KEYINPUT20), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n205_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n251_), .A2(new_n252_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n220_), .A2(new_n257_), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n258_), .B(KEYINPUT20), .C1(new_n247_), .C2(new_n220_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n256_), .B1(new_n205_), .B2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G8gat), .B(G36gat), .ZN(new_n261_));
  INV_X1    g060(.A(G92gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n261_), .B(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT18), .B(G64gat), .ZN(new_n264_));
  XOR2_X1   g063(.A(new_n263_), .B(new_n264_), .Z(new_n265_));
  AOI21_X1  g064(.A(new_n203_), .B1(new_n260_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT20), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n205_), .A2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n248_), .A2(new_n253_), .A3(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT89), .ZN(new_n270_));
  OR2_X1    g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n265_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n259_), .A2(new_n205_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n269_), .A2(new_n270_), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n271_), .A2(new_n272_), .A3(new_n273_), .A4(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n266_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT95), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n266_), .A2(KEYINPUT95), .A3(new_n275_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n271_), .A2(new_n274_), .A3(new_n273_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(new_n265_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(new_n275_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT96), .B(KEYINPUT27), .ZN(new_n283_));
  AOI22_X1  g082(.A1(new_n278_), .A2(new_n279_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(G78gat), .B(G106gat), .Z(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(G50gat), .ZN(new_n287_));
  NOR2_X1   g086(.A1(G155gat), .A2(G162gat), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT83), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G155gat), .A2(G162gat), .ZN(new_n291_));
  NOR2_X1   g090(.A1(G141gat), .A2(G148gat), .ZN(new_n292_));
  XOR2_X1   g091(.A(new_n292_), .B(KEYINPUT3), .Z(new_n293_));
  NAND2_X1  g092(.A1(G141gat), .A2(G148gat), .ZN(new_n294_));
  XOR2_X1   g093(.A(new_n294_), .B(KEYINPUT2), .Z(new_n295_));
  OAI211_X1 g094(.A(new_n290_), .B(new_n291_), .C1(new_n293_), .C2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT1), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n291_), .B(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n290_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n292_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n299_), .A2(new_n300_), .A3(new_n294_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n296_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT28), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT29), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n303_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(G22gat), .ZN(new_n307_));
  OAI21_X1  g106(.A(KEYINPUT28), .B1(new_n302_), .B2(KEYINPUT29), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n306_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n307_), .B1(new_n306_), .B2(new_n308_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n287_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NOR3_X1   g112(.A1(new_n310_), .A2(new_n287_), .A3(new_n311_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n286_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n314_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n286_), .A2(KEYINPUT87), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n316_), .A2(new_n317_), .A3(new_n312_), .ZN(new_n318_));
  AND2_X1   g117(.A1(G228gat), .A2(G233gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(KEYINPUT86), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n220_), .B1(new_n305_), .B2(new_n303_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n319_), .A2(KEYINPUT86), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n320_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n321_), .A2(KEYINPUT86), .A3(new_n319_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n315_), .A2(new_n318_), .A3(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n326_), .B1(new_n315_), .B2(new_n318_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G127gat), .B(G134gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(G120gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT82), .B(G113gat), .ZN(new_n332_));
  OR2_X1    g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n332_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(new_n302_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n333_), .A2(new_n334_), .A3(new_n301_), .A4(new_n296_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G225gat), .A2(G233gat), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n336_), .A2(KEYINPUT4), .A3(new_n337_), .ZN(new_n342_));
  OR2_X1    g141(.A1(new_n342_), .A2(KEYINPUT90), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n342_), .B(KEYINPUT90), .C1(KEYINPUT4), .C2(new_n336_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n341_), .B1(new_n345_), .B2(new_n340_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G1gat), .B(G29gat), .ZN(new_n347_));
  INV_X1    g146(.A(G85gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT0), .B(G57gat), .ZN(new_n350_));
  XOR2_X1   g149(.A(new_n349_), .B(new_n350_), .Z(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n346_), .A2(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n339_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n351_), .B1(new_n354_), .B2(new_n341_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n353_), .A2(new_n355_), .ZN(new_n356_));
  NOR3_X1   g155(.A1(new_n328_), .A2(new_n329_), .A3(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT93), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n272_), .A2(KEYINPUT32), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n358_), .B1(new_n280_), .B2(new_n360_), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n273_), .A2(new_n274_), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n362_), .A2(KEYINPUT93), .A3(new_n271_), .A4(new_n359_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n260_), .A2(new_n360_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n361_), .A2(new_n363_), .A3(new_n356_), .A4(new_n364_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(KEYINPUT91), .A2(KEYINPUT33), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n353_), .A2(new_n366_), .ZN(new_n367_));
  OAI211_X1 g166(.A(new_n346_), .B(new_n352_), .C1(KEYINPUT91), .C2(KEYINPUT33), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n340_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n351_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n370_));
  OR3_X1    g169(.A1(new_n369_), .A2(KEYINPUT92), .A3(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(KEYINPUT92), .B1(new_n369_), .B2(new_n370_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n367_), .A2(new_n368_), .A3(new_n371_), .A4(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n365_), .B1(new_n373_), .B2(new_n282_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n328_), .A2(new_n329_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  AOI22_X1  g175(.A1(new_n284_), .A2(new_n357_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n377_));
  XOR2_X1   g176(.A(KEYINPUT80), .B(KEYINPUT30), .Z(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT31), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n247_), .B(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(G43gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G71gat), .B(G99gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n335_), .B(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G227gat), .A2(G233gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(KEYINPUT81), .ZN(new_n386_));
  INV_X1    g185(.A(G15gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n386_), .B(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n384_), .B(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  OR2_X1    g189(.A1(new_n382_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n382_), .A2(new_n390_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n202_), .B1(new_n377_), .B2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n374_), .A2(new_n376_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n278_), .A2(new_n279_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n282_), .A2(new_n283_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n396_), .A2(new_n397_), .A3(new_n357_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n395_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n393_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n399_), .A2(KEYINPUT97), .A3(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n356_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n284_), .A2(new_n393_), .A3(new_n376_), .A4(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n394_), .A2(new_n401_), .A3(new_n403_), .ZN(new_n404_));
  AND3_X1   g203(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n405_));
  AOI21_X1  g204(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n406_));
  NOR3_X1   g205(.A1(new_n405_), .A2(new_n406_), .A3(KEYINPUT64), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT64), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G99gat), .A2(G106gat), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT6), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n408_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n407_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n348_), .A2(new_n262_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G85gat), .A2(G92gat), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n415_), .A2(KEYINPUT9), .A3(new_n416_), .ZN(new_n417_));
  OR2_X1    g216(.A1(new_n416_), .A2(KEYINPUT9), .ZN(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT10), .B(G99gat), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n417_), .B(new_n418_), .C1(G106gat), .C2(new_n419_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n414_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n411_), .A2(new_n412_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT7), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n423_), .B(KEYINPUT65), .C1(G99gat), .C2(G106gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(KEYINPUT65), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT65), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT7), .ZN(new_n427_));
  NOR2_X1   g226(.A1(G99gat), .A2(G106gat), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n425_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n422_), .B1(new_n424_), .B2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n415_), .A2(new_n416_), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT8), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(G99gat), .ZN(new_n433_));
  INV_X1    g232(.A(G106gat), .ZN(new_n434_));
  OAI211_X1 g233(.A(new_n433_), .B(new_n434_), .C1(new_n426_), .C2(KEYINPUT7), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n423_), .A2(KEYINPUT65), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n424_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n437_), .B1(new_n407_), .B2(new_n413_), .ZN(new_n438_));
  AND2_X1   g237(.A1(new_n415_), .A2(new_n416_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT8), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n438_), .A2(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n421_), .B1(new_n432_), .B2(new_n443_), .ZN(new_n444_));
  AND2_X1   g243(.A1(G57gat), .A2(G64gat), .ZN(new_n445_));
  NOR2_X1   g244(.A1(G57gat), .A2(G64gat), .ZN(new_n446_));
  OAI21_X1  g245(.A(KEYINPUT11), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(G57gat), .ZN(new_n448_));
  INV_X1    g247(.A(G64gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT11), .ZN(new_n451_));
  NAND2_X1  g250(.A1(G57gat), .A2(G64gat), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n450_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(G78gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(G71gat), .ZN(new_n455_));
  INV_X1    g254(.A(G71gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(G78gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n447_), .A2(new_n453_), .A3(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n450_), .A2(new_n452_), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n460_), .A2(KEYINPUT11), .A3(new_n455_), .A4(new_n457_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n459_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT66), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n459_), .A2(new_n461_), .A3(KEYINPUT66), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n464_), .A2(KEYINPUT12), .A3(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(KEYINPUT67), .B1(new_n444_), .B2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n465_), .A2(KEYINPUT12), .ZN(new_n468_));
  AOI21_X1  g267(.A(KEYINPUT66), .B1(new_n459_), .B2(new_n461_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  OR2_X1    g269(.A1(new_n419_), .A2(G106gat), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT64), .B1(new_n405_), .B2(new_n406_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n411_), .A2(new_n408_), .A3(new_n412_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n471_), .A2(new_n474_), .A3(new_n418_), .A4(new_n417_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n405_), .A2(new_n406_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n437_), .A2(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n440_), .B1(new_n477_), .B2(new_n439_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n441_), .B1(new_n474_), .B2(new_n437_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n475_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT67), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n470_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n467_), .A2(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n431_), .B1(new_n437_), .B2(new_n476_), .ZN(new_n484_));
  AOI22_X1  g283(.A1(new_n472_), .A2(new_n473_), .B1(new_n429_), .B2(new_n424_), .ZN(new_n485_));
  OAI22_X1  g284(.A1(new_n484_), .A2(new_n440_), .B1(new_n485_), .B2(new_n441_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n486_), .A2(new_n475_), .A3(new_n462_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT12), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n480_), .A2(new_n461_), .A3(new_n459_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G230gat), .A2(G233gat), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n483_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n489_), .A2(new_n487_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n493_), .A2(G230gat), .A3(G233gat), .ZN(new_n494_));
  AND2_X1   g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G120gat), .B(G148gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(G204gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(KEYINPUT5), .B(G176gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n495_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  XOR2_X1   g300(.A(new_n499_), .B(KEYINPUT68), .Z(new_n502_));
  NOR2_X1   g301(.A1(new_n495_), .A2(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n501_), .A2(new_n503_), .ZN(new_n504_));
  XOR2_X1   g303(.A(KEYINPUT69), .B(KEYINPUT13), .Z(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n500_), .B1(new_n495_), .B2(new_n502_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT69), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n507_), .B1(new_n508_), .B2(KEYINPUT13), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n506_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G1gat), .B(G8gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT75), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G15gat), .B(G22gat), .ZN(new_n514_));
  INV_X1    g313(.A(G1gat), .ZN(new_n515_));
  INV_X1    g314(.A(G8gat), .ZN(new_n516_));
  OAI21_X1  g315(.A(KEYINPUT14), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n514_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n513_), .B(new_n518_), .ZN(new_n519_));
  XOR2_X1   g318(.A(G43gat), .B(G50gat), .Z(new_n520_));
  XNOR2_X1  g319(.A(G29gat), .B(G36gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT15), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G43gat), .B(G50gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n521_), .B(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT15), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n524_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n519_), .A2(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n529_), .B1(new_n522_), .B2(new_n519_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(KEYINPUT76), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G229gat), .A2(G233gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT77), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT76), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n529_), .A2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n531_), .A2(new_n534_), .A3(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n519_), .B(new_n522_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n538_), .A2(G229gat), .A3(G233gat), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n537_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G113gat), .B(G141gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G169gat), .B(G197gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n540_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n543_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n537_), .A2(new_n539_), .A3(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n511_), .A2(new_n548_), .ZN(new_n549_));
  AND2_X1   g348(.A1(new_n404_), .A2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n519_), .B(new_n462_), .ZN(new_n551_));
  AND2_X1   g350(.A1(G231gat), .A2(G233gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(G127gat), .B(G155gat), .Z(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(G211gat), .ZN(new_n556_));
  XOR2_X1   g355(.A(KEYINPUT16), .B(G183gat), .Z(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n558_), .A2(new_n463_), .A3(KEYINPUT17), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n559_), .B1(KEYINPUT17), .B2(new_n558_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n554_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n553_), .A2(new_n559_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G232gat), .A2(G233gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT34), .ZN(new_n566_));
  XOR2_X1   g365(.A(KEYINPUT70), .B(KEYINPUT35), .Z(new_n567_));
  NOR2_X1   g366(.A1(new_n480_), .A2(new_n522_), .ZN(new_n568_));
  AOI22_X1  g367(.A1(new_n475_), .A2(new_n486_), .B1(new_n524_), .B2(new_n527_), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n566_), .B(new_n567_), .C1(new_n568_), .C2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n444_), .A2(new_n526_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n480_), .A2(new_n528_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n566_), .A2(new_n567_), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n566_), .A2(new_n567_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n571_), .A2(new_n572_), .A3(new_n573_), .A4(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n570_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT73), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n570_), .A2(KEYINPUT73), .A3(new_n575_), .ZN(new_n579_));
  XOR2_X1   g378(.A(G190gat), .B(G218gat), .Z(new_n580_));
  XNOR2_X1  g379(.A(G134gat), .B(G162gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n582_), .B(KEYINPUT36), .Z(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n578_), .A2(new_n579_), .A3(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT37), .ZN(new_n586_));
  XOR2_X1   g385(.A(KEYINPUT71), .B(KEYINPUT36), .Z(new_n587_));
  NAND2_X1  g386(.A1(new_n582_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  AND3_X1   g388(.A1(new_n570_), .A2(new_n575_), .A3(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n585_), .A2(new_n586_), .A3(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n583_), .B1(new_n570_), .B2(new_n575_), .ZN(new_n593_));
  OAI21_X1  g392(.A(KEYINPUT37), .B1(new_n590_), .B2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT72), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  OAI211_X1 g395(.A(KEYINPUT72), .B(KEYINPUT37), .C1(new_n590_), .C2(new_n593_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n592_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(KEYINPUT74), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT74), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n592_), .A2(new_n596_), .A3(new_n600_), .A4(new_n597_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n564_), .B1(new_n599_), .B2(new_n601_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n550_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n603_), .A2(new_n515_), .A3(new_n356_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT38), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT98), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n604_), .A2(new_n605_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT99), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n585_), .A2(new_n591_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n564_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n550_), .A2(new_n611_), .ZN(new_n612_));
  OAI21_X1  g411(.A(G1gat), .B1(new_n612_), .B2(new_n402_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n607_), .A2(new_n609_), .A3(new_n613_), .ZN(G1324gat));
  AND2_X1   g413(.A1(new_n550_), .A2(new_n611_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n284_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT100), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT39), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n617_), .A2(new_n618_), .A3(new_n619_), .A4(G8gat), .ZN(new_n620_));
  OAI211_X1 g419(.A(new_n619_), .B(G8gat), .C1(new_n612_), .C2(new_n284_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(KEYINPUT100), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n516_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n623_));
  OAI211_X1 g422(.A(new_n620_), .B(new_n622_), .C1(new_n619_), .C2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n603_), .A2(new_n516_), .A3(new_n616_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT102), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n626_), .A2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n624_), .A2(new_n625_), .A3(new_n628_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(G1325gat));
  OAI21_X1  g431(.A(G15gat), .B1(new_n612_), .B2(new_n400_), .ZN(new_n633_));
  OR2_X1    g432(.A1(new_n633_), .A2(KEYINPUT41), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(KEYINPUT41), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n603_), .A2(new_n387_), .A3(new_n393_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n634_), .A2(new_n635_), .A3(new_n636_), .ZN(G1326gat));
  OAI21_X1  g436(.A(G22gat), .B1(new_n612_), .B2(new_n376_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT42), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n603_), .A2(new_n307_), .A3(new_n375_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(G1327gat));
  NOR3_X1   g440(.A1(new_n511_), .A2(new_n548_), .A3(new_n563_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT43), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n599_), .A2(new_n601_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  AND3_X1   g444(.A1(new_n404_), .A2(new_n643_), .A3(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n643_), .B1(new_n404_), .B2(new_n645_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n642_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT44), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  OAI211_X1 g449(.A(KEYINPUT44), .B(new_n642_), .C1(new_n646_), .C2(new_n647_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n650_), .A2(new_n356_), .A3(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(G29gat), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n564_), .A2(new_n610_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n550_), .A2(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n402_), .A2(G29gat), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n656_), .B(KEYINPUT103), .Z(new_n657_));
  OAI21_X1  g456(.A(new_n653_), .B1(new_n655_), .B2(new_n657_), .ZN(G1328gat));
  NAND2_X1  g457(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n659_));
  NOR2_X1   g458(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT105), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n650_), .A2(new_n616_), .A3(new_n651_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n662_), .A2(G36gat), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n284_), .A2(G36gat), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n550_), .A2(new_n654_), .A3(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT45), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n665_), .B(new_n666_), .ZN(new_n667_));
  OAI211_X1 g466(.A(new_n659_), .B(new_n661_), .C1(new_n663_), .C2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n661_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n667_), .B1(new_n662_), .B2(G36gat), .ZN(new_n670_));
  INV_X1    g469(.A(new_n659_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n669_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n668_), .A2(new_n672_), .ZN(G1329gat));
  NAND4_X1  g472(.A1(new_n650_), .A2(G43gat), .A3(new_n393_), .A4(new_n651_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n381_), .B1(new_n655_), .B2(new_n400_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  XOR2_X1   g475(.A(KEYINPUT106), .B(KEYINPUT47), .Z(new_n677_));
  XNOR2_X1  g476(.A(new_n676_), .B(new_n677_), .ZN(G1330gat));
  NAND3_X1  g477(.A1(new_n650_), .A2(new_n375_), .A3(new_n651_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT107), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n287_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n681_), .B1(new_n680_), .B2(new_n679_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n375_), .A2(new_n287_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n682_), .B1(new_n655_), .B2(new_n683_), .ZN(G1331gat));
  AND3_X1   g483(.A1(new_n404_), .A2(new_n548_), .A3(new_n511_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n685_), .A2(new_n602_), .ZN(new_n686_));
  AOI21_X1  g485(.A(G57gat), .B1(new_n686_), .B2(new_n356_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n685_), .A2(new_n611_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n402_), .A2(new_n448_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n687_), .B1(new_n688_), .B2(new_n689_), .ZN(G1332gat));
  AOI21_X1  g489(.A(new_n449_), .B1(new_n688_), .B2(new_n616_), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT48), .Z(new_n692_));
  NAND3_X1  g491(.A1(new_n686_), .A2(new_n449_), .A3(new_n616_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1333gat));
  AOI21_X1  g493(.A(new_n456_), .B1(new_n688_), .B2(new_n393_), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT49), .Z(new_n696_));
  NAND3_X1  g495(.A1(new_n686_), .A2(new_n456_), .A3(new_n393_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(G1334gat));
  AOI21_X1  g497(.A(new_n454_), .B1(new_n688_), .B2(new_n375_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT50), .Z(new_n700_));
  NAND3_X1  g499(.A1(new_n686_), .A2(new_n454_), .A3(new_n375_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(G1335gat));
  NAND2_X1  g501(.A1(new_n685_), .A2(new_n654_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(G85gat), .B1(new_n704_), .B2(new_n356_), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n646_), .A2(new_n647_), .ZN(new_n706_));
  NOR3_X1   g505(.A1(new_n510_), .A2(new_n547_), .A3(new_n563_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n402_), .A2(new_n348_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n705_), .B1(new_n708_), .B2(new_n709_), .ZN(G1336gat));
  NAND2_X1  g509(.A1(new_n616_), .A2(G92gat), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT108), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n708_), .A2(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n262_), .B1(new_n703_), .B2(new_n284_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT109), .ZN(G1337gat));
  AOI21_X1  g515(.A(new_n433_), .B1(new_n708_), .B2(new_n393_), .ZN(new_n717_));
  NOR3_X1   g516(.A1(new_n703_), .A2(new_n419_), .A3(new_n400_), .ZN(new_n718_));
  OR3_X1    g517(.A1(new_n717_), .A2(KEYINPUT51), .A3(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(KEYINPUT51), .B1(new_n717_), .B2(new_n718_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(G1338gat));
  NAND3_X1  g520(.A1(new_n704_), .A2(new_n434_), .A3(new_n375_), .ZN(new_n722_));
  OAI211_X1 g521(.A(new_n375_), .B(new_n707_), .C1(new_n646_), .C2(new_n647_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(G106gat), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT110), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n724_), .A2(new_n725_), .A3(KEYINPUT52), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT52), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n723_), .A2(new_n727_), .A3(G106gat), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n725_), .B1(new_n724_), .B2(KEYINPUT52), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n722_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(KEYINPUT53), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT53), .ZN(new_n733_));
  OAI211_X1 g532(.A(new_n733_), .B(new_n722_), .C1(new_n729_), .C2(new_n730_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(G1339gat));
  NOR4_X1   g534(.A1(new_n616_), .A2(new_n400_), .A3(new_n375_), .A4(new_n402_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n491_), .B1(new_n483_), .B2(new_n490_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT55), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n492_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n483_), .A2(new_n490_), .A3(KEYINPUT55), .A4(new_n491_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n502_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT56), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n742_), .A2(KEYINPUT56), .A3(new_n743_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n531_), .A2(new_n533_), .A3(new_n536_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n545_), .B1(new_n538_), .B2(new_n534_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n546_), .A2(new_n751_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n501_), .A2(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(KEYINPUT58), .B1(new_n748_), .B2(new_n753_), .ZN(new_n754_));
  OAI21_X1  g553(.A(KEYINPUT112), .B1(new_n754_), .B2(new_n644_), .ZN(new_n755_));
  AOI21_X1  g554(.A(KEYINPUT56), .B1(new_n742_), .B2(new_n743_), .ZN(new_n756_));
  AOI211_X1 g555(.A(new_n745_), .B(new_n502_), .C1(new_n740_), .C2(new_n741_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n753_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT58), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT112), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n760_), .A2(new_n761_), .A3(new_n599_), .A4(new_n601_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n748_), .A2(KEYINPUT58), .A3(new_n753_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n755_), .A2(new_n762_), .A3(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT57), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n504_), .A2(new_n752_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n548_), .A2(new_n501_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n748_), .B2(new_n768_), .ZN(new_n769_));
  OAI211_X1 g568(.A(KEYINPUT111), .B(new_n766_), .C1(new_n769_), .C2(new_n610_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT111), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n547_), .B(new_n500_), .C1(new_n756_), .C2(new_n757_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n507_), .A2(new_n546_), .A3(new_n751_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n610_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n771_), .B1(new_n774_), .B2(KEYINPUT57), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(KEYINPUT57), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n770_), .A2(new_n775_), .A3(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n564_), .B1(new_n765_), .B2(new_n777_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n511_), .A2(new_n547_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT54), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n779_), .A2(new_n780_), .A3(new_n602_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n780_), .B1(new_n779_), .B2(new_n602_), .ZN(new_n782_));
  OR2_X1    g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n737_), .B1(new_n778_), .B2(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(G113gat), .B1(new_n784_), .B2(new_n547_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n781_), .A2(new_n782_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n766_), .B1(new_n769_), .B2(new_n610_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n764_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT114), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n764_), .A2(KEYINPUT114), .A3(new_n787_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n790_), .A2(new_n776_), .A3(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n786_), .B1(new_n792_), .B2(new_n564_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT59), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n736_), .A2(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(KEYINPUT115), .B1(new_n793_), .B2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n791_), .A2(new_n776_), .ZN(new_n797_));
  AOI21_X1  g596(.A(KEYINPUT114), .B1(new_n764_), .B2(new_n787_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n564_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n783_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT115), .ZN(new_n801_));
  INV_X1    g600(.A(new_n795_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n800_), .A2(new_n801_), .A3(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(KEYINPUT113), .B1(new_n784_), .B2(new_n794_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT113), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n764_), .A2(new_n775_), .A3(new_n770_), .A4(new_n776_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n786_), .B1(new_n806_), .B2(new_n564_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n805_), .B(KEYINPUT59), .C1(new_n807_), .C2(new_n737_), .ZN(new_n808_));
  AOI22_X1  g607(.A1(new_n796_), .A2(new_n803_), .B1(new_n804_), .B2(new_n808_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n548_), .A2(KEYINPUT116), .ZN(new_n810_));
  MUX2_X1   g609(.A(KEYINPUT116), .B(new_n810_), .S(G113gat), .Z(new_n811_));
  AOI21_X1  g610(.A(new_n785_), .B1(new_n809_), .B2(new_n811_), .ZN(G1340gat));
  INV_X1    g611(.A(G120gat), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n813_), .B1(new_n510_), .B2(KEYINPUT60), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n784_), .B(new_n814_), .C1(KEYINPUT60), .C2(new_n813_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n804_), .A2(new_n808_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n801_), .B1(new_n800_), .B2(new_n802_), .ZN(new_n817_));
  AOI211_X1 g616(.A(KEYINPUT115), .B(new_n795_), .C1(new_n799_), .C2(new_n783_), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n511_), .B(new_n816_), .C1(new_n817_), .C2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT117), .ZN(new_n820_));
  OAI21_X1  g619(.A(G120gat), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(KEYINPUT117), .B1(new_n809_), .B2(new_n511_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n815_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT118), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT118), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n825_), .B(new_n815_), .C1(new_n821_), .C2(new_n822_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n826_), .ZN(G1341gat));
  AOI21_X1  g626(.A(G127gat), .B1(new_n784_), .B2(new_n563_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n563_), .A2(G127gat), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n828_), .B1(new_n809_), .B2(new_n829_), .ZN(G1342gat));
  AOI21_X1  g629(.A(G134gat), .B1(new_n784_), .B2(new_n610_), .ZN(new_n831_));
  XNOR2_X1  g630(.A(new_n831_), .B(KEYINPUT119), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n645_), .A2(G134gat), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n832_), .B1(new_n809_), .B2(new_n833_), .ZN(G1343gat));
  NOR3_X1   g633(.A1(new_n807_), .A2(new_n393_), .A3(new_n376_), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n835_), .A2(new_n356_), .A3(new_n284_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n547_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n511_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(KEYINPUT120), .B(G148gat), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n839_), .B(new_n840_), .ZN(G1345gat));
  NAND2_X1  g640(.A1(new_n836_), .A2(new_n563_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(KEYINPUT121), .ZN(new_n843_));
  XOR2_X1   g642(.A(KEYINPUT61), .B(G155gat), .Z(new_n844_));
  XNOR2_X1  g643(.A(new_n843_), .B(new_n844_), .ZN(G1346gat));
  AOI21_X1  g644(.A(G162gat), .B1(new_n836_), .B2(new_n610_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n645_), .A2(G162gat), .ZN(new_n847_));
  XOR2_X1   g646(.A(new_n847_), .B(KEYINPUT122), .Z(new_n848_));
  AOI21_X1  g647(.A(new_n846_), .B1(new_n836_), .B2(new_n848_), .ZN(G1347gat));
  NOR2_X1   g648(.A1(new_n284_), .A2(new_n356_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n393_), .ZN(new_n851_));
  XOR2_X1   g650(.A(new_n851_), .B(KEYINPUT123), .Z(new_n852_));
  NOR3_X1   g651(.A1(new_n793_), .A2(new_n375_), .A3(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n236_), .B1(new_n853_), .B2(new_n547_), .ZN(new_n854_));
  OR2_X1    g653(.A1(new_n854_), .A2(KEYINPUT62), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(KEYINPUT62), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n853_), .A2(new_n547_), .A3(new_n231_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n855_), .A2(new_n856_), .A3(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT124), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n855_), .A2(KEYINPUT124), .A3(new_n856_), .A4(new_n857_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(G1348gat));
  NOR3_X1   g661(.A1(new_n852_), .A2(new_n807_), .A3(new_n375_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n863_), .A2(G176gat), .A3(new_n511_), .ZN(new_n864_));
  XOR2_X1   g663(.A(new_n864_), .B(KEYINPUT125), .Z(new_n865_));
  AOI21_X1  g664(.A(G176gat), .B1(new_n853_), .B2(new_n511_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n865_), .A2(new_n866_), .ZN(G1349gat));
  AOI21_X1  g666(.A(G183gat), .B1(new_n863_), .B2(new_n563_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n564_), .A2(new_n240_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n868_), .B1(new_n853_), .B2(new_n869_), .ZN(G1350gat));
  NAND3_X1  g669(.A1(new_n853_), .A2(new_n241_), .A3(new_n610_), .ZN(new_n871_));
  AND2_X1   g670(.A1(new_n853_), .A2(new_n645_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n871_), .B1(new_n872_), .B2(new_n222_), .ZN(G1351gat));
  NAND2_X1  g672(.A1(new_n835_), .A2(new_n850_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n874_), .A2(new_n548_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(new_n212_), .ZN(G1352gat));
  NOR2_X1   g675(.A1(new_n874_), .A2(new_n510_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(new_n206_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n878_), .B1(new_n209_), .B2(new_n877_), .ZN(G1353gat));
  NOR2_X1   g678(.A1(new_n874_), .A2(new_n564_), .ZN(new_n880_));
  XOR2_X1   g679(.A(KEYINPUT63), .B(G211gat), .Z(new_n881_));
  AND2_X1   g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(KEYINPUT126), .ZN(new_n883_));
  OR2_X1    g682(.A1(new_n882_), .A2(KEYINPUT126), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n880_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n883_), .B1(new_n884_), .B2(new_n885_), .ZN(G1354gat));
  INV_X1    g685(.A(new_n874_), .ZN(new_n887_));
  AOI21_X1  g686(.A(G218gat), .B1(new_n887_), .B2(new_n610_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n645_), .A2(G218gat), .ZN(new_n889_));
  XOR2_X1   g688(.A(new_n889_), .B(KEYINPUT127), .Z(new_n890_));
  AOI21_X1  g689(.A(new_n888_), .B1(new_n887_), .B2(new_n890_), .ZN(G1355gat));
endmodule


