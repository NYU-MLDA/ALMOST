//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 1 1 0 0 0 1 0 0 0 0 1 1 1 0 0 1 1 1 0 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 0 0 0 1 0 1 0 1 1 1 1 0 0 1 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n678_, new_n679_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n726_, new_n727_, new_n728_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n859_, new_n860_, new_n862_, new_n863_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n897_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_, new_n910_,
    new_n911_;
  XNOR2_X1  g000(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G226gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G169gat), .ZN(new_n205_));
  INV_X1    g004(.A(G176gat), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT24), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208_));
  MUX2_X1   g007(.A(new_n207_), .B(KEYINPUT24), .S(new_n208_), .Z(new_n209_));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT23), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT25), .B(G183gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n212_), .A2(KEYINPUT79), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT26), .B(G190gat), .ZN(new_n214_));
  INV_X1    g013(.A(G183gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT79), .B1(new_n215_), .B2(KEYINPUT25), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n209_), .B(new_n211_), .C1(new_n213_), .C2(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n211_), .B1(G183gat), .B2(G190gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n205_), .A2(new_n206_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT22), .B(G169gat), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n220_), .B1(new_n221_), .B2(new_n206_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n219_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n218_), .A2(new_n223_), .ZN(new_n224_));
  XOR2_X1   g023(.A(G197gat), .B(G204gat), .Z(new_n225_));
  INV_X1    g024(.A(KEYINPUT86), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(new_n226_), .A3(KEYINPUT21), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G211gat), .B(G218gat), .ZN(new_n228_));
  OAI211_X1 g027(.A(new_n227_), .B(new_n228_), .C1(KEYINPUT21), .C2(new_n225_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n228_), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n230_), .A2(new_n225_), .A3(new_n226_), .A4(KEYINPUT21), .ZN(new_n231_));
  AND3_X1   g030(.A1(new_n229_), .A2(KEYINPUT87), .A3(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(KEYINPUT87), .B1(new_n229_), .B2(new_n231_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n224_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n229_), .A2(new_n231_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n212_), .A2(new_n214_), .ZN(new_n239_));
  AND2_X1   g038(.A1(new_n239_), .A2(new_n211_), .ZN(new_n240_));
  AOI22_X1  g039(.A1(new_n240_), .A2(new_n209_), .B1(new_n219_), .B2(new_n222_), .ZN(new_n241_));
  OAI21_X1  g040(.A(KEYINPUT20), .B1(new_n238_), .B2(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n204_), .B1(new_n236_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT20), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n244_), .B1(new_n238_), .B2(new_n241_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n204_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n233_), .A2(new_n235_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n224_), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n245_), .B(new_n246_), .C1(new_n247_), .C2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n243_), .A2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G8gat), .B(G36gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT18), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G64gat), .B(G92gat), .ZN(new_n253_));
  XOR2_X1   g052(.A(new_n252_), .B(new_n253_), .Z(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n250_), .A2(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n243_), .A2(new_n249_), .A3(new_n254_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT98), .B(KEYINPUT27), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n246_), .B1(new_n236_), .B2(new_n242_), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n204_), .B(new_n245_), .C1(new_n247_), .C2(new_n248_), .ZN(new_n262_));
  AND2_X1   g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(new_n255_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n264_), .A2(KEYINPUT27), .A3(new_n257_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n260_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(G155gat), .A2(G162gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G155gat), .A2(G162gat), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n268_), .B1(KEYINPUT1), .B2(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n270_), .B1(KEYINPUT1), .B2(new_n269_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G141gat), .A2(G148gat), .ZN(new_n272_));
  INV_X1    g071(.A(G141gat), .ZN(new_n273_));
  INV_X1    g072(.A(G148gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n271_), .A2(new_n272_), .A3(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT83), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT3), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n278_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT2), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n272_), .A2(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n282_));
  OAI21_X1  g081(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n279_), .A2(new_n281_), .A3(new_n282_), .A4(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT82), .ZN(new_n285_));
  AND3_X1   g084(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n286_));
  AOI21_X1  g085(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT82), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n288_), .A2(new_n289_), .A3(new_n283_), .A4(new_n279_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n285_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n269_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n292_), .A2(new_n268_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n277_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n293_), .ZN(new_n295_));
  AOI211_X1 g094(.A(KEYINPUT83), .B(new_n295_), .C1(new_n285_), .C2(new_n290_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n276_), .B1(new_n294_), .B2(new_n296_), .ZN(new_n297_));
  XOR2_X1   g096(.A(G127gat), .B(G134gat), .Z(new_n298_));
  XNOR2_X1  g097(.A(G113gat), .B(G120gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  XOR2_X1   g099(.A(new_n297_), .B(new_n300_), .Z(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT4), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT4), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n297_), .A2(new_n303_), .A3(new_n300_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G225gat), .A2(G233gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(KEYINPUT93), .ZN(new_n306_));
  XOR2_X1   g105(.A(new_n306_), .B(KEYINPUT94), .Z(new_n307_));
  NAND3_X1  g106(.A1(new_n302_), .A2(new_n304_), .A3(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n301_), .A2(new_n306_), .ZN(new_n309_));
  XOR2_X1   g108(.A(G1gat), .B(G29gat), .Z(new_n310_));
  XNOR2_X1  g109(.A(G57gat), .B(G85gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(KEYINPUT95), .B(KEYINPUT0), .Z(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  AND3_X1   g114(.A1(new_n308_), .A2(new_n309_), .A3(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n315_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT97), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NOR3_X1   g119(.A1(new_n316_), .A2(new_n317_), .A3(KEYINPUT97), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n267_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT85), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n297_), .A2(new_n323_), .A3(KEYINPUT29), .ZN(new_n324_));
  AND2_X1   g123(.A1(G228gat), .A2(G233gat), .ZN(new_n325_));
  NOR3_X1   g124(.A1(new_n232_), .A2(new_n234_), .A3(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n324_), .A2(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n323_), .B1(new_n297_), .B2(KEYINPUT29), .ZN(new_n328_));
  OAI21_X1  g127(.A(KEYINPUT88), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n297_), .A2(KEYINPUT29), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT85), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT88), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n331_), .A2(new_n332_), .A3(new_n324_), .A4(new_n326_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n329_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT89), .ZN(new_n335_));
  AND3_X1   g134(.A1(new_n297_), .A2(new_n335_), .A3(KEYINPUT29), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n335_), .B1(new_n297_), .B2(KEYINPUT29), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n237_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(new_n325_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n334_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT90), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G78gat), .B(G106gat), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n340_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  AOI22_X1  g142(.A1(new_n329_), .A2(new_n333_), .B1(new_n338_), .B2(new_n325_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n342_), .ZN(new_n345_));
  OAI21_X1  g144(.A(KEYINPUT90), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(new_n345_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n343_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(KEYINPUT84), .ZN(new_n349_));
  OR2_X1    g148(.A1(new_n297_), .A2(KEYINPUT29), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT28), .ZN(new_n351_));
  XOR2_X1   g150(.A(G22gat), .B(G50gat), .Z(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n349_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT84), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n348_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n352_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n351_), .B(new_n357_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n345_), .A2(KEYINPUT91), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n344_), .A2(new_n360_), .ZN(new_n361_));
  AND3_X1   g160(.A1(new_n334_), .A2(new_n339_), .A3(new_n360_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n358_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n356_), .A2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n300_), .B(KEYINPUT31), .ZN(new_n366_));
  XOR2_X1   g165(.A(new_n224_), .B(KEYINPUT30), .Z(new_n367_));
  XOR2_X1   g166(.A(G15gat), .B(G43gat), .Z(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT80), .ZN(new_n369_));
  XOR2_X1   g168(.A(G71gat), .B(G99gat), .Z(new_n370_));
  NAND2_X1  g169(.A1(G227gat), .A2(G233gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n369_), .B(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n367_), .B(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n366_), .B1(new_n374_), .B2(KEYINPUT81), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n375_), .B1(KEYINPUT81), .B2(new_n374_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n374_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT81), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n377_), .A2(new_n378_), .A3(new_n366_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n376_), .A2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n354_), .A2(new_n365_), .A3(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n380_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n363_), .B1(new_n355_), .B2(new_n348_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n358_), .B1(new_n348_), .B2(KEYINPUT84), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n382_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n322_), .B1(new_n381_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n250_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n254_), .A2(KEYINPUT32), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(KEYINPUT96), .ZN(new_n389_));
  INV_X1    g188(.A(new_n388_), .ZN(new_n390_));
  AOI22_X1  g189(.A1(new_n387_), .A2(new_n389_), .B1(new_n263_), .B2(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n391_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n302_), .A2(new_n306_), .A3(new_n304_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n315_), .B1(new_n301_), .B2(new_n307_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n258_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n308_), .A2(KEYINPUT33), .A3(new_n309_), .A4(new_n315_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n316_), .A2(KEYINPUT33), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n392_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n380_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n400_), .B1(new_n354_), .B2(new_n365_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n386_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(KEYINPUT64), .A2(KEYINPUT6), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(KEYINPUT64), .A2(KEYINPUT6), .ZN(new_n405_));
  OAI211_X1 g204(.A(G99gat), .B(G106gat), .C1(new_n404_), .C2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT64), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT6), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(G99gat), .ZN(new_n410_));
  INV_X1    g209(.A(G106gat), .ZN(new_n411_));
  OAI211_X1 g210(.A(new_n409_), .B(new_n403_), .C1(new_n410_), .C2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n406_), .A2(new_n412_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n414_));
  NAND2_X1  g213(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n415_));
  NOR2_X1   g214(.A1(G99gat), .A2(G106gat), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n414_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n416_), .A2(new_n414_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n413_), .A2(new_n419_), .ZN(new_n420_));
  XOR2_X1   g219(.A(G85gat), .B(G92gat), .Z(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT8), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT8), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n420_), .A2(new_n424_), .A3(new_n421_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n423_), .A2(KEYINPUT69), .A3(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT69), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n424_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n421_), .ZN(new_n429_));
  AOI211_X1 g228(.A(KEYINPUT8), .B(new_n429_), .C1(new_n413_), .C2(new_n419_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n427_), .B1(new_n428_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(G85gat), .ZN(new_n432_));
  INV_X1    g231(.A(G92gat), .ZN(new_n433_));
  NOR3_X1   g232(.A1(new_n432_), .A2(new_n433_), .A3(KEYINPUT9), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n434_), .B1(new_n421_), .B2(KEYINPUT9), .ZN(new_n435_));
  XOR2_X1   g234(.A(KEYINPUT10), .B(G99gat), .Z(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(new_n411_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n435_), .A2(new_n413_), .A3(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n426_), .A2(new_n431_), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT11), .ZN(new_n440_));
  INV_X1    g239(.A(G64gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(G57gat), .ZN(new_n442_));
  INV_X1    g241(.A(G57gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(G64gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT67), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT67), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n442_), .A2(new_n444_), .A3(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n440_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n449_));
  AND3_X1   g248(.A1(new_n442_), .A2(new_n444_), .A3(new_n447_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n447_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n451_));
  NOR3_X1   g250(.A1(new_n450_), .A2(new_n451_), .A3(KEYINPUT11), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT68), .ZN(new_n453_));
  NOR2_X1   g252(.A1(KEYINPUT66), .A2(G71gat), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(G78gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(KEYINPUT66), .A2(G71gat), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n455_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n457_), .ZN(new_n459_));
  OAI21_X1  g258(.A(G78gat), .B1(new_n459_), .B2(new_n454_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n458_), .A2(new_n460_), .ZN(new_n461_));
  NOR3_X1   g260(.A1(new_n452_), .A2(new_n453_), .A3(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n461_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n446_), .A2(new_n440_), .A3(new_n448_), .ZN(new_n464_));
  AOI21_X1  g263(.A(KEYINPUT68), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n449_), .B1(new_n462_), .B2(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n453_), .B1(new_n452_), .B2(new_n461_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n463_), .A2(new_n464_), .A3(KEYINPUT68), .ZN(new_n468_));
  INV_X1    g267(.A(new_n449_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n467_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  AND2_X1   g269(.A1(new_n466_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n439_), .A2(new_n471_), .A3(KEYINPUT12), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G230gat), .A2(G233gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n466_), .A2(new_n470_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n438_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n475_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(KEYINPUT70), .B(KEYINPUT12), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n478_), .B1(new_n474_), .B2(new_n476_), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n472_), .A2(new_n473_), .A3(new_n477_), .A4(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n473_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n477_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n474_), .A2(new_n476_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n481_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G120gat), .B(G148gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT5), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G176gat), .B(G204gat), .ZN(new_n487_));
  XOR2_X1   g286(.A(new_n486_), .B(new_n487_), .Z(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n480_), .A2(new_n484_), .A3(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(KEYINPUT71), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n480_), .A2(new_n484_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(new_n488_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n491_), .B(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT13), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n491_), .A2(new_n492_), .A3(new_n488_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n493_), .A2(KEYINPUT71), .A3(new_n490_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT13), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n496_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT72), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n496_), .A2(KEYINPUT72), .A3(new_n500_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G29gat), .B(G36gat), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G43gat), .B(G50gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n508_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(new_n506_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n509_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G15gat), .B(G22gat), .ZN(new_n514_));
  INV_X1    g313(.A(G1gat), .ZN(new_n515_));
  INV_X1    g314(.A(G8gat), .ZN(new_n516_));
  OAI21_X1  g315(.A(KEYINPUT14), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n514_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G1gat), .B(G8gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n518_), .A2(new_n519_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n513_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n520_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(new_n512_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G229gat), .A2(G233gat), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT15), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n512_), .B(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(new_n523_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(new_n522_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n527_), .B1(new_n531_), .B2(new_n526_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G113gat), .B(G141gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G169gat), .B(G197gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n532_), .B(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n505_), .A2(new_n536_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n402_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n439_), .A2(new_n529_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT74), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT35), .ZN(new_n541_));
  XNOR2_X1  g340(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G232gat), .A2(G233gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  AOI22_X1  g344(.A1(new_n476_), .A2(new_n513_), .B1(new_n541_), .B2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n539_), .A2(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n545_), .A2(new_n541_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n540_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT76), .ZN(new_n550_));
  INV_X1    g349(.A(new_n548_), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n539_), .B(new_n546_), .C1(KEYINPUT74), .C2(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n549_), .A2(new_n550_), .A3(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G190gat), .B(G218gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT75), .ZN(new_n555_));
  XOR2_X1   g354(.A(G134gat), .B(G162gat), .Z(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n557_), .A2(KEYINPUT36), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n553_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n558_), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n549_), .A2(new_n550_), .A3(new_n560_), .A4(new_n552_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n549_), .A2(new_n552_), .ZN(new_n562_));
  AND2_X1   g361(.A1(new_n557_), .A2(KEYINPUT36), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n559_), .A2(new_n561_), .A3(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(KEYINPUT37), .ZN(new_n566_));
  AOI22_X1  g365(.A1(new_n553_), .A2(new_n558_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT37), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n567_), .A2(new_n568_), .A3(new_n561_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n566_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G231gat), .A2(G233gat), .ZN(new_n571_));
  XOR2_X1   g370(.A(new_n523_), .B(new_n571_), .Z(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(new_n474_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G127gat), .B(G155gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G183gat), .B(G211gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(KEYINPUT17), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n573_), .A2(new_n579_), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n578_), .B(KEYINPUT17), .Z(new_n581_));
  OAI21_X1  g380(.A(new_n580_), .B1(new_n573_), .B2(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n582_), .B(KEYINPUT78), .Z(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n570_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n538_), .A2(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n320_), .A2(new_n321_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NOR3_X1   g387(.A1(new_n586_), .A2(G1gat), .A3(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n589_), .B(KEYINPUT38), .Z(new_n590_));
  INV_X1    g389(.A(new_n322_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n380_), .B1(new_n354_), .B2(new_n365_), .ZN(new_n592_));
  NOR3_X1   g391(.A1(new_n383_), .A2(new_n384_), .A3(new_n382_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n591_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n354_), .A2(new_n365_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n595_), .A2(new_n380_), .A3(new_n399_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n594_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT99), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n565_), .A2(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n567_), .A2(KEYINPUT99), .A3(new_n561_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n536_), .ZN(new_n602_));
  AOI211_X1 g401(.A(new_n602_), .B(new_n584_), .C1(new_n503_), .C2(new_n504_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n597_), .A2(new_n601_), .A3(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(G1gat), .B1(new_n604_), .B2(new_n588_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n590_), .A2(new_n605_), .ZN(G1324gat));
  INV_X1    g405(.A(KEYINPUT40), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT102), .ZN(new_n608_));
  OAI21_X1  g407(.A(G8gat), .B1(new_n604_), .B2(new_n267_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n608_), .B1(new_n609_), .B2(KEYINPUT39), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n599_), .A2(new_n600_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n402_), .A2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n612_), .A2(new_n266_), .A3(new_n603_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT39), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n613_), .A2(KEYINPUT102), .A3(new_n614_), .A4(G8gat), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n610_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT101), .ZN(new_n617_));
  AND3_X1   g416(.A1(new_n609_), .A2(new_n617_), .A3(KEYINPUT39), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n617_), .B1(new_n609_), .B2(KEYINPUT39), .ZN(new_n619_));
  NOR3_X1   g418(.A1(new_n616_), .A2(new_n618_), .A3(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n266_), .A2(new_n516_), .ZN(new_n621_));
  OR3_X1    g420(.A1(new_n586_), .A2(KEYINPUT100), .A3(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(KEYINPUT100), .B1(new_n586_), .B2(new_n621_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n607_), .B1(new_n620_), .B2(new_n625_), .ZN(new_n626_));
  OR2_X1    g425(.A1(new_n618_), .A2(new_n619_), .ZN(new_n627_));
  OAI211_X1 g426(.A(KEYINPUT40), .B(new_n624_), .C1(new_n627_), .C2(new_n616_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(G1325gat));
  NOR3_X1   g428(.A1(new_n586_), .A2(G15gat), .A3(new_n380_), .ZN(new_n630_));
  XOR2_X1   g429(.A(new_n630_), .B(KEYINPUT103), .Z(new_n631_));
  OAI21_X1  g430(.A(G15gat), .B1(new_n604_), .B2(new_n380_), .ZN(new_n632_));
  XOR2_X1   g431(.A(new_n632_), .B(KEYINPUT41), .Z(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n633_), .ZN(G1326gat));
  XOR2_X1   g433(.A(new_n595_), .B(KEYINPUT104), .Z(new_n635_));
  OAI21_X1  g434(.A(G22gat), .B1(new_n604_), .B2(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT42), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n635_), .A2(G22gat), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT105), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n637_), .B1(new_n586_), .B2(new_n639_), .ZN(G1327gat));
  NOR2_X1   g439(.A1(new_n601_), .A2(new_n583_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n538_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(G29gat), .B1(new_n643_), .B2(new_n587_), .ZN(new_n644_));
  XOR2_X1   g443(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n645_));
  INV_X1    g444(.A(new_n570_), .ZN(new_n646_));
  OAI21_X1  g445(.A(KEYINPUT43), .B1(new_n402_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT43), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n648_), .B(new_n570_), .C1(new_n386_), .C2(new_n401_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n537_), .A2(new_n583_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n645_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(G29gat), .ZN(new_n653_));
  NOR3_X1   g452(.A1(new_n652_), .A2(new_n653_), .A3(new_n588_), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n650_), .A2(KEYINPUT44), .A3(new_n651_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n644_), .B1(new_n654_), .B2(new_n656_), .ZN(G1328gat));
  INV_X1    g456(.A(G36gat), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n266_), .A2(new_n658_), .ZN(new_n659_));
  OR3_X1    g458(.A1(new_n642_), .A2(KEYINPUT45), .A3(new_n659_), .ZN(new_n660_));
  OAI21_X1  g459(.A(KEYINPUT45), .B1(new_n642_), .B2(new_n659_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n655_), .A2(new_n652_), .A3(new_n267_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n662_), .B1(new_n663_), .B2(new_n658_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT46), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  OAI211_X1 g465(.A(KEYINPUT46), .B(new_n662_), .C1(new_n663_), .C2(new_n658_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1329gat));
  NOR2_X1   g467(.A1(new_n655_), .A2(new_n652_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n669_), .A2(G43gat), .A3(new_n382_), .ZN(new_n670_));
  INV_X1    g469(.A(G43gat), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n671_), .B1(new_n642_), .B2(new_n380_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(KEYINPUT47), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT47), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n670_), .A2(new_n675_), .A3(new_n672_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n676_), .ZN(G1330gat));
  INV_X1    g476(.A(new_n635_), .ZN(new_n678_));
  AOI21_X1  g477(.A(G50gat), .B1(new_n643_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(G50gat), .ZN(new_n680_));
  NOR3_X1   g479(.A1(new_n652_), .A2(new_n680_), .A3(new_n595_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n679_), .B1(new_n681_), .B2(new_n656_), .ZN(G1331gat));
  NOR2_X1   g481(.A1(new_n402_), .A2(new_n536_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n505_), .B1(new_n683_), .B2(KEYINPUT107), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT107), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n685_), .B1(new_n402_), .B2(new_n536_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n684_), .A2(new_n585_), .A3(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT108), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n684_), .A2(KEYINPUT108), .A3(new_n585_), .A4(new_n686_), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n689_), .A2(new_n443_), .A3(new_n587_), .A4(new_n690_), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n505_), .A2(new_n536_), .A3(new_n584_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n612_), .A2(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(G57gat), .B1(new_n693_), .B2(new_n588_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n691_), .A2(new_n694_), .ZN(G1332gat));
  OAI21_X1  g494(.A(G64gat), .B1(new_n693_), .B2(new_n267_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT48), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n266_), .A2(new_n441_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT109), .Z(new_n699_));
  NAND3_X1  g498(.A1(new_n689_), .A2(new_n690_), .A3(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n697_), .A2(new_n700_), .ZN(G1333gat));
  OAI21_X1  g500(.A(G71gat), .B1(new_n693_), .B2(new_n380_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT49), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n380_), .A2(G71gat), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n689_), .A2(new_n690_), .A3(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT110), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n703_), .A2(new_n705_), .A3(KEYINPUT110), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1334gat));
  NAND4_X1  g509(.A1(new_n689_), .A2(new_n456_), .A3(new_n678_), .A4(new_n690_), .ZN(new_n711_));
  OAI21_X1  g510(.A(G78gat), .B1(new_n693_), .B2(new_n635_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT50), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(KEYINPUT111), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT111), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n711_), .A2(new_n713_), .A3(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(G1335gat));
  NAND3_X1  g517(.A1(new_n684_), .A2(new_n641_), .A3(new_n686_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n720_), .A2(new_n432_), .A3(new_n587_), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n505_), .A2(new_n536_), .A3(new_n583_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n650_), .A2(new_n722_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n723_), .A2(new_n587_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n721_), .B1(new_n724_), .B2(new_n432_), .ZN(G1336gat));
  AOI21_X1  g524(.A(G92gat), .B1(new_n720_), .B2(new_n266_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n266_), .A2(G92gat), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT112), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n726_), .B1(new_n723_), .B2(new_n728_), .ZN(G1337gat));
  AOI21_X1  g528(.A(new_n410_), .B1(new_n723_), .B2(new_n382_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n382_), .A2(new_n436_), .ZN(new_n731_));
  OAI21_X1  g530(.A(KEYINPUT113), .B1(new_n719_), .B2(new_n731_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n730_), .A2(new_n732_), .ZN(new_n733_));
  XOR2_X1   g532(.A(KEYINPUT114), .B(KEYINPUT51), .Z(new_n734_));
  XNOR2_X1  g533(.A(new_n733_), .B(new_n734_), .ZN(G1338gat));
  INV_X1    g534(.A(new_n595_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n648_), .B1(new_n597_), .B2(new_n570_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n649_), .ZN(new_n738_));
  OAI211_X1 g537(.A(new_n736_), .B(new_n722_), .C1(new_n737_), .C2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT52), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n739_), .A2(new_n740_), .A3(G106gat), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT115), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n739_), .A2(KEYINPUT115), .A3(new_n740_), .A4(G106gat), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n739_), .A2(G106gat), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(KEYINPUT52), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n743_), .A2(new_n744_), .A3(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n720_), .A2(new_n411_), .A3(new_n736_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT53), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT53), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n747_), .A2(new_n751_), .A3(new_n748_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(G1339gat));
  NOR3_X1   g552(.A1(new_n320_), .A2(new_n321_), .A3(new_n266_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n592_), .A2(new_n754_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT121), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT119), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n490_), .A2(new_n536_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(KEYINPUT116), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT116), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n490_), .A2(new_n536_), .A3(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT117), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT55), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n480_), .A2(new_n765_), .A3(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n472_), .A2(new_n477_), .A3(new_n479_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(new_n481_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n766_), .B1(new_n480_), .B2(new_n765_), .ZN(new_n771_));
  OAI211_X1 g570(.A(KEYINPUT56), .B(new_n488_), .C1(new_n770_), .C2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n480_), .A2(new_n765_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT55), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n775_), .A2(new_n767_), .A3(new_n769_), .ZN(new_n776_));
  AOI21_X1  g575(.A(KEYINPUT56), .B1(new_n776_), .B2(new_n488_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n764_), .B1(new_n773_), .B2(new_n777_), .ZN(new_n778_));
  OR2_X1    g577(.A1(new_n532_), .A2(new_n535_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n525_), .A2(new_n526_), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n780_), .B(new_n535_), .C1(new_n531_), .C2(new_n526_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n779_), .A2(new_n781_), .ZN(new_n782_));
  AND3_X1   g581(.A1(new_n497_), .A2(new_n498_), .A3(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n611_), .B1(new_n778_), .B2(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n758_), .B1(new_n785_), .B2(KEYINPUT57), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n488_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT56), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(new_n772_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n783_), .B1(new_n790_), .B2(new_n764_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT57), .ZN(new_n792_));
  NOR4_X1   g591(.A1(new_n791_), .A2(KEYINPUT119), .A3(new_n611_), .A4(new_n792_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n782_), .A2(new_n490_), .ZN(new_n794_));
  AOI21_X1  g593(.A(KEYINPUT58), .B1(new_n790_), .B2(new_n794_), .ZN(new_n795_));
  OAI211_X1 g594(.A(KEYINPUT58), .B(new_n794_), .C1(new_n773_), .C2(new_n777_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(new_n570_), .ZN(new_n797_));
  OAI22_X1  g596(.A1(new_n786_), .A2(new_n793_), .B1(new_n795_), .B2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n785_), .A2(KEYINPUT118), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT118), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n800_), .B1(new_n791_), .B2(new_n611_), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT57), .B1(new_n799_), .B2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n584_), .B1(new_n798_), .B2(new_n802_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n585_), .A2(new_n602_), .A3(new_n500_), .A4(new_n496_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT54), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n804_), .B(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n803_), .A2(KEYINPUT120), .A3(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT120), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n797_), .A2(new_n795_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n763_), .B1(new_n789_), .B2(new_n772_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n601_), .B(KEYINPUT57), .C1(new_n783_), .C2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(KEYINPUT119), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n778_), .A2(new_n784_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n814_), .A2(new_n758_), .A3(KEYINPUT57), .A4(new_n601_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n810_), .B1(new_n813_), .B2(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(KEYINPUT118), .B1(new_n814_), .B2(new_n601_), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n791_), .A2(new_n800_), .A3(new_n611_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n792_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n583_), .B1(new_n816_), .B2(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n809_), .B1(new_n820_), .B2(new_n806_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n757_), .B1(new_n808_), .B2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(G113gat), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n822_), .A2(new_n823_), .A3(new_n536_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n803_), .A2(new_n807_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT59), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n756_), .A2(KEYINPUT122), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n756_), .A2(KEYINPUT122), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n825_), .B(new_n826_), .C1(new_n827_), .C2(new_n828_), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n536_), .B(new_n829_), .C1(new_n822_), .C2(new_n826_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n824_), .B1(new_n831_), .B2(new_n823_), .ZN(G1340gat));
  OAI21_X1  g631(.A(new_n829_), .B1(new_n822_), .B2(new_n826_), .ZN(new_n833_));
  OAI21_X1  g632(.A(G120gat), .B1(new_n833_), .B2(new_n505_), .ZN(new_n834_));
  INV_X1    g633(.A(G120gat), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n835_), .A2(KEYINPUT60), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n835_), .B1(new_n505_), .B2(KEYINPUT60), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n836_), .B1(new_n838_), .B2(KEYINPUT123), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n822_), .B(new_n839_), .C1(KEYINPUT123), .C2(new_n838_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n834_), .A2(new_n840_), .ZN(G1341gat));
  INV_X1    g640(.A(G127gat), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n584_), .A2(new_n842_), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n829_), .B(new_n843_), .C1(new_n822_), .C2(new_n826_), .ZN(new_n844_));
  AOI21_X1  g643(.A(KEYINPUT120), .B1(new_n803_), .B2(new_n807_), .ZN(new_n845_));
  NOR3_X1   g644(.A1(new_n820_), .A2(new_n809_), .A3(new_n806_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n583_), .B(new_n756_), .C1(new_n845_), .C2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n842_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n844_), .A2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(KEYINPUT124), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT124), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n844_), .A2(new_n851_), .A3(new_n848_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n852_), .ZN(G1342gat));
  AOI21_X1  g652(.A(G134gat), .B1(new_n822_), .B2(new_n611_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n833_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n570_), .A2(G134gat), .ZN(new_n856_));
  XOR2_X1   g655(.A(new_n856_), .B(KEYINPUT125), .Z(new_n857_));
  AOI21_X1  g656(.A(new_n854_), .B1(new_n855_), .B2(new_n857_), .ZN(G1343gat));
  NAND2_X1  g657(.A1(new_n808_), .A2(new_n821_), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n859_), .A2(new_n593_), .A3(new_n536_), .A4(new_n754_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g660(.A(new_n505_), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n859_), .A2(new_n593_), .A3(new_n862_), .A4(new_n754_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(G148gat), .ZN(G1345gat));
  NAND4_X1  g663(.A1(new_n859_), .A2(new_n593_), .A3(new_n583_), .A4(new_n754_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(KEYINPUT61), .B(G155gat), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n865_), .B(new_n866_), .ZN(G1346gat));
  INV_X1    g666(.A(new_n859_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n868_), .A2(new_n381_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n869_), .A2(new_n570_), .A3(new_n754_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(G162gat), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n601_), .A2(G162gat), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n869_), .A2(new_n754_), .A3(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n871_), .A2(new_n873_), .ZN(G1347gat));
  INV_X1    g673(.A(KEYINPUT62), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n587_), .A2(new_n267_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n382_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n678_), .A2(new_n877_), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n825_), .A2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n536_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n875_), .B1(new_n880_), .B2(G169gat), .ZN(new_n881_));
  AOI211_X1 g680(.A(KEYINPUT62), .B(new_n205_), .C1(new_n879_), .C2(new_n536_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n221_), .ZN(new_n883_));
  OAI22_X1  g682(.A1(new_n881_), .A2(new_n882_), .B1(new_n883_), .B2(new_n880_), .ZN(G1348gat));
  AOI21_X1  g683(.A(G176gat), .B1(new_n879_), .B2(new_n862_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n868_), .A2(new_n736_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n877_), .A2(new_n505_), .A3(new_n206_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n885_), .B1(new_n886_), .B2(new_n887_), .ZN(G1349gat));
  NAND4_X1  g687(.A1(new_n886_), .A2(new_n382_), .A3(new_n583_), .A4(new_n876_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n584_), .A2(new_n212_), .ZN(new_n890_));
  AOI22_X1  g689(.A1(new_n889_), .A2(new_n215_), .B1(new_n879_), .B2(new_n890_), .ZN(G1350gat));
  NAND3_X1  g690(.A1(new_n879_), .A2(new_n214_), .A3(new_n611_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n825_), .A2(new_n878_), .ZN(new_n893_));
  OAI21_X1  g692(.A(G190gat), .B1(new_n893_), .B2(new_n646_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n894_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(KEYINPUT126), .ZN(G1351gat));
  NAND4_X1  g695(.A1(new_n859_), .A2(new_n593_), .A3(new_n536_), .A4(new_n876_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(G197gat), .ZN(G1352gat));
  NAND4_X1  g697(.A1(new_n859_), .A2(new_n593_), .A3(new_n862_), .A4(new_n876_), .ZN(new_n899_));
  INV_X1    g698(.A(G204gat), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n899_), .A2(KEYINPUT127), .A3(new_n900_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(KEYINPUT127), .B(G204gat), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n901_), .B1(new_n899_), .B2(new_n902_), .ZN(G1353gat));
  NAND4_X1  g702(.A1(new_n859_), .A2(new_n593_), .A3(new_n583_), .A4(new_n876_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n904_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n905_));
  XOR2_X1   g704(.A(KEYINPUT63), .B(G211gat), .Z(new_n906_));
  OAI21_X1  g705(.A(new_n905_), .B1(new_n904_), .B2(new_n906_), .ZN(G1354gat));
  NAND3_X1  g706(.A1(new_n869_), .A2(new_n570_), .A3(new_n876_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(G218gat), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n601_), .A2(G218gat), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n869_), .A2(new_n876_), .A3(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n909_), .A2(new_n911_), .ZN(G1355gat));
endmodule


