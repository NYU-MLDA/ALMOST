//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 1 0 0 1 0 1 0 0 1 1 1 0 0 1 1 0 1 0 0 0 1 1 1 1 1 0 0 1 0 1 0 1 1 1 0 0 0 0 0 0 1 1 0 1 0 1 1 1 1 1 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n775_, new_n776_, new_n777_,
    new_n779_, new_n780_, new_n781_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n793_, new_n794_, new_n795_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n824_, new_n825_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n938_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n947_, new_n948_, new_n949_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n961_, new_n962_, new_n964_, new_n965_,
    new_n966_, new_n967_, new_n969_, new_n970_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n980_,
    new_n981_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n989_, new_n990_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(G113gat), .B(G141gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT76), .ZN(new_n204_));
  XOR2_X1   g003(.A(G169gat), .B(G197gat), .Z(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G15gat), .B(G22gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G1gat), .A2(G8gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT14), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(G8gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n202_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(new_n209_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n211_), .A2(new_n214_), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n208_), .A2(new_n209_), .A3(new_n210_), .A4(new_n213_), .ZN(new_n216_));
  AND2_X1   g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  XOR2_X1   g016(.A(G29gat), .B(G36gat), .Z(new_n218_));
  OR2_X1    g017(.A1(G43gat), .A2(G50gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G43gat), .A2(G50gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n218_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT74), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G29gat), .B(G36gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n224_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n222_), .A2(new_n223_), .A3(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n223_), .B1(new_n222_), .B2(new_n225_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n217_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n222_), .A2(new_n225_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT74), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n215_), .A2(new_n216_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n231_), .A2(new_n232_), .A3(new_n226_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G229gat), .A2(G233gat), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  AND3_X1   g034(.A1(new_n229_), .A2(new_n233_), .A3(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n230_), .A2(KEYINPUT15), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT15), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n222_), .A2(new_n238_), .A3(new_n225_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n237_), .A2(new_n232_), .A3(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n235_), .B1(new_n229_), .B2(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n236_), .A2(new_n241_), .ZN(new_n242_));
  AND2_X1   g041(.A1(new_n242_), .A2(KEYINPUT75), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n242_), .A2(KEYINPUT75), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n207_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n206_), .B1(new_n236_), .B2(new_n241_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT77), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  OAI211_X1 g047(.A(KEYINPUT77), .B(new_n206_), .C1(new_n236_), .C2(new_n241_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n245_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT83), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT26), .B(G190gat), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT78), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT25), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n254_), .B1(new_n255_), .B2(G183gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT25), .B(G183gat), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n253_), .B(new_n256_), .C1(new_n257_), .C2(new_n254_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G183gat), .A2(G190gat), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT23), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  AND2_X1   g060(.A1(KEYINPUT80), .A2(KEYINPUT23), .ZN(new_n262_));
  NOR2_X1   g061(.A1(KEYINPUT80), .A2(KEYINPUT23), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n261_), .B1(new_n264_), .B2(new_n259_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT24), .ZN(new_n266_));
  INV_X1    g065(.A(G169gat), .ZN(new_n267_));
  INV_X1    g066(.A(G176gat), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n266_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G169gat), .A2(G176gat), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT79), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(KEYINPUT79), .A2(G169gat), .A3(G176gat), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n271_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n258_), .A2(new_n265_), .A3(new_n269_), .A4(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(G183gat), .ZN(new_n278_));
  INV_X1    g077(.A(G190gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NOR3_X1   g079(.A1(new_n262_), .A2(new_n263_), .A3(new_n259_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n259_), .A2(KEYINPUT23), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n280_), .B1(new_n281_), .B2(new_n283_), .ZN(new_n284_));
  AND3_X1   g083(.A1(KEYINPUT79), .A2(G169gat), .A3(G176gat), .ZN(new_n285_));
  AOI21_X1  g084(.A(KEYINPUT79), .B1(G169gat), .B2(G176gat), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n267_), .A2(KEYINPUT22), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT22), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(G169gat), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n288_), .A2(new_n290_), .A3(new_n268_), .ZN(new_n291_));
  AND2_X1   g090(.A1(new_n287_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n284_), .A2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n277_), .A2(new_n293_), .A3(KEYINPUT30), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(KEYINPUT30), .B1(new_n277_), .B2(new_n293_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G227gat), .A2(G233gat), .ZN(new_n297_));
  INV_X1    g096(.A(G15gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G71gat), .B(G99gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(G43gat), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n301_), .A2(G43gat), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n300_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n304_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n306_), .A2(new_n299_), .A3(new_n302_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  NOR3_X1   g107(.A1(new_n295_), .A2(new_n296_), .A3(new_n308_), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n305_), .A2(new_n307_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n279_), .A2(KEYINPUT26), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT26), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(G190gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n256_), .A2(new_n311_), .A3(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n278_), .A2(KEYINPUT25), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n255_), .A2(G183gat), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n254_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n276_), .B1(new_n314_), .B2(new_n317_), .ZN(new_n318_));
  OR2_X1    g117(.A1(KEYINPUT80), .A2(KEYINPUT23), .ZN(new_n319_));
  NAND2_X1  g118(.A1(KEYINPUT80), .A2(KEYINPUT23), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n319_), .A2(new_n259_), .A3(new_n320_), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n321_), .B(new_n269_), .C1(new_n260_), .C2(new_n259_), .ZN(new_n322_));
  AND2_X1   g121(.A1(G183gat), .A2(G190gat), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n319_), .A2(new_n323_), .A3(new_n320_), .ZN(new_n324_));
  AOI22_X1  g123(.A1(new_n324_), .A2(new_n282_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n287_), .A2(new_n291_), .ZN(new_n326_));
  OAI22_X1  g125(.A1(new_n318_), .A2(new_n322_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT30), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n310_), .B1(new_n329_), .B2(new_n294_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n252_), .B1(new_n309_), .B2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G127gat), .B(G134gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G113gat), .B(G120gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n335_));
  XOR2_X1   g134(.A(new_n334_), .B(new_n335_), .Z(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n308_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n329_), .A2(new_n310_), .A3(new_n294_), .ZN(new_n339_));
  AOI21_X1  g138(.A(KEYINPUT82), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n331_), .B(new_n337_), .C1(new_n340_), .C2(new_n252_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n309_), .A2(new_n330_), .ZN(new_n342_));
  OAI211_X1 g141(.A(KEYINPUT83), .B(new_n336_), .C1(new_n342_), .C2(KEYINPUT82), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(G197gat), .A2(G204gat), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G197gat), .A2(G204gat), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n346_), .A2(KEYINPUT21), .A3(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT21), .ZN(new_n349_));
  INV_X1    g148(.A(new_n347_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n349_), .B1(new_n350_), .B2(new_n345_), .ZN(new_n351_));
  INV_X1    g150(.A(G218gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(G211gat), .ZN(new_n353_));
  INV_X1    g152(.A(G211gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(G218gat), .ZN(new_n355_));
  AND3_X1   g154(.A1(new_n353_), .A2(new_n355_), .A3(KEYINPUT86), .ZN(new_n356_));
  AOI21_X1  g155(.A(KEYINPUT86), .B1(new_n353_), .B2(new_n355_), .ZN(new_n357_));
  OAI211_X1 g156(.A(new_n348_), .B(new_n351_), .C1(new_n356_), .C2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n353_), .A2(new_n355_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT86), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n353_), .A2(new_n355_), .A3(KEYINPUT86), .ZN(new_n362_));
  NOR3_X1   g161(.A1(new_n350_), .A2(new_n345_), .A3(new_n349_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n361_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n358_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G228gat), .A2(G233gat), .ZN(new_n366_));
  XOR2_X1   g165(.A(new_n366_), .B(KEYINPUT85), .Z(new_n367_));
  INV_X1    g166(.A(G141gat), .ZN(new_n368_));
  INV_X1    g167(.A(G148gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT3), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(KEYINPUT3), .B1(new_n368_), .B2(new_n369_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G141gat), .A2(G148gat), .ZN(new_n374_));
  AND2_X1   g173(.A1(new_n374_), .A2(KEYINPUT2), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n374_), .A2(KEYINPUT2), .ZN(new_n376_));
  OAI22_X1  g175(.A1(new_n372_), .A2(new_n373_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  XOR2_X1   g176(.A(G155gat), .B(G162gat), .Z(new_n378_));
  INV_X1    g177(.A(G155gat), .ZN(new_n379_));
  INV_X1    g178(.A(G162gat), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT1), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT1), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n382_), .A2(G155gat), .A3(G162gat), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n381_), .B(new_n383_), .C1(G155gat), .C2(G162gat), .ZN(new_n384_));
  AND2_X1   g183(.A1(new_n370_), .A2(new_n374_), .ZN(new_n385_));
  AOI22_X1  g184(.A1(new_n377_), .A2(new_n378_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT29), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n365_), .B(new_n367_), .C1(new_n386_), .C2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT87), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n365_), .A2(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n358_), .A2(KEYINPUT87), .A3(new_n364_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n377_), .A2(new_n378_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n384_), .A2(new_n385_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  AOI22_X1  g193(.A1(new_n390_), .A2(new_n391_), .B1(KEYINPUT29), .B2(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n388_), .B1(new_n395_), .B2(new_n367_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G78gat), .B(G106gat), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n398_), .A2(KEYINPUT88), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n396_), .A2(new_n399_), .ZN(new_n400_));
  OAI221_X1 g199(.A(new_n388_), .B1(KEYINPUT88), .B2(new_n398_), .C1(new_n395_), .C2(new_n367_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n392_), .A2(new_n387_), .A3(new_n393_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT28), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT28), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n386_), .A2(new_n404_), .A3(new_n387_), .ZN(new_n405_));
  XOR2_X1   g204(.A(G22gat), .B(G50gat), .Z(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n403_), .A2(new_n405_), .A3(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n407_), .B1(new_n403_), .B2(new_n405_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n400_), .A2(new_n401_), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n396_), .A2(new_n398_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT84), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n414_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n415_));
  OAI211_X1 g214(.A(new_n388_), .B(new_n397_), .C1(new_n395_), .C2(new_n367_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n403_), .A2(new_n405_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(new_n406_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n418_), .A2(KEYINPUT84), .A3(new_n408_), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n413_), .A2(new_n415_), .A3(new_n416_), .A4(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n344_), .A2(new_n412_), .A3(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n334_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n394_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n386_), .A2(new_n334_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n424_), .A2(KEYINPUT4), .A3(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G225gat), .A2(G233gat), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  OR3_X1    g227(.A1(new_n386_), .A2(KEYINPUT4), .A3(new_n334_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n426_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n424_), .A2(new_n425_), .A3(new_n427_), .ZN(new_n431_));
  XOR2_X1   g230(.A(G1gat), .B(G29gat), .Z(new_n432_));
  XNOR2_X1  g231(.A(G57gat), .B(G85gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n432_), .B(new_n433_), .ZN(new_n434_));
  XOR2_X1   g233(.A(KEYINPUT96), .B(KEYINPUT0), .Z(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(KEYINPUT97), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n434_), .B(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n430_), .A2(new_n431_), .A3(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT33), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT33), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n430_), .A2(new_n440_), .A3(new_n431_), .A4(new_n437_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n426_), .A2(new_n427_), .A3(new_n429_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n437_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n424_), .A2(new_n425_), .A3(new_n428_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n443_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT98), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n443_), .A2(KEYINPUT98), .A3(new_n444_), .A4(new_n445_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n442_), .A2(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G8gat), .B(G36gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n452_), .B(KEYINPUT18), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G64gat), .B(G92gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n272_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n269_), .B1(new_n456_), .B2(new_n270_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n457_), .B1(new_n282_), .B2(new_n324_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n315_), .A2(new_n316_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT92), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT92), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n315_), .A2(new_n316_), .A3(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n460_), .A2(new_n253_), .A3(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n458_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT93), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT93), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n458_), .A2(new_n463_), .A3(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n465_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n365_), .ZN(new_n469_));
  OAI211_X1 g268(.A(new_n321_), .B(new_n280_), .C1(new_n260_), .C2(new_n259_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT94), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n265_), .A2(KEYINPUT94), .A3(new_n280_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n472_), .A2(new_n473_), .A3(new_n292_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n468_), .A2(new_n469_), .A3(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n327_), .A2(new_n365_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G226gat), .A2(G233gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT90), .ZN(new_n478_));
  XOR2_X1   g277(.A(KEYINPUT89), .B(KEYINPUT19), .Z(new_n479_));
  XOR2_X1   g278(.A(new_n478_), .B(new_n479_), .Z(new_n480_));
  AND3_X1   g279(.A1(new_n476_), .A2(KEYINPUT20), .A3(new_n480_), .ZN(new_n481_));
  AND3_X1   g280(.A1(new_n458_), .A2(new_n466_), .A3(new_n463_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n466_), .B1(new_n458_), .B2(new_n463_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n474_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(new_n365_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT91), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n486_), .B(KEYINPUT20), .C1(new_n327_), .C2(new_n365_), .ZN(new_n487_));
  OAI21_X1  g286(.A(KEYINPUT20), .B1(new_n327_), .B2(new_n365_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT91), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n485_), .A2(new_n487_), .A3(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n480_), .ZN(new_n491_));
  AOI221_X4 g290(.A(new_n455_), .B1(new_n475_), .B2(new_n481_), .C1(new_n490_), .C2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n455_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n489_), .A2(new_n487_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n469_), .B1(new_n468_), .B2(new_n474_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n491_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n475_), .A2(new_n481_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n493_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT95), .B1(new_n492_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n487_), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n277_), .A2(new_n293_), .A3(new_n364_), .A4(new_n358_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n486_), .B1(new_n501_), .B2(KEYINPUT20), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n500_), .A2(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n480_), .B1(new_n503_), .B2(new_n485_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n497_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n455_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT95), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n496_), .A2(new_n497_), .A3(new_n493_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n506_), .A2(new_n507_), .A3(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n451_), .B1(new_n499_), .B2(new_n509_), .ZN(new_n510_));
  AND4_X1   g309(.A1(new_n474_), .A2(new_n390_), .A3(new_n464_), .A4(new_n391_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n476_), .A2(KEYINPUT20), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  MUX2_X1   g312(.A(new_n513_), .B(new_n490_), .S(new_n480_), .Z(new_n514_));
  NAND3_X1  g313(.A1(new_n514_), .A2(KEYINPUT32), .A3(new_n493_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n493_), .A2(KEYINPUT32), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n516_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n438_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n437_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n518_), .B1(KEYINPUT99), .B2(new_n519_), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n519_), .A2(KEYINPUT99), .ZN(new_n521_));
  AOI22_X1  g320(.A1(new_n515_), .A2(new_n517_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n422_), .B1(new_n510_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n420_), .A2(new_n412_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(new_n344_), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n420_), .A2(new_n341_), .A3(new_n412_), .A4(new_n343_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT27), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n528_), .B1(new_n492_), .B2(new_n498_), .ZN(new_n529_));
  OAI211_X1 g328(.A(KEYINPUT27), .B(new_n508_), .C1(new_n514_), .C2(new_n493_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n519_), .A2(KEYINPUT99), .ZN(new_n531_));
  AND3_X1   g330(.A1(new_n521_), .A2(new_n531_), .A3(new_n438_), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n527_), .A2(new_n529_), .A3(new_n530_), .A4(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n523_), .A2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G190gat), .B(G218gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G134gat), .B(G162gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  XOR2_X1   g336(.A(new_n537_), .B(KEYINPUT36), .Z(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(KEYINPUT10), .B(G99gat), .Z(new_n540_));
  INV_X1    g339(.A(G106gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  AND3_X1   g341(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n543_));
  AOI21_X1  g342(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n542_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT9), .ZN(new_n548_));
  XNOR2_X1  g347(.A(KEYINPUT64), .B(G85gat), .ZN(new_n549_));
  INV_X1    g348(.A(G92gat), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n548_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(G85gat), .A2(G92gat), .ZN(new_n552_));
  AND2_X1   g351(.A1(G85gat), .A2(G92gat), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n552_), .B1(new_n553_), .B2(KEYINPUT9), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n551_), .A2(KEYINPUT65), .A3(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(KEYINPUT65), .B1(new_n551_), .B2(new_n554_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n547_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n553_), .A2(new_n552_), .ZN(new_n559_));
  INV_X1    g358(.A(G99gat), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n560_), .A2(new_n541_), .A3(KEYINPUT7), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT7), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n562_), .B1(G99gat), .B2(G106gat), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n559_), .B1(new_n564_), .B2(new_n545_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n553_), .A2(new_n552_), .ZN(new_n566_));
  AOI21_X1  g365(.A(KEYINPUT8), .B1(new_n566_), .B2(KEYINPUT66), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n565_), .B(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n558_), .A2(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n569_), .A2(new_n237_), .A3(new_n239_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n558_), .A2(new_n568_), .A3(new_n222_), .A4(new_n225_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G232gat), .A2(G233gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT34), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT35), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n570_), .A2(new_n571_), .A3(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n574_), .A2(new_n575_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n578_), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n570_), .A2(new_n580_), .A3(new_n571_), .A4(new_n576_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n539_), .B1(new_n579_), .B2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n537_), .A2(KEYINPUT36), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n579_), .A2(new_n584_), .A3(new_n581_), .ZN(new_n585_));
  AND3_X1   g384(.A1(new_n583_), .A2(KEYINPUT103), .A3(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(KEYINPUT103), .B1(new_n583_), .B2(new_n585_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n534_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(G230gat), .A2(G233gat), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(G64gat), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(G57gat), .ZN(new_n593_));
  INV_X1    g392(.A(G57gat), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(G64gat), .ZN(new_n595_));
  AOI21_X1  g394(.A(KEYINPUT11), .B1(new_n593_), .B2(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G71gat), .B(G78gat), .ZN(new_n597_));
  OAI21_X1  g396(.A(KEYINPUT67), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  AND2_X1   g397(.A1(G71gat), .A2(G78gat), .ZN(new_n599_));
  NOR2_X1   g398(.A1(G71gat), .A2(G78gat), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT67), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G57gat), .B(G64gat), .ZN(new_n603_));
  OAI211_X1 g402(.A(new_n601_), .B(new_n602_), .C1(new_n603_), .C2(KEYINPUT11), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(KEYINPUT11), .ZN(new_n605_));
  AND3_X1   g404(.A1(new_n598_), .A2(new_n604_), .A3(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n605_), .B1(new_n598_), .B2(new_n604_), .ZN(new_n607_));
  OAI211_X1 g406(.A(new_n558_), .B(new_n568_), .C1(new_n606_), .C2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(KEYINPUT68), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n606_), .A2(new_n607_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n569_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n608_), .A2(KEYINPUT68), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n591_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT69), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT12), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n551_), .A2(new_n554_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT65), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n546_), .B1(new_n620_), .B2(new_n555_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT8), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT66), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n622_), .B1(new_n559_), .B2(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n565_), .B(new_n624_), .ZN(new_n625_));
  OAI211_X1 g424(.A(new_n610_), .B(new_n617_), .C1(new_n621_), .C2(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n615_), .A2(new_n616_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(new_n629_));
  OAI211_X1 g428(.A(new_n610_), .B(new_n627_), .C1(new_n621_), .C2(new_n625_), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n629_), .A2(new_n590_), .A3(new_n608_), .A4(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n614_), .A2(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(G120gat), .B(G148gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT5), .ZN(new_n634_));
  XNOR2_X1  g433(.A(G176gat), .B(G204gat), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n634_), .B(new_n635_), .Z(new_n636_));
  NAND2_X1  g435(.A1(new_n632_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n636_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n614_), .A2(new_n631_), .A3(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(KEYINPUT13), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT13), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n637_), .A2(new_n642_), .A3(new_n639_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT72), .ZN(new_n645_));
  NAND2_X1  g444(.A1(G231gat), .A2(G233gat), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n610_), .B(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n232_), .B(KEYINPUT70), .ZN(new_n648_));
  OR2_X1    g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT17), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n647_), .A2(new_n648_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(G127gat), .B(G155gat), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT16), .ZN(new_n653_));
  XOR2_X1   g452(.A(G183gat), .B(G211gat), .Z(new_n654_));
  XNOR2_X1  g453(.A(new_n653_), .B(new_n654_), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n649_), .A2(new_n650_), .A3(new_n651_), .A4(new_n655_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n655_), .A2(new_n650_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n645_), .B1(new_n656_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n647_), .B(new_n648_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n661_), .A2(KEYINPUT71), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n656_), .A2(new_n645_), .A3(new_n658_), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n660_), .A2(new_n662_), .A3(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n662_), .B1(new_n660_), .B2(new_n663_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  AND4_X1   g466(.A1(new_n251_), .A2(new_n589_), .A3(new_n644_), .A4(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n520_), .A2(new_n521_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n202_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT37), .ZN(new_n671_));
  INV_X1    g470(.A(new_n585_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n671_), .B1(new_n672_), .B2(new_n582_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n583_), .A2(KEYINPUT37), .A3(new_n585_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n675_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT73), .Z(new_n677_));
  NAND2_X1  g476(.A1(new_n644_), .A2(new_n251_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n678_), .B1(new_n533_), .B2(new_n523_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT100), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT101), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n669_), .B(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n681_), .A2(new_n202_), .A3(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT38), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n670_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n681_), .A2(KEYINPUT38), .A3(new_n202_), .A4(new_n684_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n688_), .A2(KEYINPUT102), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n688_), .A2(KEYINPUT102), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n687_), .B1(new_n689_), .B2(new_n690_), .ZN(G1324gat));
  NAND2_X1  g490(.A1(new_n530_), .A2(new_n529_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n681_), .A2(new_n212_), .A3(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n668_), .A2(new_n692_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(G8gat), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n695_), .A2(KEYINPUT39), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n695_), .A2(KEYINPUT39), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n693_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT40), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n698_), .B(new_n699_), .ZN(G1325gat));
  INV_X1    g499(.A(new_n344_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n668_), .A2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(G15gat), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n703_), .A2(KEYINPUT41), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(KEYINPUT41), .ZN(new_n705_));
  INV_X1    g504(.A(new_n680_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n706_), .A2(new_n298_), .A3(new_n701_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n704_), .A2(new_n705_), .A3(new_n707_), .ZN(G1326gat));
  INV_X1    g507(.A(G22gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n709_), .B1(new_n668_), .B2(new_n524_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(KEYINPUT104), .B(KEYINPUT42), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n710_), .B(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n706_), .A2(new_n709_), .A3(new_n524_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1327gat));
  NOR2_X1   g513(.A1(new_n667_), .A2(new_n588_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n715_), .A2(new_n679_), .ZN(new_n716_));
  AOI21_X1  g515(.A(G29gat), .B1(new_n716_), .B2(new_n669_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n666_), .A2(new_n251_), .A3(new_n644_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n675_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n451_), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n492_), .A2(new_n498_), .A3(KEYINPUT95), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n507_), .B1(new_n506_), .B2(new_n508_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n721_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n515_), .A2(new_n517_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(new_n669_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n421_), .B1(new_n724_), .B2(new_n726_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n524_), .A2(new_n344_), .ZN(new_n728_));
  AOI22_X1  g527(.A1(new_n420_), .A2(new_n412_), .B1(new_n341_), .B2(new_n343_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n532_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n730_), .A2(new_n692_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n720_), .B1(new_n727_), .B2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT105), .ZN(new_n733_));
  AOI21_X1  g532(.A(KEYINPUT43), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n675_), .B1(new_n523_), .B2(new_n533_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT43), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n735_), .A2(KEYINPUT105), .A3(new_n736_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n719_), .B1(new_n734_), .B2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT44), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n738_), .A2(KEYINPUT106), .A3(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT106), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n732_), .A2(new_n733_), .A3(KEYINPUT43), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n736_), .B1(new_n735_), .B2(KEYINPUT105), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n718_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n741_), .B1(new_n744_), .B2(KEYINPUT44), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n740_), .A2(new_n745_), .ZN(new_n746_));
  OAI211_X1 g545(.A(KEYINPUT44), .B(new_n719_), .C1(new_n734_), .C2(new_n737_), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n747_), .A2(G29gat), .A3(new_n684_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n717_), .B1(new_n746_), .B2(new_n748_), .ZN(G1328gat));
  XOR2_X1   g548(.A(KEYINPUT109), .B(KEYINPUT46), .Z(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT107), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n747_), .A2(new_n692_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n745_), .B2(new_n740_), .ZN(new_n754_));
  INV_X1    g553(.A(G36gat), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n752_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n692_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n757_), .B1(new_n744_), .B2(KEYINPUT44), .ZN(new_n758_));
  AOI21_X1  g557(.A(KEYINPUT106), .B1(new_n738_), .B2(new_n739_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n744_), .A2(new_n741_), .A3(KEYINPUT44), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n758_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n761_), .A2(KEYINPUT107), .A3(G36gat), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n756_), .A2(new_n762_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n757_), .A2(G36gat), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n716_), .A2(new_n764_), .ZN(new_n765_));
  XOR2_X1   g564(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n766_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n716_), .A2(new_n764_), .A3(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n751_), .B1(new_n763_), .B2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n770_), .ZN(new_n772_));
  AOI211_X1 g571(.A(new_n772_), .B(new_n750_), .C1(new_n756_), .C2(new_n762_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n771_), .A2(new_n773_), .ZN(G1329gat));
  AOI21_X1  g573(.A(G43gat), .B1(new_n716_), .B2(new_n701_), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n747_), .A2(G43gat), .A3(new_n701_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n746_), .B2(new_n776_), .ZN(new_n777_));
  XOR2_X1   g576(.A(new_n777_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g577(.A(G50gat), .B1(new_n716_), .B2(new_n524_), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n747_), .A2(G50gat), .A3(new_n524_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n779_), .B1(new_n746_), .B2(new_n780_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT110), .ZN(G1331gat));
  NOR2_X1   g581(.A1(new_n644_), .A2(new_n251_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n589_), .A2(new_n667_), .A3(new_n783_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT112), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n785_), .A2(G57gat), .A3(new_n669_), .ZN(new_n786_));
  XOR2_X1   g585(.A(new_n786_), .B(KEYINPUT113), .Z(new_n787_));
  AND2_X1   g586(.A1(new_n783_), .A2(new_n534_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n677_), .A2(new_n788_), .ZN(new_n789_));
  XOR2_X1   g588(.A(new_n789_), .B(KEYINPUT111), .Z(new_n790_));
  AOI21_X1  g589(.A(G57gat), .B1(new_n790_), .B2(new_n684_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n787_), .A2(new_n791_), .ZN(G1332gat));
  AOI21_X1  g591(.A(new_n592_), .B1(new_n785_), .B2(new_n692_), .ZN(new_n793_));
  XOR2_X1   g592(.A(new_n793_), .B(KEYINPUT48), .Z(new_n794_));
  NAND3_X1  g593(.A1(new_n790_), .A2(new_n592_), .A3(new_n692_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(G1333gat));
  INV_X1    g595(.A(G71gat), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n797_), .B1(new_n785_), .B2(new_n701_), .ZN(new_n798_));
  XOR2_X1   g597(.A(new_n798_), .B(KEYINPUT49), .Z(new_n799_));
  NAND3_X1  g598(.A1(new_n790_), .A2(new_n797_), .A3(new_n701_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(G1334gat));
  INV_X1    g600(.A(G78gat), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n790_), .A2(new_n802_), .A3(new_n524_), .ZN(new_n803_));
  AOI211_X1 g602(.A(KEYINPUT50), .B(new_n802_), .C1(new_n785_), .C2(new_n524_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT50), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n785_), .A2(new_n524_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n805_), .B1(new_n806_), .B2(G78gat), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n803_), .B1(new_n804_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT114), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n803_), .B(KEYINPUT114), .C1(new_n804_), .C2(new_n807_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(G1335gat));
  AND2_X1   g611(.A1(new_n715_), .A2(new_n788_), .ZN(new_n813_));
  AOI21_X1  g612(.A(G85gat), .B1(new_n813_), .B2(new_n684_), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n783_), .A2(new_n666_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT115), .ZN(new_n816_));
  OR2_X1    g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n742_), .A2(new_n743_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n815_), .A2(new_n816_), .ZN(new_n819_));
  AND3_X1   g618(.A1(new_n817_), .A2(new_n818_), .A3(new_n819_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n532_), .A2(new_n549_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(KEYINPUT116), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n814_), .B1(new_n820_), .B2(new_n822_), .ZN(G1336gat));
  NAND3_X1  g622(.A1(new_n813_), .A2(new_n550_), .A3(new_n692_), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n820_), .A2(new_n692_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n824_), .B1(new_n825_), .B2(new_n550_), .ZN(G1337gat));
  AND2_X1   g625(.A1(new_n701_), .A2(new_n540_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n813_), .A2(new_n827_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n820_), .A2(new_n701_), .ZN(new_n829_));
  OAI211_X1 g628(.A(KEYINPUT117), .B(new_n828_), .C1(new_n829_), .C2(new_n560_), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n830_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g630(.A1(new_n813_), .A2(new_n541_), .A3(new_n524_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT52), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n820_), .A2(new_n524_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n833_), .B1(new_n834_), .B2(G106gat), .ZN(new_n835_));
  AOI211_X1 g634(.A(KEYINPUT52), .B(new_n541_), .C1(new_n820_), .C2(new_n524_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n832_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g637(.A1(new_n684_), .A2(new_n757_), .A3(new_n728_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n839_), .B(KEYINPUT121), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n251_), .A2(new_n639_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT55), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n631_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n629_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n630_), .A2(new_n608_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n591_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n845_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n847_), .A2(KEYINPUT55), .A3(new_n590_), .A4(new_n629_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n843_), .A2(new_n846_), .A3(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n636_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT56), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n849_), .A2(KEYINPUT56), .A3(new_n636_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n841_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n235_), .B1(new_n229_), .B2(new_n233_), .ZN(new_n855_));
  OR3_X1    g654(.A1(new_n855_), .A2(KEYINPUT118), .A3(new_n206_), .ZN(new_n856_));
  OAI21_X1  g655(.A(KEYINPUT118), .B1(new_n855_), .B2(new_n206_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n229_), .A2(new_n240_), .A3(new_n235_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n856_), .A2(new_n857_), .A3(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n250_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT119), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n250_), .A2(KEYINPUT119), .A3(new_n859_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n864_), .A2(new_n640_), .ZN(new_n865_));
  OAI211_X1 g664(.A(KEYINPUT57), .B(new_n588_), .C1(new_n854_), .C2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(KEYINPUT120), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n864_), .A2(new_n640_), .ZN(new_n868_));
  AND3_X1   g667(.A1(new_n849_), .A2(KEYINPUT56), .A3(new_n636_), .ZN(new_n869_));
  AOI21_X1  g668(.A(KEYINPUT56), .B1(new_n849_), .B2(new_n636_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n868_), .B1(new_n871_), .B2(new_n841_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT120), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n872_), .A2(new_n873_), .A3(KEYINPUT57), .A4(new_n588_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n867_), .A2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n863_), .ZN(new_n876_));
  AOI21_X1  g675(.A(KEYINPUT119), .B1(new_n250_), .B2(new_n859_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n639_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n878_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n675_), .B1(new_n879_), .B2(KEYINPUT58), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT58), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n881_), .B1(new_n871_), .B2(new_n878_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n588_), .B1(new_n854_), .B2(new_n865_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT57), .ZN(new_n884_));
  AOI22_X1  g683(.A1(new_n880_), .A2(new_n882_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n667_), .B1(new_n875_), .B2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n251_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n644_), .A2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT54), .ZN(new_n889_));
  OR3_X1    g688(.A1(new_n676_), .A2(new_n888_), .A3(new_n889_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n889_), .B1(new_n676_), .B2(new_n888_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n840_), .B1(new_n886_), .B2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(G113gat), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n894_), .A2(new_n895_), .A3(new_n251_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT59), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n894_), .A2(new_n897_), .ZN(new_n898_));
  AND3_X1   g697(.A1(new_n893_), .A2(KEYINPUT122), .A3(KEYINPUT59), .ZN(new_n899_));
  AOI21_X1  g698(.A(KEYINPUT122), .B1(new_n893_), .B2(KEYINPUT59), .ZN(new_n900_));
  OAI211_X1 g699(.A(new_n251_), .B(new_n898_), .C1(new_n899_), .C2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n896_), .B1(new_n902_), .B2(new_n895_), .ZN(G1340gat));
  INV_X1    g702(.A(new_n644_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT60), .ZN(new_n905_));
  INV_X1    g704(.A(G120gat), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n904_), .A2(new_n905_), .A3(new_n906_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n907_), .B1(new_n905_), .B2(new_n906_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n894_), .A2(new_n908_), .ZN(new_n909_));
  OAI211_X1 g708(.A(new_n904_), .B(new_n898_), .C1(new_n899_), .C2(new_n900_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n909_), .B1(new_n911_), .B2(new_n906_), .ZN(G1341gat));
  INV_X1    g711(.A(G127gat), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n666_), .A2(new_n913_), .ZN(new_n914_));
  OAI211_X1 g713(.A(new_n898_), .B(new_n914_), .C1(new_n899_), .C2(new_n900_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n913_), .B1(new_n893_), .B2(new_n666_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT123), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n915_), .A2(KEYINPUT123), .A3(new_n916_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n920_), .ZN(G1342gat));
  OR2_X1    g720(.A1(new_n893_), .A2(new_n588_), .ZN(new_n922_));
  INV_X1    g721(.A(G134gat), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT124), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n924_), .A2(new_n925_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n922_), .A2(KEYINPUT124), .A3(new_n923_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n926_), .A2(new_n927_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n899_), .A2(new_n900_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n929_), .B1(new_n897_), .B2(new_n894_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n675_), .A2(new_n923_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n928_), .B1(new_n930_), .B2(new_n931_), .ZN(G1343gat));
  OR2_X1    g731(.A1(new_n886_), .A2(new_n892_), .ZN(new_n933_));
  NOR3_X1   g732(.A1(new_n683_), .A2(new_n692_), .A3(new_n525_), .ZN(new_n934_));
  AND2_X1   g733(.A1(new_n933_), .A2(new_n934_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(new_n251_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n936_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g736(.A1(new_n935_), .A2(new_n904_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g738(.A1(new_n933_), .A2(new_n667_), .A3(new_n934_), .ZN(new_n940_));
  AND2_X1   g739(.A1(new_n940_), .A2(KEYINPUT125), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n940_), .A2(KEYINPUT125), .ZN(new_n942_));
  XNOR2_X1  g741(.A(KEYINPUT61), .B(G155gat), .ZN(new_n943_));
  OR3_X1    g742(.A1(new_n941_), .A2(new_n942_), .A3(new_n943_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n943_), .B1(new_n941_), .B2(new_n942_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n944_), .A2(new_n945_), .ZN(G1346gat));
  OAI211_X1 g745(.A(new_n935_), .B(new_n380_), .C1(new_n587_), .C2(new_n586_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n935_), .A2(new_n720_), .ZN(new_n948_));
  INV_X1    g747(.A(new_n948_), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n947_), .B1(new_n949_), .B2(new_n380_), .ZN(G1347gat));
  AND2_X1   g749(.A1(new_n933_), .A2(new_n692_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n684_), .A2(new_n526_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n951_), .A2(new_n952_), .ZN(new_n953_));
  OAI21_X1  g752(.A(G169gat), .B1(new_n953_), .B2(new_n887_), .ZN(new_n954_));
  INV_X1    g753(.A(KEYINPUT62), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n954_), .A2(new_n955_), .ZN(new_n956_));
  OAI211_X1 g755(.A(KEYINPUT62), .B(G169gat), .C1(new_n953_), .C2(new_n887_), .ZN(new_n957_));
  INV_X1    g756(.A(new_n953_), .ZN(new_n958_));
  NAND4_X1  g757(.A1(new_n958_), .A2(new_n251_), .A3(new_n288_), .A4(new_n290_), .ZN(new_n959_));
  NAND3_X1  g758(.A1(new_n956_), .A2(new_n957_), .A3(new_n959_), .ZN(G1348gat));
  AOI21_X1  g759(.A(G176gat), .B1(new_n958_), .B2(new_n904_), .ZN(new_n961_));
  NOR3_X1   g760(.A1(new_n953_), .A2(new_n268_), .A3(new_n644_), .ZN(new_n962_));
  NOR2_X1   g761(.A1(new_n961_), .A2(new_n962_), .ZN(G1349gat));
  NAND2_X1  g762(.A1(new_n278_), .A2(KEYINPUT126), .ZN(new_n964_));
  OAI21_X1  g763(.A(new_n964_), .B1(new_n953_), .B2(new_n666_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n958_), .A2(new_n667_), .ZN(new_n966_));
  OAI211_X1 g765(.A(new_n460_), .B(new_n462_), .C1(KEYINPUT126), .C2(G183gat), .ZN(new_n967_));
  OAI21_X1  g766(.A(new_n965_), .B1(new_n966_), .B2(new_n967_), .ZN(G1350gat));
  OAI21_X1  g767(.A(G190gat), .B1(new_n953_), .B2(new_n675_), .ZN(new_n969_));
  OAI21_X1  g768(.A(new_n253_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n970_));
  OAI21_X1  g769(.A(new_n969_), .B1(new_n953_), .B2(new_n970_), .ZN(G1351gat));
  XOR2_X1   g770(.A(KEYINPUT127), .B(G197gat), .Z(new_n972_));
  INV_X1    g771(.A(new_n972_), .ZN(new_n973_));
  NOR2_X1   g772(.A1(new_n525_), .A2(new_n669_), .ZN(new_n974_));
  NAND2_X1  g773(.A1(new_n951_), .A2(new_n974_), .ZN(new_n975_));
  INV_X1    g774(.A(new_n975_), .ZN(new_n976_));
  AOI21_X1  g775(.A(new_n973_), .B1(new_n976_), .B2(new_n251_), .ZN(new_n977_));
  NOR3_X1   g776(.A1(new_n975_), .A2(new_n887_), .A3(new_n972_), .ZN(new_n978_));
  NOR2_X1   g777(.A1(new_n977_), .A2(new_n978_), .ZN(G1352gat));
  OR3_X1    g778(.A1(new_n975_), .A2(G204gat), .A3(new_n644_), .ZN(new_n980_));
  OAI21_X1  g779(.A(G204gat), .B1(new_n975_), .B2(new_n644_), .ZN(new_n981_));
  NAND2_X1  g780(.A1(new_n980_), .A2(new_n981_), .ZN(G1353gat));
  INV_X1    g781(.A(KEYINPUT63), .ZN(new_n983_));
  NAND2_X1  g782(.A1(new_n983_), .A2(new_n354_), .ZN(new_n984_));
  AOI21_X1  g783(.A(new_n666_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n985_));
  NAND3_X1  g784(.A1(new_n976_), .A2(new_n984_), .A3(new_n985_), .ZN(new_n986_));
  OAI211_X1 g785(.A(new_n983_), .B(new_n354_), .C1(new_n975_), .C2(new_n666_), .ZN(new_n987_));
  AND2_X1   g786(.A1(new_n986_), .A2(new_n987_), .ZN(G1354gat));
  OAI21_X1  g787(.A(G218gat), .B1(new_n975_), .B2(new_n675_), .ZN(new_n989_));
  OAI21_X1  g788(.A(new_n352_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n990_));
  OAI21_X1  g789(.A(new_n989_), .B1(new_n975_), .B2(new_n990_), .ZN(G1355gat));
endmodule


