//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 0 1 1 1 1 1 0 0 0 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0 0 1 0 0 0 1 1 0 0 1 1 0 0 1 1 1 0 1 0 0 0 0 1 1 1 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n632_, new_n633_, new_n634_, new_n635_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n717_, new_n718_, new_n719_, new_n721_, new_n722_,
    new_n723_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n738_, new_n739_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n855_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n862_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n897_, new_n898_, new_n899_, new_n901_,
    new_n902_, new_n903_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_;
  NAND2_X1  g000(.A1(G99gat), .A2(G106gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT6), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT6), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n204_), .A2(G99gat), .A3(G106gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  XOR2_X1   g005(.A(KEYINPUT10), .B(G99gat), .Z(new_n207_));
  INV_X1    g006(.A(G106gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G85gat), .B(G92gat), .ZN(new_n210_));
  OR2_X1    g009(.A1(new_n210_), .A2(KEYINPUT9), .ZN(new_n211_));
  INV_X1    g010(.A(G92gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n210_), .B1(KEYINPUT9), .B2(new_n212_), .ZN(new_n213_));
  AND3_X1   g012(.A1(new_n211_), .A2(KEYINPUT64), .A3(new_n213_), .ZN(new_n214_));
  AOI21_X1  g013(.A(KEYINPUT64), .B1(new_n211_), .B2(new_n213_), .ZN(new_n215_));
  OAI211_X1 g014(.A(new_n206_), .B(new_n209_), .C1(new_n214_), .C2(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n217_), .B1(G99gat), .B2(G106gat), .ZN(new_n218_));
  INV_X1    g017(.A(G99gat), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n219_), .B(new_n208_), .C1(KEYINPUT65), .C2(KEYINPUT7), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(new_n206_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n210_), .ZN(new_n223_));
  OR2_X1    g022(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n224_));
  NAND2_X1  g023(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .A4(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT8), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n206_), .A2(KEYINPUT67), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT67), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n203_), .A2(new_n205_), .A3(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n228_), .A2(new_n221_), .A3(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n227_), .B1(new_n231_), .B2(new_n223_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT68), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n226_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  AOI211_X1 g033(.A(KEYINPUT68), .B(new_n227_), .C1(new_n231_), .C2(new_n223_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n216_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  XOR2_X1   g035(.A(G71gat), .B(G78gat), .Z(new_n237_));
  XNOR2_X1  g036(.A(G57gat), .B(G64gat), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n237_), .B1(KEYINPUT11), .B2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(KEYINPUT69), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT69), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n237_), .B(new_n241_), .C1(KEYINPUT11), .C2(new_n238_), .ZN(new_n242_));
  AND2_X1   g041(.A1(new_n238_), .A2(KEYINPUT11), .ZN(new_n243_));
  AND3_X1   g042(.A1(new_n240_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n243_), .B1(new_n240_), .B2(new_n242_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n236_), .A2(new_n247_), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n246_), .B(new_n216_), .C1(new_n234_), .C2(new_n235_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n248_), .A2(KEYINPUT12), .A3(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT12), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n236_), .A2(new_n247_), .A3(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G230gat), .A2(G233gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n248_), .A2(new_n249_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n254_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n255_), .A2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G120gat), .B(G148gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT5), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G176gat), .B(G204gat), .ZN(new_n262_));
  XOR2_X1   g061(.A(new_n261_), .B(new_n262_), .Z(new_n263_));
  NAND2_X1  g062(.A1(new_n259_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n263_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n255_), .A2(new_n258_), .A3(new_n265_), .ZN(new_n266_));
  AND3_X1   g065(.A1(new_n264_), .A2(KEYINPUT13), .A3(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(KEYINPUT13), .B1(new_n264_), .B2(new_n266_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(KEYINPUT70), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT70), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n271_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  XOR2_X1   g072(.A(G29gat), .B(G36gat), .Z(new_n274_));
  XOR2_X1   g073(.A(G43gat), .B(G50gat), .Z(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT15), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n236_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT74), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G232gat), .A2(G233gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT72), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT35), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n279_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n276_), .ZN(new_n286_));
  OAI211_X1 g085(.A(new_n278_), .B(new_n285_), .C1(new_n286_), .C2(new_n236_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n283_), .A2(new_n284_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G190gat), .B(G218gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT73), .ZN(new_n291_));
  XOR2_X1   g090(.A(G134gat), .B(G162gat), .Z(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT36), .ZN(new_n294_));
  AND2_X1   g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  OR2_X1    g094(.A1(new_n236_), .A2(new_n286_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n288_), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n296_), .A2(new_n297_), .A3(new_n278_), .A4(new_n285_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n289_), .A2(new_n295_), .A3(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT75), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT75), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n289_), .A2(new_n301_), .A3(new_n295_), .A4(new_n298_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n293_), .B(new_n294_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n304_), .B1(new_n289_), .B2(new_n298_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(KEYINPUT37), .B1(new_n303_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT37), .ZN(new_n308_));
  AOI211_X1 g107(.A(new_n308_), .B(new_n305_), .C1(new_n300_), .C2(new_n302_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n307_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT80), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT76), .B(G1gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(G8gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT14), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G15gat), .B(G22gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G1gat), .B(G8gat), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n316_), .B(new_n318_), .ZN(new_n319_));
  XOR2_X1   g118(.A(KEYINPUT77), .B(KEYINPUT78), .Z(new_n320_));
  NAND2_X1  g119(.A1(G231gat), .A2(G233gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n246_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n246_), .A2(new_n322_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n319_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n325_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n316_), .B(new_n317_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n327_), .A2(new_n328_), .A3(new_n323_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G127gat), .B(G155gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT16), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G183gat), .B(G211gat), .ZN(new_n332_));
  XOR2_X1   g131(.A(new_n331_), .B(new_n332_), .Z(new_n333_));
  NAND3_X1  g132(.A1(new_n326_), .A2(new_n329_), .A3(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT79), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n326_), .A2(new_n329_), .A3(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n333_), .ZN(new_n337_));
  AOI22_X1  g136(.A1(KEYINPUT17), .A2(new_n334_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n336_), .A2(KEYINPUT17), .A3(new_n337_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n311_), .B1(new_n338_), .B2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n336_), .A2(new_n337_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n334_), .A2(KEYINPUT17), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n344_), .A2(KEYINPUT80), .A3(new_n339_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n341_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n310_), .A2(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n273_), .A2(new_n348_), .ZN(new_n349_));
  XOR2_X1   g148(.A(new_n349_), .B(KEYINPUT81), .Z(new_n350_));
  INV_X1    g149(.A(KEYINPUT101), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT27), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G226gat), .A2(G233gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT19), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n356_));
  INV_X1    g155(.A(G169gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT23), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n360_), .B1(G183gat), .B2(G190gat), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT84), .ZN(new_n363_));
  INV_X1    g162(.A(G183gat), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n364_), .A2(KEYINPUT23), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n363_), .B1(new_n365_), .B2(G190gat), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n363_), .A2(new_n360_), .A3(G183gat), .A4(G190gat), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n362_), .B1(new_n366_), .B2(new_n368_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(G183gat), .A2(G190gat), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(KEYINPUT90), .B1(new_n369_), .B2(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n360_), .A2(G183gat), .A3(G190gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT84), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n361_), .B1(new_n374_), .B2(new_n367_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT90), .ZN(new_n376_));
  NOR3_X1   g175(.A1(new_n375_), .A2(new_n376_), .A3(new_n370_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n359_), .B1(new_n372_), .B2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n362_), .A2(new_n373_), .ZN(new_n379_));
  NOR3_X1   g178(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G169gat), .A2(G176gat), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n380_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n364_), .A2(KEYINPUT25), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT25), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(G183gat), .ZN(new_n387_));
  INV_X1    g186(.A(G190gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT26), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT26), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(G190gat), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n385_), .A2(new_n387_), .A3(new_n389_), .A4(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n379_), .A2(new_n384_), .A3(new_n392_), .ZN(new_n393_));
  XOR2_X1   g192(.A(G211gat), .B(G218gat), .Z(new_n394_));
  INV_X1    g193(.A(KEYINPUT88), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G197gat), .B(G204gat), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n394_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  AND2_X1   g196(.A1(new_n394_), .A2(new_n396_), .ZN(new_n398_));
  OAI21_X1  g197(.A(KEYINPUT21), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n396_), .A2(new_n395_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G211gat), .B(G218gat), .ZN(new_n401_));
  AOI21_X1  g200(.A(KEYINPUT21), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n399_), .A2(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n378_), .A2(new_n393_), .A3(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(KEYINPUT92), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT92), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n378_), .A2(new_n407_), .A3(new_n404_), .A4(new_n393_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n406_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT91), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n358_), .B1(new_n379_), .B2(new_n371_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT83), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n392_), .A2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT25), .B(G183gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(KEYINPUT26), .B(G190gat), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n414_), .A2(new_n415_), .A3(KEYINPUT83), .ZN(new_n416_));
  AND3_X1   g215(.A1(new_n413_), .A2(new_n384_), .A3(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n411_), .B1(new_n417_), .B2(new_n369_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n410_), .B1(new_n418_), .B2(new_n404_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n413_), .A2(new_n384_), .A3(new_n416_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n370_), .B1(new_n362_), .B2(new_n373_), .ZN(new_n421_));
  OAI22_X1  g220(.A1(new_n420_), .A2(new_n375_), .B1(new_n358_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n400_), .A2(new_n401_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n394_), .A2(new_n396_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n402_), .B1(new_n425_), .B2(KEYINPUT21), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n422_), .A2(new_n426_), .A3(KEYINPUT91), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n419_), .A2(KEYINPUT20), .A3(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n355_), .B1(new_n409_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT20), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n430_), .B1(new_n418_), .B2(new_n404_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n369_), .A2(KEYINPUT90), .A3(new_n371_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n376_), .B1(new_n375_), .B2(new_n370_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n358_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n393_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n426_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n431_), .A2(new_n436_), .A3(new_n354_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n429_), .A2(new_n437_), .ZN(new_n438_));
  XOR2_X1   g237(.A(G8gat), .B(G36gat), .Z(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(KEYINPUT94), .ZN(new_n440_));
  XOR2_X1   g239(.A(G64gat), .B(G92gat), .Z(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n443_));
  XOR2_X1   g242(.A(new_n442_), .B(new_n443_), .Z(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n352_), .B1(new_n438_), .B2(new_n445_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n419_), .A2(new_n405_), .A3(KEYINPUT20), .A4(new_n427_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(new_n354_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT98), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n431_), .A2(new_n436_), .A3(new_n449_), .A4(new_n355_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n431_), .A2(new_n436_), .A3(new_n355_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT98), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n448_), .A2(new_n450_), .A3(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n444_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT99), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT99), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n453_), .A2(new_n456_), .A3(new_n444_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n446_), .A2(new_n455_), .A3(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT100), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n437_), .ZN(new_n461_));
  AND2_X1   g260(.A1(new_n427_), .A2(KEYINPUT20), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n462_), .A2(new_n406_), .A3(new_n419_), .A4(new_n408_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n461_), .B1(new_n463_), .B2(new_n355_), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT27), .B1(new_n464_), .B2(new_n444_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n456_), .B1(new_n453_), .B2(new_n444_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n467_), .A2(KEYINPUT100), .A3(new_n457_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n438_), .A2(new_n445_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n464_), .A2(new_n444_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  AOI22_X1  g270(.A1(new_n460_), .A2(new_n468_), .B1(new_n352_), .B2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G78gat), .B(G106gat), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT3), .ZN(new_n474_));
  INV_X1    g273(.A(G141gat), .ZN(new_n475_));
  INV_X1    g274(.A(G148gat), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n474_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G141gat), .A2(G148gat), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT2), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n481_));
  OAI21_X1  g280(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n477_), .A2(new_n480_), .A3(new_n481_), .A4(new_n482_), .ZN(new_n483_));
  XOR2_X1   g282(.A(G155gat), .B(G162gat), .Z(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT87), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n485_), .B(new_n486_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(G155gat), .A2(G162gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G155gat), .A2(G162gat), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n488_), .B1(KEYINPUT1), .B2(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n490_), .B1(KEYINPUT1), .B2(new_n489_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n475_), .A2(new_n476_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n491_), .A2(new_n478_), .A3(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n487_), .A2(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n404_), .B1(new_n494_), .B2(KEYINPUT29), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G228gat), .A2(G233gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n495_), .A2(new_n496_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n473_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT89), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  OR2_X1    g301(.A1(new_n494_), .A2(KEYINPUT29), .ZN(new_n503_));
  XOR2_X1   g302(.A(G22gat), .B(G50gat), .Z(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(KEYINPUT28), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n503_), .B(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n499_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n473_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n507_), .A2(new_n497_), .A3(new_n508_), .ZN(new_n509_));
  AOI22_X1  g308(.A1(new_n502_), .A2(new_n506_), .B1(new_n500_), .B2(new_n509_), .ZN(new_n510_));
  AND4_X1   g309(.A1(KEYINPUT89), .A2(new_n500_), .A3(new_n509_), .A4(new_n506_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G71gat), .B(G99gat), .ZN(new_n514_));
  INV_X1    g313(.A(G43gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT30), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(new_n418_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G227gat), .A2(G233gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(G15gat), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n518_), .A2(new_n520_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n521_), .A2(KEYINPUT86), .A3(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G127gat), .B(G134gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT85), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G113gat), .B(G120gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  XOR2_X1   g326(.A(new_n527_), .B(KEYINPUT31), .Z(new_n528_));
  OR2_X1    g327(.A1(new_n523_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n523_), .A2(new_n528_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n527_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(new_n494_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n527_), .A2(new_n487_), .A3(new_n493_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(KEYINPUT4), .A3(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT4), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n533_), .A2(new_n494_), .A3(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G225gat), .A2(G233gat), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G57gat), .B(G85gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  XOR2_X1   g344(.A(G1gat), .B(G29gat), .Z(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT96), .B(KEYINPUT97), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n534_), .A2(new_n535_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n542_), .B(new_n550_), .C1(new_n541_), .C2(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n552_), .A2(new_n541_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n540_), .B1(new_n536_), .B2(new_n538_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n549_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n553_), .A2(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n532_), .A2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n472_), .A2(new_n513_), .A3(new_n558_), .ZN(new_n559_));
  AND2_X1   g358(.A1(new_n445_), .A2(KEYINPUT32), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(new_n453_), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n557_), .B(new_n561_), .C1(new_n560_), .C2(new_n464_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n550_), .B1(new_n551_), .B2(new_n540_), .ZN(new_n563_));
  AND3_X1   g362(.A1(new_n536_), .A2(new_n540_), .A3(new_n538_), .ZN(new_n564_));
  OAI21_X1  g363(.A(KEYINPUT33), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(new_n556_), .ZN(new_n566_));
  OAI211_X1 g365(.A(KEYINPUT33), .B(new_n549_), .C1(new_n554_), .C2(new_n555_), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n566_), .A2(new_n469_), .A3(new_n470_), .A4(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n512_), .B1(new_n562_), .B2(new_n568_), .ZN(new_n569_));
  NOR3_X1   g368(.A1(new_n510_), .A2(new_n557_), .A3(new_n511_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n569_), .B1(new_n472_), .B2(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n559_), .B1(new_n571_), .B2(new_n531_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n277_), .A2(new_n328_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n319_), .A2(new_n276_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G229gat), .A2(G233gat), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n573_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n328_), .A2(new_n286_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n574_), .A2(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n576_), .B1(new_n578_), .B2(new_n575_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G113gat), .B(G141gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G169gat), .B(G197gat), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n580_), .B(new_n581_), .Z(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n579_), .A2(new_n583_), .ZN(new_n584_));
  OAI211_X1 g383(.A(new_n576_), .B(new_n582_), .C1(new_n578_), .C2(new_n575_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n584_), .A2(KEYINPUT82), .A3(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT82), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n579_), .A2(new_n587_), .A3(new_n583_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n586_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n572_), .A2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n350_), .A2(new_n351_), .A3(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n349_), .B(KEYINPUT81), .ZN(new_n593_));
  INV_X1    g392(.A(new_n591_), .ZN(new_n594_));
  OAI21_X1  g393(.A(KEYINPUT101), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n592_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n557_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n597_), .A2(new_n312_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n596_), .A2(KEYINPUT38), .A3(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n303_), .A2(new_n306_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n572_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n344_), .A2(new_n339_), .ZN(new_n602_));
  AND4_X1   g401(.A1(new_n590_), .A2(new_n270_), .A3(new_n272_), .A4(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n601_), .A2(KEYINPUT102), .A3(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n603_), .A2(new_n572_), .A3(new_n600_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT102), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n604_), .A2(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(G1gat), .B1(new_n608_), .B2(new_n597_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n592_), .A2(new_n595_), .A3(new_n598_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT38), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n599_), .A2(new_n609_), .A3(new_n612_), .ZN(G1324gat));
  NOR2_X1   g412(.A1(new_n472_), .A2(G8gat), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n592_), .A2(new_n595_), .A3(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(G8gat), .B1(new_n605_), .B2(new_n472_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT39), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT40), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(G1325gat));
  INV_X1    g419(.A(KEYINPUT41), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n532_), .B1(new_n604_), .B2(new_n607_), .ZN(new_n622_));
  INV_X1    g421(.A(G15gat), .ZN(new_n623_));
  OAI21_X1  g422(.A(KEYINPUT103), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NOR3_X1   g424(.A1(new_n622_), .A2(KEYINPUT103), .A3(new_n623_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n621_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n626_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n628_), .A2(new_n624_), .A3(KEYINPUT41), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n596_), .A2(new_n623_), .A3(new_n531_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n627_), .A2(new_n629_), .A3(new_n630_), .ZN(G1326gat));
  OAI21_X1  g430(.A(G22gat), .B1(new_n608_), .B2(new_n513_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT42), .ZN(new_n633_));
  INV_X1    g432(.A(G22gat), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n596_), .A2(new_n634_), .A3(new_n512_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(G1327gat));
  INV_X1    g435(.A(new_n273_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n600_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(new_n346_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n591_), .A2(new_n637_), .A3(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(G29gat), .B1(new_n642_), .B2(new_n557_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n310_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n471_), .A2(new_n352_), .ZN(new_n645_));
  AOI21_X1  g444(.A(KEYINPUT100), .B1(new_n467_), .B2(new_n457_), .ZN(new_n646_));
  AND4_X1   g445(.A1(KEYINPUT100), .A2(new_n446_), .A3(new_n455_), .A4(new_n457_), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n570_), .B(new_n645_), .C1(new_n646_), .C2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n562_), .A2(new_n568_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(new_n513_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n531_), .B1(new_n648_), .B2(new_n650_), .ZN(new_n651_));
  OAI211_X1 g450(.A(new_n513_), .B(new_n645_), .C1(new_n646_), .C2(new_n647_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n558_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n644_), .B1(new_n651_), .B2(new_n654_), .ZN(new_n655_));
  OAI21_X1  g454(.A(KEYINPUT104), .B1(new_n307_), .B2(new_n309_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(KEYINPUT43), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n655_), .A2(new_n658_), .ZN(new_n659_));
  OAI211_X1 g458(.A(new_n644_), .B(new_n657_), .C1(new_n651_), .C2(new_n654_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n273_), .A2(new_n347_), .A3(new_n589_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n661_), .A2(KEYINPUT44), .A3(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(KEYINPUT44), .B1(new_n661_), .B2(new_n662_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n557_), .A2(G29gat), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n643_), .B1(new_n666_), .B2(new_n667_), .ZN(G1328gat));
  INV_X1    g467(.A(new_n472_), .ZN(new_n669_));
  INV_X1    g468(.A(G36gat), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  OR3_X1    g470(.A1(new_n641_), .A2(KEYINPUT45), .A3(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(KEYINPUT45), .B1(new_n641_), .B2(new_n671_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n664_), .A2(new_n665_), .A3(new_n472_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n674_), .B1(new_n675_), .B2(new_n670_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT46), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  OAI211_X1 g477(.A(new_n674_), .B(KEYINPUT46), .C1(new_n675_), .C2(new_n670_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(G1329gat));
  AOI21_X1  g479(.A(new_n657_), .B1(new_n572_), .B2(new_n644_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n660_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n662_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n532_), .A2(new_n515_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n685_), .A2(new_n663_), .A3(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT105), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n685_), .A2(KEYINPUT105), .A3(new_n663_), .A4(new_n686_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n515_), .B1(new_n641_), .B2(new_n532_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n689_), .A2(new_n690_), .A3(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(KEYINPUT47), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT47), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n689_), .A2(new_n694_), .A3(new_n690_), .A4(new_n691_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n693_), .A2(new_n695_), .ZN(G1330gat));
  AOI21_X1  g495(.A(G50gat), .B1(new_n642_), .B2(new_n512_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n512_), .A2(G50gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n697_), .B1(new_n666_), .B2(new_n698_), .ZN(G1331gat));
  AND2_X1   g498(.A1(new_n572_), .A2(new_n589_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n637_), .A2(new_n348_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(G57gat), .B1(new_n703_), .B2(new_n557_), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n341_), .A2(new_n345_), .A3(new_n589_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n273_), .A2(new_n705_), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n601_), .A2(G57gat), .A3(new_n557_), .A4(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT106), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n707_), .A2(new_n708_), .ZN(new_n710_));
  NOR3_X1   g509(.A1(new_n704_), .A2(new_n709_), .A3(new_n710_), .ZN(G1332gat));
  NAND2_X1  g510(.A1(new_n601_), .A2(new_n706_), .ZN(new_n712_));
  OAI21_X1  g511(.A(G64gat), .B1(new_n712_), .B2(new_n472_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT48), .ZN(new_n714_));
  OR2_X1    g513(.A1(new_n472_), .A2(G64gat), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n714_), .B1(new_n702_), .B2(new_n715_), .ZN(G1333gat));
  OAI21_X1  g515(.A(G71gat), .B1(new_n712_), .B2(new_n532_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT49), .ZN(new_n718_));
  OR2_X1    g517(.A1(new_n532_), .A2(G71gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n718_), .B1(new_n702_), .B2(new_n719_), .ZN(G1334gat));
  OAI21_X1  g519(.A(G78gat), .B1(new_n712_), .B2(new_n513_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT50), .ZN(new_n722_));
  OR2_X1    g521(.A1(new_n513_), .A2(G78gat), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n722_), .B1(new_n702_), .B2(new_n723_), .ZN(G1335gat));
  INV_X1    g523(.A(KEYINPUT107), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n700_), .A2(new_n725_), .A3(new_n273_), .A4(new_n640_), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n572_), .A2(new_n640_), .A3(new_n589_), .A4(new_n273_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(KEYINPUT107), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(G85gat), .B1(new_n729_), .B2(new_n557_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n661_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n273_), .A2(new_n589_), .A3(new_n346_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n557_), .A2(G85gat), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n733_), .B(KEYINPUT108), .Z(new_n734_));
  NOR3_X1   g533(.A1(new_n731_), .A2(new_n732_), .A3(new_n734_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n730_), .A2(new_n735_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT109), .ZN(G1336gat));
  NAND3_X1  g536(.A1(new_n729_), .A2(new_n212_), .A3(new_n669_), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n731_), .A2(new_n472_), .A3(new_n732_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n738_), .B1(new_n739_), .B2(new_n212_), .ZN(G1337gat));
  NAND2_X1  g539(.A1(new_n531_), .A2(new_n207_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n741_), .B1(new_n726_), .B2(new_n728_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n732_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n661_), .A2(new_n531_), .A3(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(G99gat), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(KEYINPUT110), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT110), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n744_), .A2(new_n747_), .A3(G99gat), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n742_), .B1(new_n746_), .B2(new_n748_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(KEYINPUT111), .B(KEYINPUT51), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n750_), .ZN(new_n752_));
  AOI211_X1 g551(.A(new_n742_), .B(new_n752_), .C1(new_n746_), .C2(new_n748_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n751_), .A2(new_n753_), .ZN(G1338gat));
  INV_X1    g553(.A(KEYINPUT112), .ZN(new_n755_));
  AOI211_X1 g554(.A(new_n513_), .B(new_n732_), .C1(new_n659_), .C2(new_n660_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n755_), .B1(new_n756_), .B2(new_n208_), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n512_), .B(new_n743_), .C1(new_n681_), .C2(new_n682_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n758_), .A2(KEYINPUT112), .A3(G106gat), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n757_), .A2(KEYINPUT52), .A3(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n512_), .A2(new_n208_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n761_), .B1(new_n726_), .B2(new_n728_), .ZN(new_n762_));
  AOI21_X1  g561(.A(KEYINPUT112), .B1(new_n758_), .B2(G106gat), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT52), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n762_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n760_), .A2(new_n765_), .A3(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n760_), .B2(new_n765_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n767_), .A2(new_n768_), .ZN(G1339gat));
  XNOR2_X1  g568(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n269_), .A2(new_n705_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n771_), .B2(new_n310_), .ZN(new_n772_));
  AND4_X1   g571(.A1(new_n269_), .A2(new_n310_), .A3(new_n705_), .A4(new_n770_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT58), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n250_), .A2(new_n257_), .A3(new_n252_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n255_), .A2(KEYINPUT55), .A3(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n257_), .B1(new_n250_), .B2(new_n252_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT55), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n265_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n777_), .A2(KEYINPUT56), .A3(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT56), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n250_), .A2(new_n257_), .A3(new_n252_), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n784_), .A2(new_n778_), .A3(new_n779_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n253_), .A2(new_n779_), .A3(new_n254_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(new_n263_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n783_), .B1(new_n785_), .B2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT118), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n777_), .A2(new_n780_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT118), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n790_), .A2(new_n791_), .A3(new_n783_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n782_), .B1(new_n789_), .B2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n575_), .ZN(new_n794_));
  OAI211_X1 g593(.A(KEYINPUT116), .B(new_n583_), .C1(new_n578_), .C2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT116), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n794_), .B1(new_n577_), .B2(new_n574_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n796_), .B1(new_n797_), .B2(new_n582_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n573_), .A2(new_n574_), .A3(new_n794_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n795_), .A2(new_n798_), .A3(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT117), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n800_), .A2(new_n801_), .A3(new_n585_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n801_), .B1(new_n800_), .B2(new_n585_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(new_n266_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n775_), .B1(new_n793_), .B2(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n791_), .B1(new_n790_), .B2(new_n783_), .ZN(new_n808_));
  AOI211_X1 g607(.A(KEYINPUT118), .B(KEYINPUT56), .C1(new_n777_), .C2(new_n780_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n781_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n810_), .A2(KEYINPUT58), .A3(new_n266_), .A4(new_n805_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n807_), .A2(new_n811_), .A3(new_n644_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT57), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n804_), .B1(new_n264_), .B2(new_n266_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n590_), .A2(new_n266_), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT115), .B1(new_n790_), .B2(new_n783_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n815_), .B1(new_n816_), .B2(new_n781_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n777_), .A2(new_n780_), .A3(KEYINPUT115), .A4(KEYINPUT56), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n814_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n813_), .B1(new_n819_), .B2(new_n638_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT115), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n788_), .A2(new_n821_), .A3(new_n781_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n822_), .A2(new_n590_), .A3(new_n266_), .A4(new_n818_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n814_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n825_), .A2(KEYINPUT57), .A3(new_n600_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n812_), .A2(new_n820_), .A3(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n602_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n774_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n472_), .A2(new_n557_), .A3(new_n513_), .A4(new_n531_), .ZN(new_n830_));
  OR3_X1    g629(.A1(new_n829_), .A2(KEYINPUT119), .A3(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(G113gat), .ZN(new_n832_));
  OAI21_X1  g631(.A(KEYINPUT119), .B1(new_n829_), .B2(new_n830_), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n831_), .A2(new_n832_), .A3(new_n590_), .A4(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n774_), .B1(new_n827_), .B2(new_n346_), .ZN(new_n835_));
  NOR3_X1   g634(.A1(new_n835_), .A2(KEYINPUT59), .A3(new_n830_), .ZN(new_n836_));
  OAI21_X1  g635(.A(KEYINPUT59), .B1(new_n829_), .B2(new_n830_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(KEYINPUT120), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT120), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n839_), .B(KEYINPUT59), .C1(new_n829_), .C2(new_n830_), .ZN(new_n840_));
  AOI211_X1 g639(.A(new_n589_), .B(new_n836_), .C1(new_n838_), .C2(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n834_), .B1(new_n841_), .B2(new_n832_), .ZN(G1340gat));
  INV_X1    g641(.A(G120gat), .ZN(new_n843_));
  OR2_X1    g642(.A1(new_n843_), .A2(KEYINPUT60), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n843_), .B1(new_n637_), .B2(KEYINPUT60), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n831_), .A2(new_n833_), .A3(new_n844_), .A4(new_n845_), .ZN(new_n846_));
  AOI211_X1 g645(.A(new_n637_), .B(new_n836_), .C1(new_n838_), .C2(new_n840_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n846_), .B1(new_n847_), .B2(new_n843_), .ZN(G1341gat));
  INV_X1    g647(.A(G127gat), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n831_), .A2(new_n849_), .A3(new_n347_), .A4(new_n833_), .ZN(new_n850_));
  AOI211_X1 g649(.A(new_n828_), .B(new_n836_), .C1(new_n838_), .C2(new_n840_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n850_), .B1(new_n851_), .B2(new_n849_), .ZN(G1342gat));
  INV_X1    g651(.A(G134gat), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n831_), .A2(new_n853_), .A3(new_n638_), .A4(new_n833_), .ZN(new_n854_));
  AOI211_X1 g653(.A(new_n310_), .B(new_n836_), .C1(new_n838_), .C2(new_n840_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n855_), .B2(new_n853_), .ZN(G1343gat));
  NOR2_X1   g655(.A1(new_n829_), .A2(new_n531_), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n669_), .A2(new_n597_), .A3(new_n513_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n859_), .A2(new_n589_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(new_n475_), .ZN(G1344gat));
  NOR2_X1   g660(.A1(new_n859_), .A2(new_n637_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(new_n476_), .ZN(G1345gat));
  INV_X1    g662(.A(new_n829_), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n864_), .A2(new_n532_), .A3(new_n347_), .A4(new_n858_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(KEYINPUT121), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT121), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n857_), .A2(new_n867_), .A3(new_n347_), .A4(new_n858_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(KEYINPUT61), .B(G155gat), .ZN(new_n869_));
  AND3_X1   g668(.A1(new_n866_), .A2(new_n868_), .A3(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n869_), .B1(new_n866_), .B2(new_n868_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n870_), .A2(new_n871_), .ZN(G1346gat));
  OAI21_X1  g671(.A(G162gat), .B1(new_n859_), .B2(new_n310_), .ZN(new_n873_));
  OR2_X1    g672(.A1(new_n600_), .A2(G162gat), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n873_), .B1(new_n859_), .B2(new_n874_), .ZN(G1347gat));
  NOR2_X1   g674(.A1(new_n472_), .A2(new_n653_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n513_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n835_), .A2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n590_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT62), .ZN(new_n880_));
  AND4_X1   g679(.A1(KEYINPUT122), .A2(new_n879_), .A3(new_n880_), .A4(G169gat), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT122), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n357_), .B1(new_n882_), .B2(KEYINPUT62), .ZN(new_n883_));
  AOI22_X1  g682(.A1(new_n879_), .A2(new_n883_), .B1(KEYINPUT122), .B2(new_n880_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n878_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(KEYINPUT22), .B(G169gat), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n590_), .A2(new_n886_), .ZN(new_n887_));
  XOR2_X1   g686(.A(new_n887_), .B(KEYINPUT123), .Z(new_n888_));
  OAI22_X1  g687(.A1(new_n881_), .A2(new_n884_), .B1(new_n885_), .B2(new_n888_), .ZN(G1348gat));
  AOI21_X1  g688(.A(G176gat), .B1(new_n878_), .B2(new_n273_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n829_), .A2(new_n512_), .ZN(new_n891_));
  AND3_X1   g690(.A1(new_n273_), .A2(G176gat), .A3(new_n876_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n890_), .B1(new_n891_), .B2(new_n892_), .ZN(G1349gat));
  NAND3_X1  g692(.A1(new_n891_), .A2(new_n347_), .A3(new_n876_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n828_), .A2(new_n414_), .ZN(new_n895_));
  AOI22_X1  g694(.A1(new_n894_), .A2(new_n364_), .B1(new_n878_), .B2(new_n895_), .ZN(G1350gat));
  OAI21_X1  g695(.A(G190gat), .B1(new_n885_), .B2(new_n310_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n638_), .A2(new_n415_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(KEYINPUT124), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n897_), .B1(new_n885_), .B2(new_n899_), .ZN(G1351gat));
  NAND2_X1  g699(.A1(new_n669_), .A2(new_n570_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n857_), .A2(new_n590_), .A3(new_n902_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g703(.A1(new_n857_), .A2(new_n273_), .A3(new_n902_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(G204gat), .ZN(G1353gat));
  XNOR2_X1  g705(.A(KEYINPUT63), .B(G211gat), .ZN(new_n907_));
  NAND4_X1  g706(.A1(new_n857_), .A2(new_n602_), .A3(new_n902_), .A4(new_n907_), .ZN(new_n908_));
  NOR4_X1   g707(.A1(new_n829_), .A2(new_n531_), .A3(new_n828_), .A4(new_n901_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n908_), .B1(new_n909_), .B2(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(KEYINPUT125), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT125), .ZN(new_n913_));
  OAI211_X1 g712(.A(new_n908_), .B(new_n913_), .C1(new_n909_), .C2(new_n910_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n912_), .A2(new_n914_), .ZN(G1354gat));
  NAND2_X1  g714(.A1(new_n857_), .A2(new_n902_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n644_), .A2(G218gat), .ZN(new_n917_));
  XOR2_X1   g716(.A(new_n917_), .B(KEYINPUT127), .Z(new_n918_));
  NOR2_X1   g717(.A1(new_n916_), .A2(new_n918_), .ZN(new_n919_));
  OAI21_X1  g718(.A(KEYINPUT126), .B1(new_n916_), .B2(new_n600_), .ZN(new_n920_));
  NOR4_X1   g719(.A1(new_n829_), .A2(new_n531_), .A3(new_n600_), .A4(new_n901_), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT126), .ZN(new_n922_));
  AOI21_X1  g721(.A(G218gat), .B1(new_n921_), .B2(new_n922_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n919_), .B1(new_n920_), .B2(new_n923_), .ZN(G1355gat));
endmodule


