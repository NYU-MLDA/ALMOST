//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 0 1 1 1 0 1 1 1 0 0 1 0 1 0 0 1 1 1 0 0 1 1 1 0 1 0 1 1 0 0 0 1 1 1 1 1 1 1 1 0 0 1 1 0 1 0 1 1 1 1 1 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n596_, new_n597_, new_n598_, new_n599_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n677_, new_n678_, new_n679_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n688_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n804_, new_n805_, new_n806_, new_n808_,
    new_n809_, new_n810_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n817_, new_n819_, new_n820_, new_n822_, new_n823_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n837_, new_n838_,
    new_n840_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n864_, new_n865_, new_n866_;
  XOR2_X1   g000(.A(G190gat), .B(G218gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G134gat), .B(G162gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT36), .ZN(new_n205_));
  AND2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  XOR2_X1   g005(.A(G29gat), .B(G36gat), .Z(new_n207_));
  XNOR2_X1  g006(.A(G43gat), .B(G50gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  XOR2_X1   g008(.A(new_n209_), .B(KEYINPUT15), .Z(new_n210_));
  AND3_X1   g009(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n211_));
  AOI21_X1  g010(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G99gat), .ZN(new_n214_));
  INV_X1    g013(.A(G106gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n214_), .A2(new_n215_), .A3(KEYINPUT65), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT7), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT7), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n218_), .A2(new_n214_), .A3(new_n215_), .A4(KEYINPUT65), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n213_), .A2(new_n217_), .A3(new_n219_), .ZN(new_n220_));
  AND2_X1   g019(.A1(G85gat), .A2(G92gat), .ZN(new_n221_));
  NOR2_X1   g020(.A1(G85gat), .A2(G92gat), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n220_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n220_), .A2(KEYINPUT66), .A3(KEYINPUT8), .A4(new_n223_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT9), .ZN(new_n228_));
  INV_X1    g027(.A(G85gat), .ZN(new_n229_));
  INV_X1    g028(.A(G92gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G85gat), .A2(G92gat), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n228_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n228_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT64), .B1(new_n233_), .B2(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(KEYINPUT10), .B(G99gat), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n237_), .A2(G106gat), .ZN(new_n238_));
  OAI21_X1  g037(.A(KEYINPUT9), .B1(new_n221_), .B2(new_n222_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT64), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(new_n240_), .A3(new_n234_), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n236_), .A2(new_n213_), .A3(new_n238_), .A4(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n226_), .A2(new_n227_), .A3(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n210_), .A2(new_n243_), .ZN(new_n244_));
  XOR2_X1   g043(.A(KEYINPUT68), .B(KEYINPUT34), .Z(new_n245_));
  NAND2_X1  g044(.A1(G232gat), .A2(G233gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  OAI221_X1 g046(.A(new_n244_), .B1(KEYINPUT35), .B2(new_n247_), .C1(new_n209_), .C2(new_n243_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(KEYINPUT35), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n249_), .B1(new_n244_), .B2(KEYINPUT69), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n248_), .B(new_n250_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n204_), .A2(new_n205_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n206_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT70), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n251_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n251_), .B(new_n254_), .C1(new_n206_), .C2(new_n252_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT37), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G15gat), .B(G22gat), .ZN(new_n260_));
  INV_X1    g059(.A(G1gat), .ZN(new_n261_));
  INV_X1    g060(.A(G8gat), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT14), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n260_), .A2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G1gat), .B(G8gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n264_), .B(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G231gat), .A2(G233gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G57gat), .B(G64gat), .ZN(new_n269_));
  OR2_X1    g068(.A1(new_n269_), .A2(KEYINPUT11), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(KEYINPUT11), .ZN(new_n271_));
  XOR2_X1   g070(.A(G71gat), .B(G78gat), .Z(new_n272_));
  NAND3_X1  g071(.A1(new_n270_), .A2(new_n271_), .A3(new_n272_), .ZN(new_n273_));
  OR2_X1    g072(.A1(new_n271_), .A2(new_n272_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n268_), .B(new_n276_), .ZN(new_n277_));
  XOR2_X1   g076(.A(G127gat), .B(G155gat), .Z(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT16), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G183gat), .B(G211gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT17), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  AND2_X1   g082(.A1(new_n281_), .A2(new_n282_), .ZN(new_n284_));
  OR3_X1    g083(.A1(new_n277_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n277_), .A2(new_n283_), .ZN(new_n286_));
  AND2_X1   g085(.A1(new_n286_), .A2(KEYINPUT71), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n286_), .A2(KEYINPUT71), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n285_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  OR2_X1    g088(.A1(new_n289_), .A2(KEYINPUT72), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(KEYINPUT72), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  AND4_X1   g091(.A1(new_n275_), .A2(new_n226_), .A3(new_n227_), .A4(new_n242_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT12), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n294_), .A2(KEYINPUT67), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n295_), .B1(new_n243_), .B2(new_n276_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(KEYINPUT67), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n293_), .B1(new_n296_), .B2(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n240_), .B1(new_n239_), .B2(new_n234_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n213_), .B1(G106gat), .B2(new_n237_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  AOI22_X1  g101(.A1(new_n302_), .A2(new_n241_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n275_), .B1(new_n303_), .B2(new_n227_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n297_), .B1(new_n304_), .B2(new_n295_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G230gat), .A2(G233gat), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n299_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n306_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n308_), .B1(new_n304_), .B2(new_n293_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G120gat), .B(G148gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT5), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G176gat), .B(G204gat), .ZN(new_n313_));
  XOR2_X1   g112(.A(new_n312_), .B(new_n313_), .Z(new_n314_));
  NAND2_X1  g113(.A1(new_n310_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n314_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n307_), .A2(new_n309_), .A3(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  OR2_X1    g117(.A1(new_n318_), .A2(KEYINPUT13), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(KEYINPUT13), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NOR3_X1   g121(.A1(new_n259_), .A2(new_n292_), .A3(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT73), .ZN(new_n324_));
  AND2_X1   g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n323_), .A2(new_n324_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n210_), .A2(new_n266_), .ZN(new_n327_));
  OR2_X1    g126(.A1(new_n266_), .A2(new_n209_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G229gat), .A2(G233gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT74), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n328_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n266_), .A2(new_n209_), .ZN(new_n334_));
  MUX2_X1   g133(.A(new_n332_), .B(new_n333_), .S(new_n334_), .Z(new_n335_));
  OAI21_X1  g134(.A(new_n331_), .B1(new_n335_), .B2(new_n330_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G113gat), .B(G141gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G169gat), .B(G197gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n336_), .B(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G141gat), .A2(G148gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT2), .ZN(new_n342_));
  NOR2_X1   g141(.A1(G141gat), .A2(G148gat), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT3), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT3), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n343_), .A2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n342_), .A2(new_n345_), .A3(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT79), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G155gat), .A2(G162gat), .ZN(new_n351_));
  NOR2_X1   g150(.A1(G155gat), .A2(G162gat), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n350_), .A2(new_n351_), .A3(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT29), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n352_), .B1(KEYINPUT1), .B2(new_n351_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n356_), .B1(KEYINPUT1), .B2(new_n351_), .ZN(new_n357_));
  AND3_X1   g156(.A1(new_n357_), .A2(new_n341_), .A3(new_n344_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n354_), .A2(new_n355_), .A3(new_n359_), .ZN(new_n360_));
  XOR2_X1   g159(.A(G22gat), .B(G50gat), .Z(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G78gat), .B(G106gat), .ZN(new_n364_));
  AND3_X1   g163(.A1(new_n350_), .A2(new_n351_), .A3(new_n353_), .ZN(new_n365_));
  OAI21_X1  g164(.A(KEYINPUT29), .B1(new_n365_), .B2(new_n358_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G211gat), .B(G218gat), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n367_), .A2(KEYINPUT21), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G197gat), .B(G204gat), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n367_), .A2(KEYINPUT21), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(KEYINPUT81), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n373_), .A2(G228gat), .A3(G233gat), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n366_), .A2(new_n372_), .A3(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n374_), .B1(new_n366_), .B2(new_n372_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n364_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n377_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n364_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n379_), .A2(new_n375_), .A3(new_n380_), .ZN(new_n381_));
  XOR2_X1   g180(.A(KEYINPUT80), .B(KEYINPUT28), .Z(new_n382_));
  AND3_X1   g181(.A1(new_n378_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n382_), .B1(new_n378_), .B2(new_n381_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n363_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n378_), .A2(new_n381_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n382_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n378_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n388_), .A2(new_n362_), .A3(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n385_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT27), .ZN(new_n392_));
  XOR2_X1   g191(.A(KEYINPUT82), .B(KEYINPUT19), .Z(new_n393_));
  NAND2_X1  g192(.A1(G226gat), .A2(G233gat), .ZN(new_n394_));
  XOR2_X1   g193(.A(new_n393_), .B(new_n394_), .Z(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(KEYINPUT83), .ZN(new_n396_));
  INV_X1    g195(.A(G183gat), .ZN(new_n397_));
  INV_X1    g196(.A(G190gat), .ZN(new_n398_));
  OAI21_X1  g197(.A(KEYINPUT23), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT23), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n400_), .A2(G183gat), .A3(G190gat), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n399_), .A2(KEYINPUT77), .A3(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT77), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n403_), .A2(new_n400_), .A3(G183gat), .A4(G190gat), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n405_), .B1(G183gat), .B2(G190gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G169gat), .A2(G176gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(KEYINPUT22), .B(G169gat), .ZN(new_n408_));
  INV_X1    g207(.A(G176gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n406_), .A2(new_n407_), .A3(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(KEYINPUT26), .B(G190gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT76), .ZN(new_n413_));
  OR3_X1    g212(.A1(new_n398_), .A2(KEYINPUT76), .A3(KEYINPUT26), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT25), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT75), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n415_), .B1(new_n416_), .B2(new_n397_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(KEYINPUT75), .A2(KEYINPUT25), .A3(G183gat), .ZN(new_n418_));
  AOI22_X1  g217(.A1(new_n413_), .A2(new_n414_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  OR2_X1    g218(.A1(G169gat), .A2(G176gat), .ZN(new_n420_));
  OR2_X1    g219(.A1(new_n420_), .A2(KEYINPUT24), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n399_), .A2(new_n401_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n420_), .A2(KEYINPUT24), .A3(new_n407_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n421_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  OR2_X1    g223(.A1(new_n419_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n411_), .A2(new_n425_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n426_), .A2(new_n372_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT20), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n422_), .B1(G183gat), .B2(G190gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n407_), .B(KEYINPUT85), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n430_), .A2(new_n410_), .A3(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n405_), .A2(KEYINPUT84), .A3(new_n421_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(KEYINPUT25), .B(G183gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n412_), .A2(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n433_), .A2(new_n423_), .A3(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(KEYINPUT84), .B1(new_n405_), .B2(new_n421_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n432_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(new_n372_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n396_), .B1(new_n429_), .B2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n426_), .A2(new_n372_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT86), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT86), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n426_), .A2(new_n443_), .A3(new_n372_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n395_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT20), .B1(new_n438_), .B2(new_n372_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT87), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT87), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n445_), .A2(new_n447_), .A3(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n440_), .B1(new_n449_), .B2(new_n451_), .ZN(new_n452_));
  XOR2_X1   g251(.A(G8gat), .B(G36gat), .Z(new_n453_));
  XNOR2_X1  g252(.A(G64gat), .B(G92gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(KEYINPUT88), .B(KEYINPUT18), .ZN(new_n456_));
  XOR2_X1   g255(.A(new_n455_), .B(new_n456_), .Z(new_n457_));
  NOR2_X1   g256(.A1(new_n452_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n457_), .ZN(new_n459_));
  AOI211_X1 g258(.A(new_n459_), .B(new_n440_), .C1(new_n449_), .C2(new_n451_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n392_), .B1(new_n458_), .B2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n429_), .A2(new_n439_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n396_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n442_), .A2(new_n444_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT93), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n446_), .A2(new_n466_), .ZN(new_n467_));
  OAI211_X1 g266(.A(KEYINPUT93), .B(KEYINPUT20), .C1(new_n438_), .C2(new_n372_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n465_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n464_), .B1(new_n469_), .B2(new_n395_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(new_n459_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n452_), .A2(new_n457_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n472_), .A2(new_n473_), .A3(KEYINPUT27), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n391_), .A2(new_n461_), .A3(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n426_), .B(KEYINPUT30), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G71gat), .B(G99gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(G43gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G227gat), .A2(G233gat), .ZN(new_n479_));
  INV_X1    g278(.A(G15gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n478_), .B(new_n481_), .ZN(new_n482_));
  XOR2_X1   g281(.A(new_n476_), .B(new_n482_), .Z(new_n483_));
  INV_X1    g282(.A(KEYINPUT31), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n476_), .B(new_n482_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT31), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n485_), .A2(new_n487_), .ZN(new_n488_));
  XOR2_X1   g287(.A(G127gat), .B(G134gat), .Z(new_n489_));
  XOR2_X1   g288(.A(G113gat), .B(G120gat), .Z(new_n490_));
  OR2_X1    g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  OR2_X1    g290(.A1(new_n491_), .A2(KEYINPUT78), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(KEYINPUT78), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n489_), .A2(new_n490_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n492_), .A2(new_n493_), .A3(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n488_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n495_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n485_), .A2(new_n497_), .A3(new_n487_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n497_), .B1(new_n365_), .B2(new_n358_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n491_), .A2(new_n494_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n354_), .A2(new_n359_), .A3(new_n501_), .ZN(new_n502_));
  AND2_X1   g301(.A1(new_n500_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G225gat), .A2(G233gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(KEYINPUT89), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n503_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT4), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n508_), .B(new_n497_), .C1(new_n365_), .C2(new_n358_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT90), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n500_), .A2(KEYINPUT4), .A3(new_n502_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(new_n505_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n507_), .B1(new_n511_), .B2(new_n513_), .ZN(new_n514_));
  XOR2_X1   g313(.A(G1gat), .B(G29gat), .Z(new_n515_));
  XNOR2_X1  g314(.A(G57gat), .B(G85gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(KEYINPUT91), .B(KEYINPUT0), .ZN(new_n518_));
  XOR2_X1   g317(.A(new_n517_), .B(new_n518_), .Z(new_n519_));
  NAND2_X1  g318(.A1(new_n514_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n519_), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n507_), .B(new_n521_), .C1(new_n511_), .C2(new_n513_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT96), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT96), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n520_), .A2(new_n525_), .A3(new_n522_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n499_), .A2(new_n524_), .A3(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n475_), .A2(new_n527_), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n461_), .A2(new_n474_), .A3(new_n524_), .A4(new_n526_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n391_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n499_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n457_), .A2(KEYINPUT32), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT92), .ZN(new_n533_));
  AOI22_X1  g332(.A1(new_n520_), .A2(new_n522_), .B1(new_n452_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT94), .ZN(new_n535_));
  INV_X1    g334(.A(new_n532_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n535_), .B1(new_n471_), .B2(new_n536_), .ZN(new_n537_));
  NOR3_X1   g336(.A1(new_n470_), .A2(KEYINPUT94), .A3(new_n532_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n534_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT95), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT33), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n522_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n509_), .B(KEYINPUT90), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n543_), .A2(new_n505_), .A3(new_n512_), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n544_), .A2(KEYINPUT33), .A3(new_n507_), .A4(new_n521_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n521_), .B1(new_n503_), .B2(new_n505_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n512_), .A2(new_n506_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n546_), .B1(new_n511_), .B2(new_n547_), .ZN(new_n548_));
  AND3_X1   g347(.A1(new_n542_), .A2(new_n545_), .A3(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n458_), .A2(new_n460_), .ZN(new_n550_));
  AOI22_X1  g349(.A1(new_n549_), .A2(new_n550_), .B1(new_n385_), .B2(new_n390_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT95), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n534_), .B(new_n552_), .C1(new_n537_), .C2(new_n538_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n540_), .A2(new_n551_), .A3(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n528_), .B1(new_n531_), .B2(new_n554_), .ZN(new_n555_));
  NOR4_X1   g354(.A1(new_n325_), .A2(new_n326_), .A3(new_n340_), .A4(new_n555_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n524_), .A2(new_n526_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n556_), .A2(new_n261_), .A3(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT38), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n561_), .B(KEYINPUT97), .Z(new_n562_));
  NOR2_X1   g361(.A1(new_n555_), .A2(new_n258_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n322_), .A2(new_n340_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n292_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT98), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n563_), .A2(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(G1gat), .B1(new_n568_), .B2(new_n557_), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n569_), .B(KEYINPUT99), .Z(new_n570_));
  NAND2_X1  g369(.A1(new_n559_), .A2(new_n560_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n562_), .A2(new_n570_), .A3(new_n571_), .ZN(G1324gat));
  INV_X1    g371(.A(KEYINPUT39), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n461_), .A2(new_n474_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  OAI211_X1 g374(.A(new_n573_), .B(G8gat), .C1(new_n568_), .C2(new_n575_), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n576_), .A2(KEYINPUT100), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(KEYINPUT100), .ZN(new_n578_));
  INV_X1    g377(.A(new_n568_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n262_), .B1(new_n579_), .B2(new_n574_), .ZN(new_n580_));
  OAI211_X1 g379(.A(new_n577_), .B(new_n578_), .C1(new_n573_), .C2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n556_), .A2(new_n262_), .A3(new_n574_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  XOR2_X1   g382(.A(KEYINPUT101), .B(KEYINPUT40), .Z(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n584_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n581_), .A2(new_n582_), .A3(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n587_), .ZN(G1325gat));
  NAND3_X1  g387(.A1(new_n556_), .A2(new_n480_), .A3(new_n499_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT102), .ZN(new_n590_));
  INV_X1    g389(.A(new_n499_), .ZN(new_n591_));
  OAI21_X1  g390(.A(G15gat), .B1(new_n568_), .B2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(KEYINPUT41), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n592_), .A2(KEYINPUT41), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n590_), .A2(new_n593_), .A3(new_n594_), .ZN(G1326gat));
  OAI21_X1  g394(.A(G22gat), .B1(new_n568_), .B2(new_n391_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT42), .ZN(new_n597_));
  INV_X1    g396(.A(G22gat), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n556_), .A2(new_n598_), .A3(new_n530_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(new_n599_), .ZN(G1327gat));
  NAND2_X1  g399(.A1(new_n292_), .A2(new_n258_), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n601_), .B(KEYINPUT103), .Z(new_n602_));
  AND2_X1   g401(.A1(new_n602_), .A2(new_n564_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n531_), .A2(new_n554_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n528_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n603_), .A2(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(G29gat), .B1(new_n607_), .B2(new_n558_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT43), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n606_), .A2(new_n609_), .A3(new_n259_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n259_), .ZN(new_n611_));
  OAI21_X1  g410(.A(KEYINPUT43), .B1(new_n555_), .B2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n564_), .A2(new_n292_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(KEYINPUT44), .B1(new_n613_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT44), .ZN(new_n617_));
  AOI211_X1 g416(.A(new_n617_), .B(new_n614_), .C1(new_n610_), .C2(new_n612_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n558_), .A2(G29gat), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n608_), .B1(new_n619_), .B2(new_n620_), .ZN(G1328gat));
  INV_X1    g420(.A(G36gat), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n607_), .A2(new_n622_), .A3(new_n574_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT45), .ZN(new_n624_));
  NOR3_X1   g423(.A1(new_n616_), .A2(new_n618_), .A3(new_n575_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n624_), .B1(new_n625_), .B2(new_n622_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT46), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(G1329gat));
  INV_X1    g427(.A(G43gat), .ZN(new_n629_));
  INV_X1    g428(.A(new_n607_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n629_), .B1(new_n630_), .B2(new_n591_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT104), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n591_), .A2(new_n629_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n632_), .B1(new_n619_), .B2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n633_), .ZN(new_n635_));
  NOR4_X1   g434(.A1(new_n616_), .A2(new_n618_), .A3(KEYINPUT104), .A4(new_n635_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n631_), .B1(new_n634_), .B2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(KEYINPUT47), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT47), .ZN(new_n639_));
  OAI211_X1 g438(.A(new_n639_), .B(new_n631_), .C1(new_n634_), .C2(new_n636_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n638_), .A2(new_n640_), .ZN(G1330gat));
  NOR3_X1   g440(.A1(new_n616_), .A2(new_n618_), .A3(new_n391_), .ZN(new_n642_));
  INV_X1    g441(.A(G50gat), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n391_), .A2(G50gat), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n644_), .B(KEYINPUT105), .Z(new_n645_));
  OAI22_X1  g444(.A1(new_n642_), .A2(new_n643_), .B1(new_n630_), .B2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT106), .ZN(G1331gat));
  INV_X1    g446(.A(new_n340_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n555_), .A2(KEYINPUT107), .A3(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n649_), .A2(new_n321_), .ZN(new_n650_));
  OAI21_X1  g449(.A(KEYINPUT107), .B1(new_n555_), .B2(new_n648_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n259_), .A2(new_n292_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(G57gat), .B1(new_n655_), .B2(new_n558_), .ZN(new_n656_));
  NOR3_X1   g455(.A1(new_n292_), .A2(new_n321_), .A3(new_n648_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n563_), .A2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n658_), .A2(G57gat), .A3(new_n558_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(KEYINPUT108), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n659_), .A2(KEYINPUT108), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n656_), .B1(new_n660_), .B2(new_n661_), .ZN(G1332gat));
  INV_X1    g461(.A(new_n658_), .ZN(new_n663_));
  OAI21_X1  g462(.A(G64gat), .B1(new_n663_), .B2(new_n575_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT48), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n575_), .A2(G64gat), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT109), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n665_), .B1(new_n654_), .B2(new_n667_), .ZN(G1333gat));
  NAND2_X1  g467(.A1(new_n658_), .A2(new_n499_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(G71gat), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n670_), .A2(KEYINPUT49), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n670_), .A2(KEYINPUT49), .ZN(new_n672_));
  OR2_X1    g471(.A1(new_n591_), .A2(G71gat), .ZN(new_n673_));
  OAI22_X1  g472(.A1(new_n671_), .A2(new_n672_), .B1(new_n654_), .B2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT110), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n674_), .B(new_n675_), .ZN(G1334gat));
  OAI21_X1  g475(.A(G78gat), .B1(new_n663_), .B2(new_n391_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT50), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n391_), .A2(G78gat), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n678_), .B1(new_n654_), .B2(new_n679_), .ZN(G1335gat));
  NAND3_X1  g479(.A1(new_n650_), .A2(new_n602_), .A3(new_n651_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n682_), .A2(new_n229_), .A3(new_n558_), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n565_), .A2(new_n321_), .A3(new_n648_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n613_), .A2(new_n684_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n685_), .A2(new_n558_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n683_), .B1(new_n686_), .B2(new_n229_), .ZN(G1336gat));
  AOI21_X1  g486(.A(G92gat), .B1(new_n682_), .B2(new_n574_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n574_), .A2(G92gat), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n689_), .B(KEYINPUT111), .Z(new_n690_));
  AOI21_X1  g489(.A(new_n688_), .B1(new_n685_), .B2(new_n690_), .ZN(G1337gat));
  OR3_X1    g490(.A1(new_n681_), .A2(new_n237_), .A3(new_n591_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n685_), .A2(new_n499_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(G99gat), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT51), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n695_), .A2(KEYINPUT112), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n692_), .A2(new_n694_), .A3(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(KEYINPUT112), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n697_), .B(new_n698_), .ZN(G1338gat));
  NAND3_X1  g498(.A1(new_n682_), .A2(new_n215_), .A3(new_n530_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n613_), .A2(new_n530_), .A3(new_n684_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT52), .ZN(new_n702_));
  AND3_X1   g501(.A1(new_n701_), .A2(new_n702_), .A3(G106gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n702_), .B1(new_n701_), .B2(G106gat), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n700_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  XOR2_X1   g504(.A(KEYINPUT113), .B(KEYINPUT53), .Z(new_n706_));
  XNOR2_X1  g505(.A(new_n705_), .B(new_n706_), .ZN(G1339gat));
  NOR2_X1   g506(.A1(new_n475_), .A2(new_n591_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n335_), .A2(new_n330_), .ZN(new_n709_));
  OAI211_X1 g508(.A(new_n709_), .B(new_n339_), .C1(new_n330_), .C2(new_n329_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT119), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n710_), .A2(new_n711_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n339_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n336_), .A2(new_n714_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n712_), .A2(new_n713_), .A3(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(new_n317_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT117), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n299_), .A2(new_n718_), .A3(new_n305_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n718_), .B1(new_n299_), .B2(new_n305_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n308_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT55), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n307_), .A2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT116), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n307_), .A2(new_n725_), .A3(new_n722_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n307_), .B2(new_n722_), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n721_), .B(new_n724_), .C1(new_n726_), .C2(new_n727_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n728_), .A2(KEYINPUT118), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT118), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n299_), .A2(new_n305_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(KEYINPUT117), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n299_), .A2(new_n305_), .A3(new_n718_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n723_), .B1(new_n734_), .B2(new_n308_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n307_), .A2(new_n722_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(KEYINPUT116), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n307_), .A2(new_n725_), .A3(new_n722_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n730_), .B1(new_n735_), .B2(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n314_), .B1(new_n729_), .B2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT56), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n728_), .A2(KEYINPUT118), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n735_), .A2(new_n739_), .A3(new_n730_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n746_), .A2(KEYINPUT56), .A3(new_n314_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n717_), .B1(new_n743_), .B2(new_n747_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n259_), .B1(new_n748_), .B2(KEYINPUT58), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT120), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT120), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n751_), .B(new_n259_), .C1(new_n748_), .C2(KEYINPUT58), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n748_), .A2(KEYINPUT58), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n750_), .A2(new_n752_), .A3(new_n753_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n648_), .A2(new_n317_), .ZN(new_n755_));
  AOI21_X1  g554(.A(KEYINPUT56), .B1(new_n746_), .B2(new_n314_), .ZN(new_n756_));
  AOI211_X1 g555(.A(new_n742_), .B(new_n316_), .C1(new_n744_), .C2(new_n745_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n755_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n716_), .A2(new_n318_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n258_), .ZN(new_n761_));
  AOI21_X1  g560(.A(KEYINPUT57), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT57), .ZN(new_n763_));
  AOI211_X1 g562(.A(new_n763_), .B(new_n258_), .C1(new_n758_), .C2(new_n759_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n762_), .A2(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n565_), .B1(new_n754_), .B2(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n290_), .A2(new_n291_), .A3(new_n340_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT114), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n290_), .A2(KEYINPUT114), .A3(new_n291_), .A4(new_n340_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n321_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT115), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n771_), .A2(KEYINPUT115), .A3(new_n321_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n774_), .A2(new_n611_), .A3(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT54), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n774_), .A2(KEYINPUT54), .A3(new_n611_), .A4(new_n775_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n558_), .B(new_n708_), .C1(new_n766_), .C2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(G113gat), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n782_), .A2(new_n783_), .A3(new_n648_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT121), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n785_), .B1(new_n781_), .B2(KEYINPUT122), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n754_), .A2(new_n765_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n292_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n780_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n790_), .A2(KEYINPUT121), .A3(new_n558_), .A4(new_n708_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n786_), .A2(KEYINPUT59), .A3(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT59), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n785_), .B(new_n793_), .C1(new_n781_), .C2(KEYINPUT122), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n340_), .B1(new_n792_), .B2(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n784_), .B1(new_n795_), .B2(new_n783_), .ZN(G1340gat));
  INV_X1    g595(.A(KEYINPUT60), .ZN(new_n797_));
  INV_X1    g596(.A(G120gat), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n322_), .A2(new_n797_), .A3(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n799_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n782_), .A2(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n321_), .B1(new_n792_), .B2(new_n794_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n801_), .B1(new_n802_), .B2(new_n798_), .ZN(G1341gat));
  INV_X1    g602(.A(G127gat), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n782_), .A2(new_n804_), .A3(new_n565_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n292_), .B1(new_n792_), .B2(new_n794_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n805_), .B1(new_n806_), .B2(new_n804_), .ZN(G1342gat));
  INV_X1    g606(.A(G134gat), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n782_), .A2(new_n808_), .A3(new_n258_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n611_), .B1(new_n792_), .B2(new_n794_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n809_), .B1(new_n810_), .B2(new_n808_), .ZN(G1343gat));
  NAND2_X1  g610(.A1(new_n530_), .A2(new_n591_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n812_), .A2(new_n574_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n790_), .A2(new_n558_), .A3(new_n813_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n814_), .A2(new_n340_), .ZN(new_n815_));
  XOR2_X1   g614(.A(new_n815_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g615(.A1(new_n814_), .A2(new_n321_), .ZN(new_n817_));
  XOR2_X1   g616(.A(new_n817_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g617(.A1(new_n814_), .A2(new_n292_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(KEYINPUT61), .B(G155gat), .ZN(new_n820_));
  XOR2_X1   g619(.A(new_n819_), .B(new_n820_), .Z(G1346gat));
  OAI21_X1  g620(.A(G162gat), .B1(new_n814_), .B2(new_n611_), .ZN(new_n822_));
  OR2_X1    g621(.A1(new_n761_), .A2(G162gat), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n822_), .B1(new_n814_), .B2(new_n823_), .ZN(G1347gat));
  NOR3_X1   g623(.A1(new_n575_), .A2(new_n527_), .A3(new_n530_), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n648_), .B(new_n825_), .C1(new_n766_), .C2(new_n780_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(G169gat), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT62), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n826_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n790_), .A2(new_n648_), .A3(new_n408_), .A4(new_n825_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n829_), .A2(new_n830_), .A3(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT123), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n829_), .A2(KEYINPUT123), .A3(new_n830_), .A4(new_n831_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(G1348gat));
  AND2_X1   g635(.A1(new_n790_), .A2(new_n825_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n322_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n565_), .ZN(new_n840_));
  MUX2_X1   g639(.A(new_n434_), .B(G183gat), .S(new_n840_), .Z(G1350gat));
  NAND3_X1  g640(.A1(new_n837_), .A2(new_n412_), .A3(new_n258_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT124), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n837_), .A2(new_n259_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n843_), .B1(new_n844_), .B2(G190gat), .ZN(new_n845_));
  AOI211_X1 g644(.A(KEYINPUT124), .B(new_n398_), .C1(new_n837_), .C2(new_n259_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n842_), .B1(new_n845_), .B2(new_n846_), .ZN(G1351gat));
  NOR3_X1   g646(.A1(new_n812_), .A2(new_n558_), .A3(new_n575_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n790_), .A2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n648_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n322_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g652(.A(KEYINPUT126), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n292_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(KEYINPUT125), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n849_), .A2(new_n856_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n854_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n858_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n849_), .A2(KEYINPUT126), .A3(new_n860_), .A4(new_n856_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n857_), .A2(new_n858_), .ZN(new_n862_));
  AND3_X1   g661(.A1(new_n859_), .A2(new_n861_), .A3(new_n862_), .ZN(G1354gat));
  NAND2_X1  g662(.A1(new_n849_), .A2(new_n258_), .ZN(new_n864_));
  XOR2_X1   g663(.A(KEYINPUT127), .B(G218gat), .Z(new_n865_));
  NOR2_X1   g664(.A1(new_n611_), .A2(new_n865_), .ZN(new_n866_));
  AOI22_X1  g665(.A1(new_n864_), .A2(new_n865_), .B1(new_n849_), .B2(new_n866_), .ZN(G1355gat));
endmodule


