//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1 1 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 1 1 0 0 0 1 1 0 1 0 1 0 1 0 1 1 1 1 0 1 1 0 0 0 1 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n662_, new_n663_, new_n664_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n717_, new_n718_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n762_, new_n763_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n911_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n923_, new_n924_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n958_, new_n959_, new_n961_,
    new_n962_, new_n963_, new_n965_, new_n966_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n973_, new_n974_;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G127gat), .B(G134gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT82), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G113gat), .B(G120gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT83), .ZN(new_n208_));
  INV_X1    g007(.A(new_n206_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n205_), .B(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT83), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213_));
  OR2_X1    g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214_));
  OR2_X1    g013(.A1(G141gat), .A2(G148gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT2), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G141gat), .A2(G148gat), .ZN(new_n217_));
  AOI22_X1  g016(.A1(new_n215_), .A2(KEYINPUT3), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n218_), .B1(KEYINPUT3), .B2(new_n215_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n220_));
  XOR2_X1   g019(.A(new_n220_), .B(KEYINPUT85), .Z(new_n221_));
  OAI211_X1 g020(.A(new_n213_), .B(new_n214_), .C1(new_n219_), .C2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT84), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n223_), .B1(new_n213_), .B2(KEYINPUT1), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n213_), .A2(KEYINPUT1), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(new_n225_), .A3(new_n214_), .ZN(new_n226_));
  NOR3_X1   g025(.A1(new_n213_), .A2(new_n223_), .A3(KEYINPUT1), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n217_), .B(new_n215_), .C1(new_n226_), .C2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n222_), .A2(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n208_), .A2(new_n212_), .A3(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT4), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n207_), .A2(new_n228_), .A3(new_n222_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n231_), .B1(new_n230_), .B2(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n203_), .B1(new_n232_), .B2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G1gat), .B(G29gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(G85gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(KEYINPUT0), .B(G57gat), .ZN(new_n238_));
  XOR2_X1   g037(.A(new_n237_), .B(new_n238_), .Z(new_n239_));
  NAND3_X1  g038(.A1(new_n230_), .A2(new_n202_), .A3(new_n233_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT92), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n230_), .A2(KEYINPUT92), .A3(new_n202_), .A4(new_n233_), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n235_), .A2(new_n239_), .A3(new_n242_), .A4(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT94), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n242_), .A2(new_n243_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n248_), .A2(KEYINPUT94), .A3(new_n239_), .A4(new_n235_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n239_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n235_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n250_), .B1(new_n251_), .B2(new_n247_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n246_), .A2(new_n249_), .A3(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT95), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G183gat), .A2(G190gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT23), .ZN(new_n256_));
  INV_X1    g055(.A(G169gat), .ZN(new_n257_));
  INV_X1    g056(.A(G176gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  OR2_X1    g058(.A1(new_n259_), .A2(KEYINPUT24), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n256_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT79), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G169gat), .A2(G176gat), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n259_), .A2(KEYINPUT24), .A3(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(G183gat), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n266_), .A2(KEYINPUT25), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT77), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n266_), .A2(KEYINPUT25), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n267_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(G190gat), .ZN(new_n271_));
  OR3_X1    g070(.A1(new_n271_), .A2(KEYINPUT78), .A3(KEYINPUT26), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n266_), .A2(KEYINPUT77), .A3(KEYINPUT25), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT26), .B1(new_n271_), .B2(KEYINPUT78), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n270_), .A2(new_n272_), .A3(new_n273_), .A4(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n256_), .A2(new_n260_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(KEYINPUT79), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n263_), .A2(new_n265_), .A3(new_n275_), .A4(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT22), .B(G169gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(new_n258_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT80), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n256_), .B1(G183gat), .B2(G190gat), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n281_), .A2(new_n282_), .A3(new_n264_), .ZN(new_n283_));
  AND2_X1   g082(.A1(new_n278_), .A2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT30), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT81), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G71gat), .B(G99gat), .ZN(new_n288_));
  INV_X1    g087(.A(G43gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G227gat), .A2(G233gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(G15gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n290_), .B(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n287_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(KEYINPUT31), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n278_), .A2(new_n283_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT30), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT81), .ZN(new_n298_));
  AND2_X1   g097(.A1(new_n208_), .A2(new_n212_), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT31), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n287_), .A2(new_n301_), .A3(new_n293_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n298_), .A2(new_n299_), .ZN(new_n303_));
  AND4_X1   g102(.A1(new_n295_), .A2(new_n300_), .A3(new_n302_), .A4(new_n303_), .ZN(new_n304_));
  AOI22_X1  g103(.A1(new_n295_), .A2(new_n302_), .B1(new_n300_), .B2(new_n303_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT95), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n246_), .A2(new_n249_), .A3(new_n252_), .A4(new_n307_), .ZN(new_n308_));
  AND3_X1   g107(.A1(new_n254_), .A2(new_n306_), .A3(new_n308_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n229_), .A2(KEYINPUT29), .ZN(new_n310_));
  XOR2_X1   g109(.A(new_n310_), .B(KEYINPUT28), .Z(new_n311_));
  XOR2_X1   g110(.A(G211gat), .B(G218gat), .Z(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT87), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT21), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G197gat), .B(G204gat), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n314_), .B1(new_n315_), .B2(KEYINPUT88), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n316_), .B1(KEYINPUT88), .B2(new_n315_), .ZN(new_n317_));
  OR2_X1    g116(.A1(new_n313_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(G197gat), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n319_), .A2(KEYINPUT86), .A3(G204gat), .ZN(new_n320_));
  INV_X1    g119(.A(new_n315_), .ZN(new_n321_));
  OAI211_X1 g120(.A(KEYINPUT21), .B(new_n320_), .C1(new_n321_), .C2(KEYINPUT86), .ZN(new_n322_));
  OAI211_X1 g121(.A(new_n313_), .B(new_n322_), .C1(KEYINPUT21), .C2(new_n321_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n318_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n325_), .B1(KEYINPUT29), .B2(new_n229_), .ZN(new_n326_));
  OR2_X1    g125(.A1(new_n311_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n311_), .A2(new_n326_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G228gat), .A2(G233gat), .ZN(new_n330_));
  INV_X1    g129(.A(G78gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(G106gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G22gat), .B(G50gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n329_), .A2(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n327_), .A2(new_n328_), .A3(new_n336_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n325_), .A2(new_n284_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n264_), .B(KEYINPUT91), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n282_), .A2(new_n280_), .A3(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT26), .B(G190gat), .ZN(new_n346_));
  OR2_X1    g145(.A1(new_n266_), .A2(KEYINPUT25), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n346_), .A2(new_n347_), .A3(new_n269_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n261_), .A2(new_n265_), .A3(new_n348_), .ZN(new_n349_));
  OR2_X1    g148(.A1(new_n349_), .A2(KEYINPUT90), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(KEYINPUT90), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n345_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  OAI211_X1 g151(.A(new_n342_), .B(KEYINPUT20), .C1(new_n325_), .C2(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G226gat), .A2(G233gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n353_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G8gat), .B(G36gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT18), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G64gat), .B(G92gat), .ZN(new_n360_));
  XOR2_X1   g159(.A(new_n359_), .B(new_n360_), .Z(new_n361_));
  NAND2_X1  g160(.A1(new_n352_), .A2(new_n325_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n356_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT20), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n364_), .B1(new_n296_), .B2(new_n324_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n362_), .A2(new_n363_), .A3(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n357_), .A2(new_n361_), .A3(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT27), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n350_), .A2(new_n351_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(new_n344_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n364_), .B1(new_n370_), .B2(new_n324_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n371_), .A2(new_n363_), .A3(new_n342_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n325_), .A2(new_n344_), .A3(new_n349_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n363_), .B1(new_n373_), .B2(new_n365_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n361_), .B1(new_n372_), .B2(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n368_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT96), .ZN(new_n379_));
  INV_X1    g178(.A(new_n361_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n363_), .B1(new_n371_), .B2(new_n342_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n366_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n380_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(new_n367_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT27), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n379_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  AOI211_X1 g185(.A(KEYINPUT96), .B(KEYINPUT27), .C1(new_n383_), .C2(new_n367_), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n341_), .B(new_n378_), .C1(new_n386_), .C2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT97), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n309_), .A2(new_n389_), .A3(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n254_), .A2(new_n306_), .A3(new_n308_), .ZN(new_n392_));
  OAI21_X1  g191(.A(KEYINPUT97), .B1(new_n392_), .B2(new_n388_), .ZN(new_n393_));
  NOR3_X1   g192(.A1(new_n381_), .A2(new_n382_), .A3(new_n380_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n361_), .B1(new_n357_), .B2(new_n366_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT33), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n244_), .A2(new_n397_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n202_), .B1(new_n232_), .B2(new_n234_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n230_), .A2(new_n233_), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n399_), .B(new_n250_), .C1(new_n202_), .C2(new_n400_), .ZN(new_n401_));
  AND3_X1   g200(.A1(new_n396_), .A2(new_n398_), .A3(new_n401_), .ZN(new_n402_));
  OR2_X1    g201(.A1(new_n244_), .A2(new_n397_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT93), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n361_), .A2(KEYINPUT32), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n353_), .A2(new_n356_), .ZN(new_n407_));
  OAI211_X1 g206(.A(new_n404_), .B(new_n406_), .C1(new_n407_), .C2(new_n374_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n357_), .A2(new_n405_), .A3(new_n366_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n372_), .A2(new_n375_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n404_), .B1(new_n411_), .B2(new_n406_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n410_), .A2(new_n412_), .ZN(new_n413_));
  AOI22_X1  g212(.A1(new_n402_), .A2(new_n403_), .B1(new_n253_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n254_), .A2(new_n308_), .ZN(new_n415_));
  OAI211_X1 g214(.A(new_n340_), .B(new_n378_), .C1(new_n386_), .C2(new_n387_), .ZN(new_n416_));
  OAI22_X1  g215(.A1(new_n414_), .A2(new_n340_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n306_), .ZN(new_n418_));
  AOI22_X1  g217(.A1(new_n391_), .A2(new_n393_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G113gat), .B(G141gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(KEYINPUT75), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G169gat), .B(G197gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  XOR2_X1   g223(.A(G1gat), .B(G8gat), .Z(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  OR2_X1    g225(.A1(G15gat), .A2(G22gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G15gat), .A2(G22gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G1gat), .A2(G8gat), .ZN(new_n429_));
  AOI22_X1  g228(.A1(new_n427_), .A2(new_n428_), .B1(KEYINPUT14), .B2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT73), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  AND2_X1   g231(.A1(G15gat), .A2(G22gat), .ZN(new_n433_));
  NOR2_X1   g232(.A1(G15gat), .A2(G22gat), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT14), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n436_), .B1(G1gat), .B2(G8gat), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT73), .B1(new_n435_), .B2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT74), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n432_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n439_), .B1(new_n432_), .B2(new_n438_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n426_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n430_), .A2(new_n431_), .ZN(new_n444_));
  NOR3_X1   g243(.A1(new_n435_), .A2(new_n437_), .A3(KEYINPUT73), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT74), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n446_), .A2(new_n425_), .A3(new_n440_), .ZN(new_n447_));
  INV_X1    g246(.A(G36gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(G29gat), .ZN(new_n449_));
  INV_X1    g248(.A(G29gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(G36gat), .ZN(new_n451_));
  AOI21_X1  g250(.A(KEYINPUT70), .B1(new_n449_), .B2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n449_), .A2(new_n451_), .A3(KEYINPUT70), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G43gat), .B(G50gat), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n453_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n455_), .ZN(new_n457_));
  AND3_X1   g256(.A1(new_n449_), .A2(new_n451_), .A3(KEYINPUT70), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n457_), .B1(new_n458_), .B2(new_n452_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n456_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n443_), .A2(new_n447_), .A3(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G229gat), .A2(G233gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT15), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n460_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n456_), .A2(new_n459_), .A3(KEYINPUT15), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n467_), .B1(new_n447_), .B2(new_n443_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n463_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n460_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n447_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n425_), .B1(new_n446_), .B2(new_n440_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n470_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n462_), .B1(new_n473_), .B2(new_n461_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n424_), .B1(new_n469_), .B2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT76), .ZN(new_n476_));
  INV_X1    g275(.A(new_n462_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n461_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n460_), .B1(new_n443_), .B2(new_n447_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n477_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n471_), .A2(new_n472_), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n461_), .B(new_n462_), .C1(new_n481_), .C2(new_n467_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n480_), .A2(new_n482_), .A3(new_n423_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n475_), .A2(new_n476_), .A3(new_n483_), .ZN(new_n484_));
  OAI211_X1 g283(.A(KEYINPUT76), .B(new_n424_), .C1(new_n469_), .C2(new_n474_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n419_), .A2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G120gat), .B(G148gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(KEYINPUT5), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G176gat), .B(G204gat), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n489_), .B(new_n490_), .Z(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT65), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G57gat), .B(G64gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G71gat), .B(G78gat), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n494_), .A2(new_n495_), .A3(KEYINPUT11), .ZN(new_n496_));
  INV_X1    g295(.A(G64gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(G57gat), .ZN(new_n498_));
  INV_X1    g297(.A(G57gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(G64gat), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n498_), .A2(new_n500_), .A3(KEYINPUT11), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n331_), .A2(G71gat), .ZN(new_n502_));
  INV_X1    g301(.A(G71gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(G78gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n502_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n501_), .A2(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(KEYINPUT11), .B1(new_n498_), .B2(new_n500_), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n493_), .B(new_n496_), .C1(new_n506_), .C2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT12), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n498_), .A2(new_n500_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT11), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n512_), .A2(new_n501_), .A3(new_n505_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n493_), .B1(new_n513_), .B2(new_n496_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n509_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(G85gat), .ZN(new_n516_));
  INV_X1    g315(.A(G92gat), .ZN(new_n517_));
  NOR3_X1   g316(.A1(new_n516_), .A2(new_n517_), .A3(KEYINPUT9), .ZN(new_n518_));
  AND2_X1   g317(.A1(G85gat), .A2(G92gat), .ZN(new_n519_));
  NOR2_X1   g318(.A1(G85gat), .A2(G92gat), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n518_), .B1(KEYINPUT9), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT64), .ZN(new_n523_));
  OR2_X1    g322(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n523_), .B1(new_n526_), .B2(G106gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G99gat), .A2(G106gat), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT6), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT6), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n530_), .A2(G99gat), .A3(G106gat), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n529_), .A2(new_n531_), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n524_), .A2(KEYINPUT64), .A3(new_n333_), .A4(new_n525_), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n522_), .A2(new_n527_), .A3(new_n532_), .A4(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G85gat), .B(G92gat), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NOR3_X1   g336(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  AOI211_X1 g338(.A(KEYINPUT8), .B(new_n535_), .C1(new_n539_), .C2(new_n532_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT8), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT7), .ZN(new_n542_));
  INV_X1    g341(.A(G99gat), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n542_), .A2(new_n543_), .A3(new_n333_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n530_), .B1(G99gat), .B2(G106gat), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n528_), .A2(KEYINPUT6), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n536_), .B(new_n544_), .C1(new_n545_), .C2(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n541_), .B1(new_n547_), .B2(new_n521_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n534_), .B1(new_n540_), .B2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n515_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(KEYINPUT66), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G230gat), .A2(G233gat), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n549_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n513_), .A2(new_n496_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n553_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n555_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n549_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT12), .ZN(new_n559_));
  AOI22_X1  g358(.A1(new_n558_), .A2(new_n559_), .B1(new_n515_), .B2(new_n549_), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n551_), .B(new_n556_), .C1(new_n560_), .C2(KEYINPUT66), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n554_), .A2(new_n555_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n558_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n553_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n492_), .B1(new_n561_), .B2(new_n565_), .ZN(new_n566_));
  XOR2_X1   g365(.A(new_n566_), .B(KEYINPUT67), .Z(new_n567_));
  NAND3_X1  g366(.A1(new_n561_), .A2(new_n565_), .A3(new_n492_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(KEYINPUT68), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT68), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n561_), .A2(new_n565_), .A3(new_n570_), .A4(new_n492_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n567_), .A2(new_n572_), .ZN(new_n573_));
  XOR2_X1   g372(.A(KEYINPUT69), .B(KEYINPUT13), .Z(new_n574_));
  OR2_X1    g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n573_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n575_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n554_), .A2(new_n460_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n467_), .A2(new_n554_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G232gat), .A2(G233gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT34), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n584_), .A2(KEYINPUT35), .ZN(new_n585_));
  NOR3_X1   g384(.A1(new_n581_), .A2(new_n582_), .A3(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(KEYINPUT35), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  OAI211_X1 g387(.A(KEYINPUT35), .B(new_n584_), .C1(new_n581_), .C2(new_n582_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G190gat), .B(G218gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G134gat), .B(G162gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n593_), .B(KEYINPUT36), .Z(new_n594_));
  NAND2_X1  g393(.A1(new_n590_), .A2(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n593_), .A2(KEYINPUT36), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n588_), .A2(new_n589_), .A3(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(KEYINPUT37), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(KEYINPUT71), .ZN(new_n600_));
  INV_X1    g399(.A(new_n594_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n601_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n602_), .A2(KEYINPUT72), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT37), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(KEYINPUT72), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n603_), .A2(new_n604_), .A3(new_n597_), .A4(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT71), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n598_), .A2(new_n607_), .A3(KEYINPUT37), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n600_), .A2(new_n606_), .A3(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(G231gat), .A2(G233gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n481_), .B(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(new_n557_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G127gat), .B(G155gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT16), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G183gat), .B(G211gat), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n615_), .B(new_n616_), .Z(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n618_), .A2(KEYINPUT17), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT17), .ZN(new_n620_));
  NOR3_X1   g419(.A1(new_n617_), .A2(new_n493_), .A3(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n613_), .B1(new_n619_), .B2(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n622_), .B1(new_n613_), .B2(new_n621_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n610_), .A2(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n579_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n487_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n415_), .ZN(new_n627_));
  OR3_X1    g426(.A1(new_n626_), .A2(G1gat), .A3(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT38), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n603_), .A2(new_n597_), .A3(new_n605_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n419_), .A2(new_n632_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n484_), .A2(new_n485_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n578_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n623_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n633_), .A2(new_n637_), .ZN(new_n638_));
  OAI21_X1  g437(.A(G1gat), .B1(new_n638_), .B2(new_n627_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n628_), .A2(new_n629_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n630_), .A2(new_n639_), .A3(new_n640_), .ZN(G1324gat));
  INV_X1    g440(.A(KEYINPUT39), .ZN(new_n642_));
  INV_X1    g441(.A(new_n638_), .ZN(new_n643_));
  OAI21_X1  g442(.A(KEYINPUT96), .B1(new_n396_), .B2(KEYINPUT27), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n384_), .A2(new_n379_), .A3(new_n385_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n377_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n643_), .A2(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n642_), .B1(new_n648_), .B2(G8gat), .ZN(new_n649_));
  INV_X1    g448(.A(G8gat), .ZN(new_n650_));
  AOI211_X1 g449(.A(KEYINPUT39), .B(new_n650_), .C1(new_n643_), .C2(new_n647_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n647_), .A2(new_n650_), .ZN(new_n652_));
  OAI22_X1  g451(.A1(new_n649_), .A2(new_n651_), .B1(new_n626_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT40), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n653_), .B(new_n654_), .ZN(G1325gat));
  NOR3_X1   g454(.A1(new_n626_), .A2(G15gat), .A3(new_n418_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT98), .ZN(new_n657_));
  OAI21_X1  g456(.A(G15gat), .B1(new_n638_), .B2(new_n418_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(KEYINPUT41), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n658_), .A2(KEYINPUT41), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n657_), .A2(new_n659_), .A3(new_n660_), .ZN(G1326gat));
  OAI21_X1  g460(.A(G22gat), .B1(new_n638_), .B2(new_n341_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT42), .ZN(new_n663_));
  OR2_X1    g462(.A1(new_n341_), .A2(G22gat), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n663_), .B1(new_n626_), .B2(new_n664_), .ZN(G1327gat));
  OAI21_X1  g464(.A(KEYINPUT43), .B1(new_n419_), .B2(new_n610_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT43), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n390_), .B1(new_n309_), .B2(new_n389_), .ZN(new_n668_));
  NOR3_X1   g467(.A1(new_n392_), .A2(new_n388_), .A3(KEYINPUT97), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  OR2_X1    g469(.A1(new_n415_), .A2(new_n416_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n402_), .A2(new_n403_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n253_), .A2(new_n413_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(new_n341_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n306_), .B1(new_n671_), .B2(new_n675_), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n667_), .B(new_n609_), .C1(new_n670_), .C2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n666_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT44), .ZN(new_n679_));
  AOI211_X1 g478(.A(new_n623_), .B(new_n635_), .C1(KEYINPUT99), .C2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT99), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n681_), .A2(new_n682_), .A3(KEYINPUT44), .ZN(new_n683_));
  OAI211_X1 g482(.A(new_n678_), .B(new_n680_), .C1(KEYINPUT99), .C2(new_n679_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n450_), .B1(new_n685_), .B2(new_n415_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n636_), .A2(new_n632_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n579_), .A2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n487_), .A2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n415_), .A2(new_n450_), .ZN(new_n690_));
  XOR2_X1   g489(.A(new_n690_), .B(KEYINPUT100), .Z(new_n691_));
  NOR2_X1   g490(.A1(new_n689_), .A2(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(KEYINPUT101), .B1(new_n686_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT101), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n627_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n695_));
  OAI221_X1 g494(.A(new_n694_), .B1(new_n689_), .B2(new_n691_), .C1(new_n695_), .C2(new_n450_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n693_), .A2(new_n696_), .ZN(G1328gat));
  INV_X1    g496(.A(KEYINPUT46), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n448_), .B1(new_n685_), .B2(new_n647_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n689_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n646_), .B(KEYINPUT102), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n700_), .A2(new_n448_), .A3(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT45), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n703_), .B(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n698_), .B1(new_n699_), .B2(new_n705_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n703_), .B(KEYINPUT45), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n646_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n708_));
  OAI211_X1 g507(.A(new_n707_), .B(KEYINPUT46), .C1(new_n448_), .C2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n706_), .A2(new_n709_), .ZN(G1329gat));
  NOR2_X1   g509(.A1(new_n418_), .A2(new_n289_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n685_), .A2(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n289_), .B1(new_n689_), .B2(new_n418_), .ZN(new_n713_));
  AND3_X1   g512(.A1(new_n712_), .A2(KEYINPUT47), .A3(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(KEYINPUT47), .B1(new_n712_), .B2(new_n713_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1330gat));
  AOI21_X1  g515(.A(G50gat), .B1(new_n700_), .B2(new_n340_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n340_), .A2(G50gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n685_), .B2(new_n718_), .ZN(G1331gat));
  NOR2_X1   g518(.A1(new_n419_), .A2(new_n634_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n624_), .A2(new_n578_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(KEYINPUT103), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT103), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n627_), .B1(new_n722_), .B2(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(G57gat), .B1(new_n724_), .B2(new_n726_), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n633_), .A2(new_n486_), .A3(new_n579_), .A4(new_n623_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT104), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n728_), .B(new_n729_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n627_), .A2(new_n499_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n727_), .B1(new_n730_), .B2(new_n731_), .ZN(G1332gat));
  NAND3_X1  g531(.A1(new_n723_), .A2(new_n497_), .A3(new_n702_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n728_), .B(KEYINPUT104), .ZN(new_n734_));
  OAI21_X1  g533(.A(G64gat), .B1(new_n734_), .B2(new_n701_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n735_), .A2(KEYINPUT48), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n735_), .A2(KEYINPUT48), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n733_), .B1(new_n736_), .B2(new_n737_), .ZN(G1333gat));
  NAND3_X1  g537(.A1(new_n723_), .A2(new_n503_), .A3(new_n306_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n730_), .A2(new_n306_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(KEYINPUT105), .B(KEYINPUT49), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n740_), .A2(G71gat), .A3(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n740_), .B2(G71gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n739_), .B1(new_n742_), .B2(new_n743_), .ZN(G1334gat));
  NAND3_X1  g543(.A1(new_n723_), .A2(new_n331_), .A3(new_n340_), .ZN(new_n745_));
  OAI21_X1  g544(.A(G78gat), .B1(new_n734_), .B2(new_n341_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n746_), .A2(KEYINPUT50), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n746_), .A2(KEYINPUT50), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n745_), .B1(new_n747_), .B2(new_n748_), .ZN(G1335gat));
  NOR2_X1   g548(.A1(new_n578_), .A2(new_n687_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n720_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n752_), .A2(new_n516_), .A3(new_n415_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n623_), .A2(new_n634_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n579_), .A2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n678_), .A2(KEYINPUT106), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT106), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n666_), .A2(new_n677_), .A3(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n755_), .B1(new_n756_), .B2(new_n758_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n759_), .A2(new_n415_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n753_), .B1(new_n760_), .B2(new_n516_), .ZN(G1336gat));
  NAND3_X1  g560(.A1(new_n752_), .A2(new_n517_), .A3(new_n647_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n759_), .A2(new_n702_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n762_), .B1(new_n763_), .B2(new_n517_), .ZN(G1337gat));
  NAND2_X1  g563(.A1(new_n756_), .A2(new_n758_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n755_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n765_), .A2(new_n306_), .A3(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(G99gat), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT107), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n751_), .A2(new_n418_), .A3(new_n526_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n768_), .A2(new_n769_), .A3(KEYINPUT51), .A4(new_n771_), .ZN(new_n772_));
  OR2_X1    g571(.A1(new_n769_), .A2(KEYINPUT51), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n769_), .A2(KEYINPUT51), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n543_), .B1(new_n759_), .B2(new_n306_), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n773_), .B(new_n774_), .C1(new_n775_), .C2(new_n770_), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n772_), .A2(new_n776_), .ZN(G1338gat));
  NAND3_X1  g576(.A1(new_n752_), .A2(new_n333_), .A3(new_n340_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n755_), .A2(new_n341_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n780_), .B1(new_n666_), .B2(new_n677_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n333_), .B1(new_n781_), .B2(KEYINPUT108), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n678_), .A2(new_n779_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT108), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n782_), .A2(new_n785_), .A3(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n782_), .B2(new_n785_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n778_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(KEYINPUT109), .B(KEYINPUT53), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n791_), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n778_), .B(new_n790_), .C1(new_n787_), .C2(new_n788_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(G1339gat));
  NOR3_X1   g593(.A1(new_n627_), .A2(new_n418_), .A3(new_n388_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT59), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT115), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n798_), .A2(KEYINPUT57), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n462_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n461_), .A2(new_n477_), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n800_), .B(new_n424_), .C1(new_n468_), .C2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n483_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n803_), .B1(new_n567_), .B2(new_n572_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805_));
  OAI21_X1  g604(.A(KEYINPUT114), .B1(new_n561_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT66), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n807_), .B1(new_n515_), .B2(new_n549_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n550_), .B1(new_n564_), .B2(KEYINPUT12), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n808_), .B1(new_n809_), .B2(new_n807_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT114), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n810_), .A2(new_n811_), .A3(KEYINPUT55), .A4(new_n556_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT112), .ZN(new_n813_));
  AND3_X1   g612(.A1(new_n561_), .A2(new_n813_), .A3(new_n805_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n813_), .B1(new_n561_), .B2(new_n805_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n806_), .B(new_n812_), .C1(new_n814_), .C2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT113), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n810_), .A2(new_n817_), .A3(new_n562_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n551_), .B1(new_n560_), .B2(KEYINPUT66), .ZN(new_n819_));
  OAI21_X1  g618(.A(KEYINPUT113), .B1(new_n819_), .B2(new_n563_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n552_), .B1(new_n818_), .B2(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n491_), .B1(new_n816_), .B2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT56), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  OAI211_X1 g623(.A(KEYINPUT56), .B(new_n491_), .C1(new_n816_), .C2(new_n821_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n569_), .A2(new_n571_), .ZN(new_n827_));
  NOR3_X1   g626(.A1(new_n827_), .A2(new_n486_), .A3(KEYINPUT111), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT111), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n829_), .B1(new_n634_), .B2(new_n572_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n828_), .A2(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n804_), .B1(new_n826_), .B2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n799_), .B1(new_n832_), .B2(new_n632_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n799_), .ZN(new_n834_));
  OAI21_X1  g633(.A(KEYINPUT111), .B1(new_n827_), .B2(new_n486_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n634_), .A2(new_n829_), .A3(new_n572_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n837_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n631_), .B(new_n834_), .C1(new_n838_), .C2(new_n804_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n833_), .A2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n572_), .A2(new_n483_), .A3(new_n802_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n842_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n609_), .B1(new_n843_), .B2(KEYINPUT58), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(KEYINPUT116), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(KEYINPUT58), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT116), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n609_), .B(new_n847_), .C1(new_n843_), .C2(KEYINPUT58), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n845_), .A2(new_n846_), .A3(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n841_), .A2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n636_), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n578_), .A2(new_n486_), .A3(new_n623_), .A4(new_n610_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(KEYINPUT110), .B(KEYINPUT54), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n852_), .B(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n797_), .B1(new_n851_), .B2(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n840_), .B1(new_n849_), .B2(KEYINPUT117), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT117), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n845_), .A2(new_n859_), .A3(new_n846_), .A4(new_n848_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n623_), .B1(new_n858_), .B2(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n795_), .B1(new_n861_), .B2(new_n855_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n857_), .B1(new_n862_), .B2(KEYINPUT59), .ZN(new_n863_));
  INV_X1    g662(.A(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(G113gat), .B1(new_n864_), .B2(new_n486_), .ZN(new_n865_));
  OR2_X1    g664(.A1(new_n486_), .A2(G113gat), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(new_n862_), .B2(new_n866_), .ZN(G1340gat));
  NAND2_X1  g666(.A1(new_n851_), .A2(new_n856_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n868_), .A2(new_n796_), .A3(new_n795_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n795_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n849_), .A2(KEYINPUT117), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n871_), .A2(new_n841_), .A3(new_n860_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n636_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n870_), .B1(new_n873_), .B2(new_n856_), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n869_), .B(new_n579_), .C1(new_n874_), .C2(new_n796_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(KEYINPUT118), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n863_), .A2(new_n877_), .A3(new_n579_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n876_), .A2(G120gat), .A3(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(G120gat), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n880_), .B1(new_n578_), .B2(KEYINPUT60), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n874_), .B(new_n881_), .C1(KEYINPUT60), .C2(new_n880_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n879_), .A2(new_n882_), .ZN(G1341gat));
  INV_X1    g682(.A(KEYINPUT119), .ZN(new_n884_));
  INV_X1    g683(.A(G127gat), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n885_), .B1(new_n863_), .B2(new_n623_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n862_), .A2(G127gat), .A3(new_n636_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n884_), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n869_), .B(new_n623_), .C1(new_n874_), .C2(new_n796_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(G127gat), .ZN(new_n890_));
  INV_X1    g689(.A(new_n887_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n890_), .A2(KEYINPUT119), .A3(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n888_), .A2(new_n892_), .ZN(G1342gat));
  OAI21_X1  g692(.A(G134gat), .B1(new_n864_), .B2(new_n610_), .ZN(new_n894_));
  OR2_X1    g693(.A1(new_n631_), .A2(G134gat), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n862_), .B2(new_n895_), .ZN(G1343gat));
  XNOR2_X1  g695(.A(KEYINPUT120), .B(G141gat), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n855_), .B1(new_n872_), .B2(new_n636_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n306_), .A2(new_n341_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n701_), .A2(new_n415_), .A3(new_n900_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n899_), .A2(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT121), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n902_), .A2(new_n903_), .A3(new_n634_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n903_), .B1(new_n902_), .B2(new_n634_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n898_), .B1(new_n905_), .B2(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n906_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n908_), .A2(new_n904_), .A3(new_n897_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n907_), .A2(new_n909_), .ZN(G1344gat));
  NAND2_X1  g709(.A1(new_n902_), .A2(new_n579_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g711(.A(KEYINPUT122), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n873_), .A2(new_n856_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n901_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n913_), .B1(new_n916_), .B2(new_n636_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n902_), .A2(KEYINPUT122), .A3(new_n623_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(KEYINPUT61), .B(G155gat), .ZN(new_n919_));
  AND3_X1   g718(.A1(new_n917_), .A2(new_n918_), .A3(new_n919_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n919_), .B1(new_n917_), .B2(new_n918_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n920_), .A2(new_n921_), .ZN(G1346gat));
  OR3_X1    g721(.A1(new_n916_), .A2(G162gat), .A3(new_n631_), .ZN(new_n923_));
  OAI21_X1  g722(.A(G162gat), .B1(new_n916_), .B2(new_n610_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(new_n924_), .ZN(G1347gat));
  NOR2_X1   g724(.A1(new_n701_), .A2(new_n392_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(KEYINPUT123), .ZN(new_n927_));
  NAND4_X1  g726(.A1(new_n868_), .A2(new_n341_), .A3(new_n634_), .A4(new_n927_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n928_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n927_), .A2(new_n341_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n930_), .B1(new_n856_), .B2(new_n851_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n931_), .A2(new_n279_), .A3(new_n634_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n929_), .A2(new_n932_), .ZN(new_n933_));
  AOI21_X1  g732(.A(KEYINPUT62), .B1(new_n928_), .B2(G169gat), .ZN(new_n934_));
  OAI21_X1  g733(.A(KEYINPUT124), .B1(new_n933_), .B2(new_n934_), .ZN(new_n935_));
  INV_X1    g734(.A(new_n934_), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT124), .ZN(new_n937_));
  NAND4_X1  g736(.A1(new_n936_), .A2(new_n937_), .A3(new_n932_), .A4(new_n929_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n935_), .A2(new_n938_), .ZN(G1348gat));
  AOI21_X1  g738(.A(G176gat), .B1(new_n931_), .B2(new_n579_), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT125), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n941_), .B1(new_n899_), .B2(new_n340_), .ZN(new_n942_));
  OAI211_X1 g741(.A(KEYINPUT125), .B(new_n341_), .C1(new_n861_), .C2(new_n855_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n942_), .A2(new_n943_), .ZN(new_n944_));
  INV_X1    g743(.A(new_n927_), .ZN(new_n945_));
  NOR3_X1   g744(.A1(new_n945_), .A2(new_n258_), .A3(new_n578_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n940_), .B1(new_n944_), .B2(new_n946_), .ZN(G1349gat));
  NAND3_X1  g746(.A1(new_n868_), .A2(new_n341_), .A3(new_n927_), .ZN(new_n948_));
  AOI211_X1 g747(.A(new_n636_), .B(new_n948_), .C1(new_n347_), .C2(new_n269_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n945_), .A2(new_n636_), .ZN(new_n950_));
  INV_X1    g749(.A(new_n950_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n951_), .B1(new_n942_), .B2(new_n943_), .ZN(new_n952_));
  AOI21_X1  g751(.A(G183gat), .B1(new_n952_), .B2(KEYINPUT126), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n944_), .A2(new_n950_), .ZN(new_n954_));
  INV_X1    g753(.A(KEYINPUT126), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n954_), .A2(new_n955_), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n949_), .B1(new_n953_), .B2(new_n956_), .ZN(G1350gat));
  OAI21_X1  g756(.A(G190gat), .B1(new_n948_), .B2(new_n610_), .ZN(new_n958_));
  NAND3_X1  g757(.A1(new_n931_), .A2(new_n346_), .A3(new_n632_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n958_), .A2(new_n959_), .ZN(G1351gat));
  NOR4_X1   g759(.A1(new_n701_), .A2(new_n306_), .A3(new_n341_), .A4(new_n415_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n914_), .A2(new_n961_), .ZN(new_n962_));
  NOR2_X1   g761(.A1(new_n962_), .A2(new_n486_), .ZN(new_n963_));
  XNOR2_X1  g762(.A(new_n963_), .B(new_n319_), .ZN(G1352gat));
  INV_X1    g763(.A(new_n962_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n965_), .A2(new_n579_), .ZN(new_n966_));
  XNOR2_X1  g765(.A(new_n966_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g766(.A(new_n636_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n965_), .A2(new_n968_), .ZN(new_n969_));
  NOR2_X1   g768(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n970_));
  XNOR2_X1  g769(.A(new_n970_), .B(KEYINPUT127), .ZN(new_n971_));
  XNOR2_X1  g770(.A(new_n969_), .B(new_n971_), .ZN(G1354gat));
  OR3_X1    g771(.A1(new_n962_), .A2(G218gat), .A3(new_n631_), .ZN(new_n973_));
  OAI21_X1  g772(.A(G218gat), .B1(new_n962_), .B2(new_n610_), .ZN(new_n974_));
  NAND2_X1  g773(.A1(new_n973_), .A2(new_n974_), .ZN(G1355gat));
endmodule


