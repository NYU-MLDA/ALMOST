//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 0 1 1 1 1 1 0 0 0 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0 0 1 0 0 0 1 1 0 0 1 1 0 0 1 1 1 0 1 0 0 0 0 1 1 1 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n685_, new_n686_, new_n687_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n694_, new_n695_, new_n696_, new_n697_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n848_, new_n849_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n879_, new_n880_, new_n882_,
    new_n883_, new_n884_, new_n886_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XOR2_X1   g002(.A(KEYINPUT10), .B(G99gat), .Z(new_n204_));
  INV_X1    g003(.A(G106gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  AND3_X1   g005(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n207_));
  AOI21_X1  g006(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  AOI21_X1  g008(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G85gat), .B(G92gat), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n210_), .B1(new_n211_), .B2(KEYINPUT9), .ZN(new_n212_));
  AND2_X1   g011(.A1(new_n212_), .A2(KEYINPUT64), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n212_), .A2(KEYINPUT64), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n206_), .B(new_n209_), .C1(new_n213_), .C2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT65), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT7), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n216_), .B(new_n217_), .C1(G99gat), .C2(G106gat), .ZN(new_n218_));
  INV_X1    g017(.A(G99gat), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n219_), .B(new_n205_), .C1(KEYINPUT65), .C2(KEYINPUT7), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(new_n209_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n211_), .ZN(new_n223_));
  OR2_X1    g022(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n224_));
  NAND2_X1  g023(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .A4(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT8), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT67), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n228_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G99gat), .A2(G106gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT6), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n232_), .A2(KEYINPUT67), .A3(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n221_), .A2(new_n229_), .A3(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n227_), .B1(new_n235_), .B2(new_n223_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT68), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n226_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  AOI211_X1 g037(.A(KEYINPUT68), .B(new_n227_), .C1(new_n235_), .C2(new_n223_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n215_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(G64gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(G57gat), .ZN(new_n242_));
  INV_X1    g041(.A(G57gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(G64gat), .ZN(new_n244_));
  AOI21_X1  g043(.A(KEYINPUT11), .B1(new_n242_), .B2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G71gat), .B(G78gat), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT69), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  AND2_X1   g046(.A1(G71gat), .A2(G78gat), .ZN(new_n248_));
  NOR2_X1   g047(.A1(G71gat), .A2(G78gat), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT69), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G57gat), .B(G64gat), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n250_), .B(new_n251_), .C1(new_n252_), .C2(KEYINPUT11), .ZN(new_n253_));
  AND2_X1   g052(.A1(new_n252_), .A2(KEYINPUT11), .ZN(new_n254_));
  AND3_X1   g053(.A1(new_n247_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n254_), .B1(new_n247_), .B2(new_n253_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n240_), .A2(new_n258_), .ZN(new_n259_));
  OAI211_X1 g058(.A(new_n257_), .B(new_n215_), .C1(new_n238_), .C2(new_n239_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n259_), .A2(KEYINPUT12), .A3(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT12), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n240_), .A2(new_n262_), .A3(new_n258_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n203_), .B1(new_n261_), .B2(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n202_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G120gat), .B(G148gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT5), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G176gat), .B(G204gat), .ZN(new_n269_));
  XOR2_X1   g068(.A(new_n268_), .B(new_n269_), .Z(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n266_), .A2(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n270_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n273_));
  AND3_X1   g072(.A1(new_n272_), .A2(KEYINPUT13), .A3(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(KEYINPUT13), .B1(new_n272_), .B2(new_n273_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n276_), .A2(KEYINPUT70), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(KEYINPUT70), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  XOR2_X1   g078(.A(G190gat), .B(G218gat), .Z(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT73), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G134gat), .B(G162gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT36), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  XOR2_X1   g084(.A(G29gat), .B(G36gat), .Z(new_n286_));
  XOR2_X1   g085(.A(G43gat), .B(G50gat), .Z(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT15), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT15), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n288_), .A2(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n240_), .A2(new_n290_), .A3(new_n292_), .ZN(new_n293_));
  AOI22_X1  g092(.A1(new_n209_), .A2(KEYINPUT67), .B1(new_n218_), .B2(new_n220_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n211_), .B1(new_n294_), .B2(new_n229_), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT68), .B1(new_n295_), .B2(new_n227_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n236_), .A2(new_n237_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n296_), .A2(new_n297_), .A3(new_n226_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n298_), .A2(new_n215_), .A3(new_n288_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT74), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G232gat), .A2(G233gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT72), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT35), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n300_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n293_), .A2(new_n299_), .A3(new_n306_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n304_), .A2(new_n305_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n308_), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n293_), .A2(new_n310_), .A3(new_n299_), .A4(new_n306_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n285_), .B1(new_n309_), .B2(new_n311_), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n283_), .A2(new_n284_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n309_), .A2(new_n313_), .A3(new_n311_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT75), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT75), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n309_), .A2(new_n316_), .A3(new_n313_), .A4(new_n311_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n312_), .B1(new_n315_), .B2(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n318_), .A2(KEYINPUT37), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT37), .ZN(new_n320_));
  AOI211_X1 g119(.A(new_n320_), .B(new_n312_), .C1(new_n315_), .C2(new_n317_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  XOR2_X1   g121(.A(KEYINPUT76), .B(G1gat), .Z(new_n323_));
  INV_X1    g122(.A(G8gat), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT14), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G15gat), .B(G22gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G1gat), .B(G8gat), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n325_), .A2(new_n326_), .A3(new_n328_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  XOR2_X1   g131(.A(KEYINPUT77), .B(KEYINPUT78), .Z(new_n333_));
  NAND2_X1  g132(.A1(G231gat), .A2(G233gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n332_), .B(new_n335_), .ZN(new_n336_));
  OR2_X1    g135(.A1(new_n336_), .A2(new_n257_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT79), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n336_), .A2(new_n257_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n337_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G127gat), .B(G155gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT16), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G183gat), .B(G211gat), .ZN(new_n343_));
  XOR2_X1   g142(.A(new_n342_), .B(new_n343_), .Z(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n340_), .A2(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n337_), .A2(new_n339_), .A3(new_n344_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT17), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n340_), .A2(KEYINPUT17), .A3(new_n345_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT80), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n349_), .A2(KEYINPUT80), .A3(new_n350_), .ZN(new_n354_));
  AND2_X1   g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n322_), .A2(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n279_), .A2(new_n356_), .ZN(new_n357_));
  OR2_X1    g156(.A1(new_n357_), .A2(KEYINPUT81), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(KEYINPUT81), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n290_), .A2(new_n331_), .A3(new_n292_), .A4(new_n330_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n332_), .A2(new_n288_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G229gat), .A2(G233gat), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n360_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n332_), .B(new_n289_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n363_), .B1(new_n364_), .B2(new_n362_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G113gat), .B(G141gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G169gat), .B(G197gat), .ZN(new_n367_));
  XOR2_X1   g166(.A(new_n366_), .B(new_n367_), .Z(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n365_), .A2(new_n369_), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n363_), .B(new_n368_), .C1(new_n364_), .C2(new_n362_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n370_), .A2(KEYINPUT82), .A3(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT82), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n365_), .A2(new_n373_), .A3(new_n369_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n372_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT2), .ZN(new_n376_));
  INV_X1    g175(.A(G141gat), .ZN(new_n377_));
  INV_X1    g176(.A(G148gat), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n376_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT3), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n380_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n382_));
  OAI21_X1  g181(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n379_), .A2(new_n381_), .A3(new_n382_), .A4(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(G155gat), .ZN(new_n385_));
  INV_X1    g184(.A(G162gat), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(G155gat), .A2(G162gat), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n384_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT87), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n384_), .A2(KEYINPUT87), .A3(new_n389_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT1), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n388_), .B1(new_n387_), .B2(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n395_), .B1(new_n394_), .B2(new_n387_), .ZN(new_n396_));
  XOR2_X1   g195(.A(G141gat), .B(G148gat), .Z(new_n397_));
  AOI22_X1  g196(.A1(new_n392_), .A2(new_n393_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G127gat), .B(G134gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT85), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G113gat), .B(G120gat), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  OR2_X1    g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n401_), .A2(new_n403_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n399_), .A2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n398_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n408_));
  AND2_X1   g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G225gat), .A2(G233gat), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n407_), .A2(KEYINPUT4), .A3(new_n408_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT4), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n399_), .A2(new_n414_), .A3(new_n406_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n410_), .B1(new_n413_), .B2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G57gat), .B(G85gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n417_), .B(new_n418_), .ZN(new_n419_));
  XOR2_X1   g218(.A(G1gat), .B(G29gat), .Z(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT96), .B(KEYINPUT97), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  OR3_X1    g222(.A1(new_n412_), .A2(new_n416_), .A3(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n423_), .B1(new_n412_), .B2(new_n416_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G71gat), .B(G99gat), .ZN(new_n427_));
  INV_X1    g226(.A(G43gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n427_), .B(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(KEYINPUT30), .ZN(new_n430_));
  NAND2_X1  g229(.A1(G227gat), .A2(G233gat), .ZN(new_n431_));
  INV_X1    g230(.A(G15gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n431_), .B(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n430_), .B(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(KEYINPUT25), .B(G183gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT26), .B(G190gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(KEYINPUT83), .ZN(new_n438_));
  INV_X1    g237(.A(G183gat), .ZN(new_n439_));
  INV_X1    g238(.A(G190gat), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT23), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT23), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n443_), .A2(G183gat), .A3(G190gat), .ZN(new_n444_));
  OR2_X1    g243(.A1(new_n444_), .A2(KEYINPUT84), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(KEYINPUT84), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n442_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(G169gat), .ZN(new_n448_));
  INV_X1    g247(.A(G176gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G169gat), .A2(G176gat), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n450_), .A2(KEYINPUT24), .A3(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n452_), .B1(KEYINPUT24), .B2(new_n450_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n447_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n438_), .A2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(KEYINPUT22), .B(G169gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(new_n449_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(new_n451_), .ZN(new_n458_));
  AND2_X1   g257(.A1(new_n441_), .A2(new_n444_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(G183gat), .A2(G190gat), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n455_), .B1(new_n458_), .B2(new_n461_), .ZN(new_n462_));
  OR2_X1    g261(.A1(new_n434_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n434_), .A2(new_n462_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n463_), .A2(KEYINPUT86), .A3(new_n464_), .ZN(new_n465_));
  XOR2_X1   g264(.A(new_n406_), .B(KEYINPUT31), .Z(new_n466_));
  XOR2_X1   g265(.A(new_n465_), .B(new_n466_), .Z(new_n467_));
  INV_X1    g266(.A(G50gat), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT29), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n398_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT28), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(G22gat), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n398_), .A2(KEYINPUT28), .A3(new_n469_), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n472_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n473_), .B1(new_n472_), .B2(new_n474_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n468_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n472_), .A2(new_n474_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(G22gat), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n472_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n479_), .A2(G50gat), .A3(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G78gat), .B(G106gat), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G228gat), .A2(G233gat), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n398_), .A2(new_n469_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G211gat), .B(G218gat), .ZN(new_n487_));
  XOR2_X1   g286(.A(G197gat), .B(G204gat), .Z(new_n488_));
  OAI21_X1  g287(.A(new_n487_), .B1(new_n488_), .B2(KEYINPUT88), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n489_), .A2(KEYINPUT21), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n488_), .A2(new_n487_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT21), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n490_), .B1(new_n489_), .B2(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n485_), .B1(new_n486_), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n493_), .A2(new_n489_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n496_), .B1(KEYINPUT21), .B2(new_n489_), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n497_), .B(new_n484_), .C1(new_n469_), .C2(new_n398_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n483_), .B1(new_n495_), .B2(new_n498_), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n477_), .B(new_n481_), .C1(KEYINPUT89), .C2(new_n499_), .ZN(new_n500_));
  AND3_X1   g299(.A1(new_n495_), .A2(new_n498_), .A3(new_n483_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n501_), .A2(new_n499_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n500_), .A2(new_n503_), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n499_), .A2(KEYINPUT89), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n505_), .A2(new_n502_), .A3(new_n477_), .A4(new_n481_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n467_), .A2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n465_), .B(new_n466_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n509_), .A2(new_n506_), .A3(new_n504_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n426_), .B1(new_n508_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT27), .ZN(new_n512_));
  INV_X1    g311(.A(new_n460_), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n445_), .A2(new_n446_), .ZN(new_n514_));
  OAI211_X1 g313(.A(KEYINPUT90), .B(new_n513_), .C1(new_n514_), .C2(new_n442_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT90), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n516_), .B1(new_n447_), .B2(new_n460_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n458_), .B1(new_n515_), .B2(new_n517_), .ZN(new_n518_));
  AOI211_X1 g317(.A(new_n459_), .B(new_n453_), .C1(new_n435_), .C2(new_n436_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n497_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT20), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n461_), .A2(new_n458_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n522_), .B1(new_n438_), .B2(new_n454_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n521_), .B1(new_n523_), .B2(new_n494_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n520_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G226gat), .A2(G233gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT19), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n525_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NOR3_X1   g329(.A1(new_n518_), .A2(new_n497_), .A3(new_n519_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT92), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n531_), .A2(new_n532_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n462_), .A2(KEYINPUT91), .A3(new_n497_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT91), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n536_), .B1(new_n523_), .B2(new_n494_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n535_), .A2(new_n537_), .A3(KEYINPUT20), .ZN(new_n538_));
  NOR3_X1   g337(.A1(new_n533_), .A2(new_n534_), .A3(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n530_), .B1(new_n539_), .B2(new_n527_), .ZN(new_n540_));
  XOR2_X1   g339(.A(G8gat), .B(G36gat), .Z(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT94), .ZN(new_n542_));
  XOR2_X1   g341(.A(G64gat), .B(G92gat), .Z(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n545_));
  XOR2_X1   g344(.A(new_n544_), .B(new_n545_), .Z(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n512_), .B1(new_n540_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT100), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n527_), .B1(new_n538_), .B2(new_n531_), .ZN(new_n550_));
  OAI21_X1  g349(.A(KEYINPUT98), .B1(new_n525_), .B2(new_n527_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT98), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n520_), .A2(new_n552_), .A3(new_n524_), .A4(new_n528_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n550_), .A2(new_n551_), .A3(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(KEYINPUT99), .B1(new_n554_), .B2(new_n546_), .ZN(new_n555_));
  AND3_X1   g354(.A1(new_n554_), .A2(KEYINPUT99), .A3(new_n546_), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n548_), .B(new_n549_), .C1(new_n555_), .C2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n540_), .A2(new_n547_), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n546_), .B(new_n530_), .C1(new_n539_), .C2(new_n527_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(new_n512_), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n558_), .B(KEYINPUT27), .C1(new_n556_), .C2(new_n555_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(KEYINPUT100), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n511_), .A2(new_n557_), .A3(new_n561_), .A4(new_n563_), .ZN(new_n564_));
  AND2_X1   g363(.A1(new_n547_), .A2(KEYINPUT32), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n554_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n540_), .ZN(new_n567_));
  OAI211_X1 g366(.A(new_n426_), .B(new_n566_), .C1(new_n567_), .C2(new_n565_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT33), .ZN(new_n569_));
  OR2_X1    g368(.A1(new_n425_), .A2(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n413_), .A2(new_n410_), .A3(new_n415_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n423_), .B1(new_n409_), .B2(new_n411_), .ZN(new_n572_));
  AOI22_X1  g371(.A1(new_n425_), .A2(new_n569_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n570_), .A2(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n568_), .B1(new_n560_), .B2(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n575_), .A2(new_n507_), .A3(new_n509_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n375_), .B1(new_n564_), .B2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n358_), .A2(new_n359_), .A3(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(KEYINPUT101), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT101), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n358_), .A2(new_n580_), .A3(new_n359_), .A4(new_n577_), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n426_), .A2(new_n323_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n582_), .A2(KEYINPUT38), .A3(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n351_), .ZN(new_n585_));
  NOR3_X1   g384(.A1(new_n279_), .A2(new_n585_), .A3(new_n375_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n318_), .B1(new_n564_), .B2(new_n576_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n586_), .A2(KEYINPUT102), .A3(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(KEYINPUT102), .B1(new_n586_), .B2(new_n587_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n426_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(G1gat), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n579_), .A2(new_n581_), .A3(new_n583_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT38), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n584_), .A2(new_n592_), .A3(new_n595_), .ZN(G1324gat));
  NAND2_X1  g395(.A1(new_n586_), .A2(new_n587_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n563_), .A2(new_n557_), .A3(new_n561_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  OAI21_X1  g398(.A(G8gat), .B1(new_n597_), .B2(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT39), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n579_), .A2(new_n324_), .A3(new_n598_), .A4(new_n581_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT40), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n601_), .A2(new_n602_), .A3(KEYINPUT40), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(G1325gat));
  INV_X1    g406(.A(KEYINPUT102), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n597_), .A2(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n509_), .B1(new_n609_), .B2(new_n588_), .ZN(new_n610_));
  OAI21_X1  g409(.A(KEYINPUT103), .B1(new_n610_), .B2(new_n432_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n467_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT103), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n612_), .A2(new_n613_), .A3(G15gat), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n611_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT41), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n582_), .A2(new_n432_), .A3(new_n467_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n611_), .A2(new_n614_), .A3(KEYINPUT41), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n617_), .A2(new_n618_), .A3(new_n619_), .ZN(G1326gat));
  INV_X1    g419(.A(new_n507_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n582_), .A2(new_n473_), .A3(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT42), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n621_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n623_), .B1(new_n624_), .B2(G22gat), .ZN(new_n625_));
  AND3_X1   g424(.A1(new_n624_), .A2(new_n623_), .A3(G22gat), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n622_), .B1(new_n625_), .B2(new_n626_), .ZN(G1327gat));
  NOR3_X1   g426(.A1(new_n279_), .A2(new_n355_), .A3(new_n375_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT104), .ZN(new_n629_));
  AOI221_X4 g428(.A(new_n322_), .B1(new_n629_), .B2(KEYINPUT43), .C1(new_n564_), .C2(new_n576_), .ZN(new_n630_));
  OAI21_X1  g429(.A(KEYINPUT43), .B1(new_n322_), .B2(new_n629_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n508_), .A2(new_n510_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n426_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n576_), .B1(new_n598_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n322_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n631_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n628_), .B1(new_n630_), .B2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT44), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n628_), .B(KEYINPUT44), .C1(new_n630_), .C2(new_n637_), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n640_), .A2(G29gat), .A3(new_n426_), .A4(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(G29gat), .ZN(new_n643_));
  INV_X1    g442(.A(new_n318_), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n279_), .A2(new_n644_), .A3(new_n355_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(new_n577_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n643_), .B1(new_n646_), .B2(new_n633_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n642_), .A2(new_n647_), .ZN(G1328gat));
  OR2_X1    g447(.A1(new_n599_), .A2(G36gat), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n646_), .A2(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT45), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n640_), .A2(new_n598_), .A3(new_n641_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(G36gat), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT46), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n651_), .A2(new_n653_), .A3(KEYINPUT46), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(G1329gat));
  NOR2_X1   g457(.A1(new_n509_), .A2(new_n428_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n640_), .A2(new_n641_), .A3(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT105), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n640_), .A2(KEYINPUT105), .A3(new_n641_), .A4(new_n659_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n428_), .B1(new_n646_), .B2(new_n509_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n662_), .A2(new_n663_), .A3(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(KEYINPUT47), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT47), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n662_), .A2(new_n667_), .A3(new_n663_), .A4(new_n664_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(G1330gat));
  NAND4_X1  g468(.A1(new_n640_), .A2(G50gat), .A3(new_n621_), .A4(new_n641_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n468_), .B1(new_n646_), .B2(new_n507_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n670_), .A2(new_n671_), .ZN(G1331gat));
  AND3_X1   g471(.A1(new_n353_), .A2(new_n354_), .A3(new_n375_), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n587_), .A2(new_n279_), .A3(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n674_), .A2(G57gat), .A3(new_n426_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT106), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n675_), .A2(new_n676_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n375_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n679_), .B1(new_n564_), .B2(new_n576_), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n680_), .A2(new_n279_), .A3(new_n322_), .A4(new_n355_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(G57gat), .B1(new_n682_), .B2(new_n426_), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n677_), .A2(new_n678_), .A3(new_n683_), .ZN(G1332gat));
  AOI21_X1  g483(.A(new_n241_), .B1(new_n674_), .B2(new_n598_), .ZN(new_n685_));
  XOR2_X1   g484(.A(new_n685_), .B(KEYINPUT48), .Z(new_n686_));
  NAND3_X1  g485(.A1(new_n682_), .A2(new_n241_), .A3(new_n598_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(G1333gat));
  INV_X1    g487(.A(G71gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n689_), .B1(new_n674_), .B2(new_n467_), .ZN(new_n690_));
  XOR2_X1   g489(.A(new_n690_), .B(KEYINPUT49), .Z(new_n691_));
  NAND3_X1  g490(.A1(new_n682_), .A2(new_n689_), .A3(new_n467_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(G1334gat));
  INV_X1    g492(.A(G78gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n694_), .B1(new_n674_), .B2(new_n621_), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT50), .Z(new_n696_));
  NAND3_X1  g495(.A1(new_n682_), .A2(new_n694_), .A3(new_n621_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(G1335gat));
  OR2_X1    g497(.A1(new_n630_), .A2(new_n637_), .ZN(new_n699_));
  AOI211_X1 g498(.A(new_n355_), .B(new_n679_), .C1(new_n277_), .C2(new_n278_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n426_), .A2(G85gat), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT108), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n699_), .A2(new_n700_), .A3(new_n702_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n355_), .A2(new_n644_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n680_), .A2(new_n279_), .A3(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(KEYINPUT107), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT107), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n680_), .A2(new_n707_), .A3(new_n279_), .A4(new_n704_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n633_), .B1(new_n706_), .B2(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n703_), .B1(new_n709_), .B2(G85gat), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT109), .Z(G1336gat));
  INV_X1    g510(.A(G92gat), .ZN(new_n712_));
  INV_X1    g511(.A(new_n706_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n708_), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n712_), .B(new_n598_), .C1(new_n713_), .C2(new_n714_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n699_), .A2(new_n598_), .A3(new_n700_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n715_), .B1(new_n717_), .B2(new_n712_), .ZN(G1337gat));
  XNOR2_X1  g517(.A(KEYINPUT111), .B(KEYINPUT51), .ZN(new_n719_));
  OAI211_X1 g518(.A(new_n467_), .B(new_n700_), .C1(new_n630_), .C2(new_n637_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(G99gat), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT110), .ZN(new_n722_));
  OAI211_X1 g521(.A(new_n204_), .B(new_n467_), .C1(new_n713_), .C2(new_n714_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n719_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n721_), .A2(KEYINPUT110), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT110), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n726_), .B1(new_n720_), .B2(G99gat), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n723_), .B(new_n719_), .C1(new_n725_), .C2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n724_), .A2(new_n729_), .ZN(G1338gat));
  OAI211_X1 g529(.A(new_n621_), .B(new_n700_), .C1(new_n630_), .C2(new_n637_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(G106gat), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT112), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n731_), .A2(KEYINPUT112), .A3(G106gat), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n734_), .A2(KEYINPUT52), .A3(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n621_), .A2(new_n205_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n737_), .B1(new_n706_), .B2(new_n708_), .ZN(new_n738_));
  AOI21_X1  g537(.A(KEYINPUT112), .B1(new_n731_), .B2(G106gat), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT52), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n738_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n742_));
  AND3_X1   g541(.A1(new_n736_), .A2(new_n741_), .A3(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n736_), .B2(new_n741_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n743_), .A2(new_n744_), .ZN(G1339gat));
  XNOR2_X1  g544(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n673_), .A2(new_n276_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n747_), .B1(new_n748_), .B2(new_n636_), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n673_), .A2(new_n322_), .A3(new_n276_), .A4(new_n746_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n362_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n369_), .B1(new_n364_), .B2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT116), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  OAI211_X1 g554(.A(KEYINPUT116), .B(new_n369_), .C1(new_n364_), .C2(new_n752_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n360_), .A2(new_n361_), .A3(new_n752_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n755_), .A2(new_n756_), .A3(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(new_n371_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(KEYINPUT117), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT117), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n758_), .A2(new_n761_), .A3(new_n371_), .ZN(new_n762_));
  AOI22_X1  g561(.A1(new_n760_), .A2(new_n762_), .B1(new_n273_), .B2(new_n272_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n261_), .A2(new_n203_), .A3(new_n263_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT55), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n261_), .A2(new_n263_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n765_), .B1(new_n766_), .B2(new_n202_), .ZN(new_n767_));
  AOI211_X1 g566(.A(KEYINPUT55), .B(new_n203_), .C1(new_n261_), .C2(new_n263_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n764_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n769_), .A2(KEYINPUT115), .A3(KEYINPUT56), .A4(new_n270_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n375_), .B1(new_n266_), .B2(new_n271_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT56), .ZN(new_n773_));
  INV_X1    g572(.A(new_n764_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n260_), .A2(KEYINPUT12), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n257_), .B1(new_n298_), .B2(new_n215_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n263_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n202_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT55), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n264_), .A2(new_n765_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n774_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n773_), .B1(new_n782_), .B2(new_n271_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT115), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n769_), .A2(KEYINPUT56), .A3(new_n270_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n783_), .A2(new_n784_), .A3(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n763_), .B1(new_n772_), .B2(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(KEYINPUT57), .B1(new_n787_), .B2(new_n318_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT57), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n770_), .A2(new_n771_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n780_), .A2(new_n781_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n271_), .B1(new_n791_), .B2(new_n764_), .ZN(new_n792_));
  AOI21_X1  g591(.A(KEYINPUT115), .B1(new_n792_), .B2(KEYINPUT56), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n790_), .B1(new_n793_), .B2(new_n783_), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n789_), .B(new_n644_), .C1(new_n794_), .C2(new_n763_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT118), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n796_), .B(new_n773_), .C1(new_n782_), .C2(new_n271_), .ZN(new_n797_));
  AOI22_X1  g596(.A1(new_n760_), .A2(new_n762_), .B1(new_n266_), .B2(new_n271_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n785_), .A2(KEYINPUT118), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT56), .B1(new_n769_), .B2(new_n270_), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n797_), .B(new_n798_), .C1(new_n799_), .C2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT58), .ZN(new_n802_));
  OR2_X1    g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n322_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n804_));
  AOI22_X1  g603(.A1(new_n788_), .A2(new_n795_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n751_), .B1(new_n805_), .B2(new_n355_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT59), .ZN(new_n807_));
  NOR3_X1   g606(.A1(new_n598_), .A2(new_n633_), .A3(new_n508_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n806_), .A2(new_n807_), .A3(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT120), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n751_), .B1(new_n805_), .B2(new_n351_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n808_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n810_), .B1(new_n812_), .B2(KEYINPUT59), .ZN(new_n813_));
  AOI211_X1 g612(.A(KEYINPUT120), .B(new_n807_), .C1(new_n811_), .C2(new_n808_), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n679_), .B(new_n809_), .C1(new_n813_), .C2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(G113gat), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT119), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n812_), .B(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(G113gat), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n818_), .A2(new_n819_), .A3(new_n679_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n816_), .A2(new_n820_), .ZN(G1340gat));
  OAI211_X1 g620(.A(new_n279_), .B(new_n809_), .C1(new_n813_), .C2(new_n814_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(G120gat), .ZN(new_n823_));
  INV_X1    g622(.A(G120gat), .ZN(new_n824_));
  OR2_X1    g623(.A1(new_n824_), .A2(KEYINPUT60), .ZN(new_n825_));
  INV_X1    g624(.A(new_n279_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n824_), .B1(new_n826_), .B2(KEYINPUT60), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n818_), .A2(new_n825_), .A3(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n823_), .A2(new_n828_), .ZN(G1341gat));
  OAI211_X1 g628(.A(new_n351_), .B(new_n809_), .C1(new_n813_), .C2(new_n814_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(G127gat), .ZN(new_n831_));
  INV_X1    g630(.A(G127gat), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n818_), .A2(new_n832_), .A3(new_n355_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(G1342gat));
  OAI211_X1 g633(.A(new_n636_), .B(new_n809_), .C1(new_n813_), .C2(new_n814_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(G134gat), .ZN(new_n836_));
  INV_X1    g635(.A(G134gat), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n818_), .A2(new_n837_), .A3(new_n318_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n838_), .ZN(G1343gat));
  INV_X1    g638(.A(new_n510_), .ZN(new_n840_));
  AND2_X1   g639(.A1(new_n811_), .A2(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n598_), .A2(new_n633_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n844_), .A2(new_n377_), .A3(new_n679_), .ZN(new_n845_));
  OAI21_X1  g644(.A(G141gat), .B1(new_n843_), .B2(new_n375_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(G1344gat));
  NAND3_X1  g646(.A1(new_n844_), .A2(new_n378_), .A3(new_n279_), .ZN(new_n848_));
  OAI21_X1  g647(.A(G148gat), .B1(new_n843_), .B2(new_n826_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(G1345gat));
  NAND4_X1  g649(.A1(new_n811_), .A2(new_n355_), .A3(new_n840_), .A4(new_n842_), .ZN(new_n851_));
  OR2_X1    g650(.A1(new_n851_), .A2(KEYINPUT121), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(KEYINPUT121), .ZN(new_n853_));
  XNOR2_X1  g652(.A(KEYINPUT61), .B(G155gat), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n852_), .A2(new_n853_), .A3(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n854_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n855_), .A2(new_n856_), .ZN(G1346gat));
  OAI21_X1  g656(.A(G162gat), .B1(new_n843_), .B2(new_n322_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n318_), .A2(new_n386_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n843_), .B2(new_n859_), .ZN(G1347gat));
  NOR2_X1   g659(.A1(new_n599_), .A2(new_n426_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n467_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n862_), .A2(new_n621_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n806_), .A2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n679_), .A2(new_n456_), .ZN(new_n865_));
  XOR2_X1   g664(.A(new_n865_), .B(KEYINPUT123), .Z(new_n866_));
  NOR2_X1   g665(.A1(new_n864_), .A2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT122), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n448_), .B1(new_n868_), .B2(KEYINPUT62), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n869_), .B1(new_n864_), .B2(new_n375_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n868_), .A2(KEYINPUT62), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n867_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n872_), .B1(new_n870_), .B2(new_n871_), .ZN(G1348gat));
  INV_X1    g672(.A(new_n864_), .ZN(new_n874_));
  AOI21_X1  g673(.A(G176gat), .B1(new_n874_), .B2(new_n279_), .ZN(new_n875_));
  AND2_X1   g674(.A1(new_n811_), .A2(new_n507_), .ZN(new_n876_));
  NOR3_X1   g675(.A1(new_n862_), .A2(new_n826_), .A3(new_n449_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n875_), .B1(new_n876_), .B2(new_n877_), .ZN(G1349gat));
  NOR3_X1   g677(.A1(new_n864_), .A2(new_n585_), .A3(new_n435_), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n876_), .A2(new_n355_), .A3(new_n467_), .A4(new_n861_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n879_), .B1(new_n880_), .B2(new_n439_), .ZN(G1350gat));
  OAI21_X1  g680(.A(G190gat), .B1(new_n864_), .B2(new_n322_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n318_), .A2(new_n436_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(KEYINPUT124), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n882_), .B1(new_n864_), .B2(new_n884_), .ZN(G1351gat));
  NAND3_X1  g684(.A1(new_n841_), .A2(new_n679_), .A3(new_n861_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(G197gat), .ZN(G1352gat));
  AND3_X1   g686(.A1(new_n841_), .A2(new_n279_), .A3(new_n861_), .ZN(new_n888_));
  INV_X1    g687(.A(G204gat), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n888_), .B(new_n889_), .ZN(G1353gat));
  AOI21_X1  g689(.A(new_n585_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n811_), .A2(new_n840_), .A3(new_n861_), .A4(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(KEYINPUT125), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n892_), .A2(KEYINPUT125), .ZN(new_n895_));
  OAI22_X1  g694(.A1(new_n894_), .A2(new_n895_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n896_));
  INV_X1    g695(.A(new_n895_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n897_), .A2(new_n898_), .A3(new_n893_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n896_), .A2(new_n899_), .ZN(G1354gat));
  NAND3_X1  g699(.A1(new_n841_), .A2(new_n318_), .A3(new_n861_), .ZN(new_n901_));
  OR2_X1    g700(.A1(new_n901_), .A2(KEYINPUT126), .ZN(new_n902_));
  AOI21_X1  g701(.A(G218gat), .B1(new_n901_), .B2(KEYINPUT126), .ZN(new_n903_));
  AND2_X1   g702(.A1(new_n841_), .A2(new_n861_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n636_), .A2(G218gat), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(KEYINPUT127), .ZN(new_n906_));
  AOI22_X1  g705(.A1(new_n902_), .A2(new_n903_), .B1(new_n904_), .B2(new_n906_), .ZN(G1355gat));
endmodule


