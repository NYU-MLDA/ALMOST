//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 1 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 0 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 1 1 1 0 0 0 1 0 1 1 0 0 0 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n753_, new_n754_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n800_, new_n801_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n907_, new_n909_, new_n910_, new_n912_, new_n913_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n930_, new_n931_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n939_, new_n940_, new_n941_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n952_, new_n953_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n961_, new_n962_;
  XNOR2_X1  g000(.A(G176gat), .B(G204gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G120gat), .B(G148gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT6), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT6), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n209_), .A2(G99gat), .A3(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G85gat), .A2(G92gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT9), .ZN(new_n213_));
  AOI22_X1  g012(.A1(new_n208_), .A2(new_n210_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(G106gat), .ZN(new_n215_));
  INV_X1    g014(.A(G99gat), .ZN(new_n216_));
  AND2_X1   g015(.A1(new_n216_), .A2(KEYINPUT10), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n216_), .A2(KEYINPUT10), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n215_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G85gat), .A2(G92gat), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(KEYINPUT9), .A3(new_n211_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n214_), .A2(new_n219_), .A3(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n208_), .A2(new_n210_), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT7), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n226_), .A2(new_n216_), .A3(new_n215_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n224_), .A2(new_n225_), .A3(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT8), .ZN(new_n229_));
  NOR3_X1   g028(.A1(new_n212_), .A2(new_n220_), .A3(KEYINPUT66), .ZN(new_n230_));
  AND3_X1   g029(.A1(new_n228_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n229_), .B1(new_n228_), .B2(new_n230_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n223_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(G71gat), .B(G78gat), .Z(new_n234_));
  INV_X1    g033(.A(G57gat), .ZN(new_n235_));
  INV_X1    g034(.A(G64gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT11), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G57gat), .A2(G64gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n237_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n234_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n237_), .A2(new_n239_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n242_), .B1(new_n243_), .B2(KEYINPUT11), .ZN(new_n244_));
  AND2_X1   g043(.A1(G57gat), .A2(G64gat), .ZN(new_n245_));
  NOR2_X1   g044(.A1(G57gat), .A2(G64gat), .ZN(new_n246_));
  OAI211_X1 g045(.A(new_n242_), .B(KEYINPUT11), .C1(new_n245_), .C2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n241_), .B1(new_n244_), .B2(new_n248_), .ZN(new_n249_));
  OAI21_X1  g048(.A(KEYINPUT11), .B1(new_n245_), .B2(new_n246_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT67), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n251_), .A2(new_n240_), .A3(new_n234_), .A4(new_n247_), .ZN(new_n252_));
  AND2_X1   g051(.A1(new_n249_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n233_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT68), .ZN(new_n255_));
  AND2_X1   g054(.A1(new_n208_), .A2(new_n210_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n227_), .A2(new_n225_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n230_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT8), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n228_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n249_), .A2(new_n252_), .ZN(new_n262_));
  AND4_X1   g061(.A1(new_n255_), .A2(new_n261_), .A3(new_n223_), .A4(new_n262_), .ZN(new_n263_));
  AND3_X1   g062(.A1(new_n214_), .A2(new_n219_), .A3(new_n222_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n264_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n255_), .B1(new_n265_), .B2(new_n262_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n254_), .B1(new_n263_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G230gat), .A2(G233gat), .ZN(new_n268_));
  XOR2_X1   g067(.A(new_n268_), .B(KEYINPUT64), .Z(new_n269_));
  XOR2_X1   g068(.A(new_n269_), .B(KEYINPUT65), .Z(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n267_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT12), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n273_), .B1(new_n265_), .B2(new_n262_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n233_), .A2(new_n253_), .A3(KEYINPUT12), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n265_), .A2(new_n262_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n274_), .A2(new_n275_), .A3(new_n276_), .A4(new_n270_), .ZN(new_n277_));
  AOI21_X1  g076(.A(KEYINPUT69), .B1(new_n272_), .B2(new_n277_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n265_), .A2(new_n262_), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT68), .B1(new_n233_), .B2(new_n253_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n265_), .A2(new_n255_), .A3(new_n262_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n279_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  OAI211_X1 g081(.A(KEYINPUT69), .B(new_n277_), .C1(new_n282_), .C2(new_n270_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n206_), .B1(new_n278_), .B2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(KEYINPUT71), .ZN(new_n286_));
  INV_X1    g085(.A(new_n206_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n272_), .A2(new_n277_), .A3(new_n287_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n277_), .B1(new_n282_), .B2(new_n270_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT69), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(new_n283_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT71), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n292_), .A2(new_n293_), .A3(new_n206_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n286_), .A2(new_n288_), .A3(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(KEYINPUT13), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT13), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n286_), .A2(new_n297_), .A3(new_n288_), .A4(new_n294_), .ZN(new_n298_));
  AND3_X1   g097(.A1(new_n296_), .A2(KEYINPUT72), .A3(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(KEYINPUT72), .B1(new_n296_), .B2(new_n298_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(G50gat), .ZN(new_n302_));
  OR2_X1    g101(.A1(G29gat), .A2(G36gat), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT73), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G29gat), .A2(G36gat), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n303_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n304_), .B1(new_n303_), .B2(new_n305_), .ZN(new_n308_));
  NOR3_X1   g107(.A1(new_n307_), .A2(G43gat), .A3(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(G43gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n303_), .A2(new_n305_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(KEYINPUT73), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n310_), .B1(new_n312_), .B2(new_n306_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n302_), .B1(new_n309_), .B2(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(G43gat), .B1(new_n307_), .B2(new_n308_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n312_), .A2(new_n310_), .A3(new_n306_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n315_), .A2(G50gat), .A3(new_n316_), .ZN(new_n317_));
  AND2_X1   g116(.A1(new_n314_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(G1gat), .ZN(new_n319_));
  INV_X1    g118(.A(G8gat), .ZN(new_n320_));
  OAI21_X1  g119(.A(KEYINPUT14), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT76), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G15gat), .B(G22gat), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT76), .ZN(new_n324_));
  OAI211_X1 g123(.A(new_n324_), .B(KEYINPUT14), .C1(new_n319_), .C2(new_n320_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n322_), .A2(new_n323_), .A3(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G1gat), .B(G8gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  AND2_X1   g127(.A1(new_n318_), .A2(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n318_), .A2(new_n328_), .ZN(new_n330_));
  OAI211_X1 g129(.A(G229gat), .B(G233gat), .C1(new_n329_), .C2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n330_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G229gat), .A2(G233gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n314_), .A2(new_n317_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT15), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n314_), .A2(KEYINPUT15), .A3(new_n317_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n336_), .A2(new_n328_), .A3(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n332_), .A2(new_n333_), .A3(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n331_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G113gat), .B(G141gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT80), .ZN(new_n342_));
  INV_X1    g141(.A(G169gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(G197gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n340_), .A2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n331_), .A2(new_n339_), .A3(new_n346_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n301_), .A2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G1gat), .B(G29gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(G85gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT0), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(new_n235_), .ZN(new_n355_));
  INV_X1    g154(.A(G141gat), .ZN(new_n356_));
  INV_X1    g155(.A(G148gat), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n356_), .A2(new_n357_), .A3(KEYINPUT89), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(KEYINPUT3), .ZN(new_n359_));
  NAND3_X1  g158(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT3), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n361_), .A2(new_n356_), .A3(new_n357_), .A4(KEYINPUT89), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT2), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n363_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n359_), .A2(new_n360_), .A3(new_n362_), .A4(new_n364_), .ZN(new_n365_));
  OR2_X1    g164(.A1(G155gat), .A2(G162gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G155gat), .A2(G162gat), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n365_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT88), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n367_), .A2(KEYINPUT1), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT1), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n372_), .A2(G155gat), .A3(G162gat), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n371_), .A2(new_n373_), .A3(new_n366_), .ZN(new_n374_));
  XOR2_X1   g173(.A(G141gat), .B(G148gat), .Z(new_n375_));
  AOI21_X1  g174(.A(new_n370_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  AND3_X1   g175(.A1(new_n374_), .A2(new_n375_), .A3(new_n370_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n369_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G127gat), .A2(G134gat), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(G127gat), .A2(G134gat), .ZN(new_n381_));
  OAI21_X1  g180(.A(G113gat), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(G127gat), .ZN(new_n383_));
  INV_X1    g182(.A(G134gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(G113gat), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(new_n386_), .A3(new_n379_), .ZN(new_n387_));
  AND3_X1   g186(.A1(new_n382_), .A2(new_n387_), .A3(G120gat), .ZN(new_n388_));
  AOI21_X1  g187(.A(G120gat), .B1(new_n382_), .B2(new_n387_), .ZN(new_n389_));
  OR2_X1    g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n378_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n374_), .A2(new_n375_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(KEYINPUT88), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n374_), .A2(new_n375_), .A3(new_n370_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n388_), .A2(new_n389_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n395_), .A2(new_n396_), .A3(new_n369_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n391_), .A2(KEYINPUT95), .A3(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT95), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n378_), .A2(new_n390_), .A3(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n398_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT4), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G225gat), .A2(G233gat), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n391_), .A2(KEYINPUT4), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n402_), .A2(new_n404_), .A3(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT96), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n408_), .B1(new_n401_), .B2(new_n403_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n407_), .A2(new_n410_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n402_), .A2(KEYINPUT96), .A3(new_n404_), .A4(new_n406_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n355_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT4), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n415_), .B1(new_n398_), .B2(new_n400_), .ZN(new_n416_));
  NOR3_X1   g215(.A1(new_n416_), .A2(new_n403_), .A3(new_n405_), .ZN(new_n417_));
  OAI211_X1 g216(.A(new_n412_), .B(new_n355_), .C1(new_n417_), .C2(new_n409_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n414_), .A2(new_n418_), .ZN(new_n419_));
  XOR2_X1   g218(.A(G78gat), .B(G106gat), .Z(new_n420_));
  XNOR2_X1  g219(.A(G22gat), .B(G50gat), .ZN(new_n421_));
  NOR3_X1   g220(.A1(new_n378_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT28), .ZN(new_n423_));
  AOI22_X1  g222(.A1(new_n393_), .A2(new_n394_), .B1(new_n368_), .B2(new_n365_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT29), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n423_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n421_), .B1(new_n422_), .B2(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT28), .B1(new_n378_), .B2(KEYINPUT29), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n424_), .A2(new_n423_), .A3(new_n425_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n421_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n428_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n427_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT94), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT21), .ZN(new_n434_));
  INV_X1    g233(.A(G204gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(G197gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n345_), .A2(G204gat), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n434_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  AND2_X1   g237(.A1(G211gat), .A2(G218gat), .ZN(new_n439_));
  NOR2_X1   g238(.A1(G211gat), .A2(G218gat), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT90), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(G211gat), .ZN(new_n442_));
  INV_X1    g241(.A(G218gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT90), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G211gat), .A2(G218gat), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n444_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n438_), .A2(new_n441_), .A3(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT92), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT92), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n438_), .A2(new_n441_), .A3(new_n447_), .A4(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n449_), .A2(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n345_), .A2(G204gat), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n435_), .A2(G197gat), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT21), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n436_), .A2(new_n437_), .A3(new_n434_), .ZN(new_n456_));
  NOR3_X1   g255(.A1(new_n439_), .A2(new_n440_), .A3(KEYINPUT90), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n445_), .B1(new_n444_), .B2(new_n446_), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n455_), .B(new_n456_), .C1(new_n457_), .C2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT91), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G197gat), .B(G204gat), .ZN(new_n462_));
  AOI22_X1  g261(.A1(new_n441_), .A2(new_n447_), .B1(new_n462_), .B2(new_n434_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n463_), .A2(KEYINPUT91), .A3(new_n455_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n452_), .B1(new_n461_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G228gat), .A2(G233gat), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n425_), .B1(new_n395_), .B2(new_n369_), .ZN(new_n468_));
  NOR3_X1   g267(.A1(new_n465_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n461_), .A2(new_n464_), .ZN(new_n470_));
  AND2_X1   g269(.A1(new_n449_), .A2(new_n451_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT93), .B(KEYINPUT29), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n378_), .A2(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n466_), .B1(new_n472_), .B2(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n433_), .B1(new_n469_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n473_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n477_), .B1(new_n395_), .B2(new_n369_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n467_), .B1(new_n465_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n378_), .A2(KEYINPUT29), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n472_), .A2(new_n466_), .A3(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n479_), .A2(KEYINPUT94), .A3(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n432_), .B1(new_n476_), .B2(new_n482_), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n432_), .A2(new_n482_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n420_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  AND2_X1   g284(.A1(new_n427_), .A2(new_n431_), .ZN(new_n486_));
  AND3_X1   g285(.A1(new_n479_), .A2(KEYINPUT94), .A3(new_n481_), .ZN(new_n487_));
  AOI21_X1  g286(.A(KEYINPUT94), .B1(new_n479_), .B2(new_n481_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n486_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n420_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n432_), .A2(new_n482_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n489_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT83), .ZN(new_n493_));
  INV_X1    g292(.A(G176gat), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n493_), .A2(new_n343_), .A3(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G169gat), .A2(G176gat), .ZN(new_n496_));
  OAI21_X1  g295(.A(KEYINPUT83), .B1(G169gat), .B2(G176gat), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n495_), .A2(KEYINPUT24), .A3(new_n496_), .A4(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(KEYINPUT82), .A2(G183gat), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT81), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n499_), .A2(new_n500_), .A3(KEYINPUT25), .ZN(new_n501_));
  NOR2_X1   g300(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n502_));
  AND2_X1   g301(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n501_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT25), .ZN(new_n505_));
  OAI21_X1  g304(.A(KEYINPUT81), .B1(new_n505_), .B2(G183gat), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n505_), .A2(KEYINPUT82), .A3(G183gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n498_), .B1(new_n504_), .B2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT84), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G183gat), .A2(G190gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(KEYINPUT23), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT23), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n514_), .A2(G183gat), .A3(G190gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  OAI211_X1 g315(.A(KEYINPUT84), .B(new_n498_), .C1(new_n504_), .C2(new_n508_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT24), .ZN(new_n518_));
  INV_X1    g317(.A(new_n497_), .ZN(new_n519_));
  NOR3_X1   g318(.A1(KEYINPUT83), .A2(G169gat), .A3(G176gat), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n518_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n511_), .A2(new_n516_), .A3(new_n517_), .A4(new_n521_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(new_n343_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n513_), .A2(new_n515_), .A3(KEYINPUT85), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT85), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n512_), .A2(new_n527_), .A3(KEYINPUT23), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n526_), .A2(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(G183gat), .A2(G190gat), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n525_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n522_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(G99gat), .ZN(new_n533_));
  INV_X1    g332(.A(new_n531_), .ZN(new_n534_));
  AND2_X1   g333(.A1(new_n517_), .A2(new_n521_), .ZN(new_n535_));
  AOI22_X1  g334(.A1(new_n509_), .A2(new_n510_), .B1(new_n513_), .B2(new_n515_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n534_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(new_n216_), .ZN(new_n538_));
  XOR2_X1   g337(.A(G15gat), .B(G43gat), .Z(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT86), .ZN(new_n540_));
  XOR2_X1   g339(.A(KEYINPUT30), .B(G71gat), .Z(new_n541_));
  NAND2_X1  g340(.A1(G227gat), .A2(G233gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n540_), .B(new_n543_), .ZN(new_n544_));
  AND3_X1   g343(.A1(new_n533_), .A2(new_n538_), .A3(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n544_), .B1(new_n533_), .B2(new_n538_), .ZN(new_n546_));
  OAI21_X1  g345(.A(KEYINPUT87), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n544_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n532_), .A2(G99gat), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n537_), .A2(new_n216_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n548_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT87), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n533_), .A2(new_n538_), .A3(new_n544_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n551_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n396_), .B(KEYINPUT31), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n547_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n555_), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n551_), .A2(new_n552_), .A3(new_n553_), .A4(new_n557_), .ZN(new_n558_));
  AND4_X1   g357(.A1(new_n485_), .A2(new_n492_), .A3(new_n556_), .A4(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT99), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G8gat), .B(G36gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT18), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(G64gat), .ZN(new_n563_));
  INV_X1    g362(.A(G92gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n530_), .B1(new_n513_), .B2(new_n515_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n524_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(KEYINPUT26), .B(G190gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(KEYINPUT25), .B(G183gat), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  AND3_X1   g370(.A1(new_n521_), .A2(new_n571_), .A3(new_n498_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n529_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n568_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n470_), .A2(new_n574_), .A3(new_n471_), .ZN(new_n575_));
  OAI211_X1 g374(.A(new_n575_), .B(KEYINPUT20), .C1(new_n537_), .C2(new_n465_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G226gat), .A2(G233gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT19), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n576_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT20), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n581_), .B1(new_n537_), .B2(new_n465_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n521_), .A2(new_n571_), .A3(new_n498_), .ZN(new_n583_));
  OAI22_X1  g382(.A1(new_n583_), .A2(new_n529_), .B1(new_n524_), .B2(new_n567_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n459_), .A2(new_n460_), .ZN(new_n585_));
  AOI21_X1  g384(.A(KEYINPUT91), .B1(new_n463_), .B2(new_n455_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n584_), .B1(new_n587_), .B2(new_n452_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n582_), .A2(new_n578_), .A3(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n566_), .B1(new_n580_), .B2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n576_), .A2(new_n578_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n582_), .A2(new_n579_), .A3(new_n588_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n565_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT27), .ZN(new_n594_));
  NOR3_X1   g393(.A1(new_n590_), .A2(new_n593_), .A3(new_n594_), .ZN(new_n595_));
  XOR2_X1   g394(.A(KEYINPUT98), .B(KEYINPUT27), .Z(new_n596_));
  AOI21_X1  g395(.A(new_n581_), .B1(new_n532_), .B2(new_n472_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n578_), .B1(new_n597_), .B2(new_n575_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n522_), .A2(new_n470_), .A3(new_n471_), .A4(new_n531_), .ZN(new_n599_));
  AND4_X1   g398(.A1(KEYINPUT20), .A2(new_n588_), .A3(new_n578_), .A4(new_n599_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n565_), .B1(new_n598_), .B2(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n580_), .A2(new_n589_), .A3(new_n566_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n596_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n560_), .B1(new_n595_), .B2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n593_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n605_), .A2(new_n601_), .A3(KEYINPUT27), .ZN(new_n606_));
  INV_X1    g405(.A(new_n596_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n602_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n607_), .B1(new_n608_), .B2(new_n590_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n606_), .A2(new_n609_), .A3(KEYINPUT99), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n559_), .A2(new_n604_), .A3(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n485_), .A2(new_n492_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n556_), .A2(new_n558_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n612_), .A2(new_n613_), .A3(new_n609_), .A4(new_n606_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n419_), .B1(new_n611_), .B2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n612_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(new_n613_), .ZN(new_n617_));
  NOR4_X1   g416(.A1(new_n416_), .A2(new_n408_), .A3(new_n403_), .A4(new_n405_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n618_), .B1(new_n407_), .B2(new_n410_), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n619_), .A2(KEYINPUT97), .A3(KEYINPUT33), .A4(new_n355_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT97), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT33), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n621_), .B1(new_n418_), .B2(new_n622_), .ZN(new_n623_));
  NOR3_X1   g422(.A1(new_n416_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n403_), .B1(new_n398_), .B2(new_n400_), .ZN(new_n625_));
  NOR3_X1   g424(.A1(new_n624_), .A2(new_n355_), .A3(new_n625_), .ZN(new_n626_));
  NOR3_X1   g425(.A1(new_n626_), .A2(new_n590_), .A3(new_n608_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n418_), .A2(new_n622_), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n620_), .A2(new_n623_), .A3(new_n627_), .A4(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n565_), .A2(KEYINPUT32), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n630_), .B1(new_n598_), .B2(new_n600_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n591_), .A2(new_n592_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n632_), .A2(KEYINPUT32), .A3(new_n565_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n418_), .ZN(new_n634_));
  OAI211_X1 g433(.A(new_n631_), .B(new_n633_), .C1(new_n634_), .C2(new_n413_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n617_), .B1(new_n629_), .B2(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n615_), .A2(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n351_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(G231gat), .A2(G233gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n328_), .B(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(new_n262_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(G183gat), .B(G211gat), .ZN(new_n642_));
  XNOR2_X1  g441(.A(G127gat), .B(G155gat), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n642_), .B(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n644_), .B(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT78), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n641_), .A2(new_n647_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n648_), .B1(new_n641_), .B2(new_n646_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(KEYINPUT17), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT17), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n648_), .A2(new_n651_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n650_), .A2(new_n652_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n336_), .A2(new_n337_), .A3(new_n233_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(KEYINPUT74), .ZN(new_n655_));
  NAND2_X1  g454(.A1(G232gat), .A2(G233gat), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT34), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n655_), .A2(KEYINPUT35), .A3(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n334_), .A2(new_n265_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n654_), .A2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n654_), .A2(new_n659_), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n662_), .A2(KEYINPUT35), .A3(new_n657_), .A4(new_n655_), .ZN(new_n663_));
  OR2_X1    g462(.A1(new_n657_), .A2(KEYINPUT35), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n661_), .A2(new_n663_), .A3(new_n664_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(G190gat), .B(G218gat), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(G134gat), .ZN(new_n667_));
  INV_X1    g466(.A(G162gat), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n667_), .B(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n670_), .A2(KEYINPUT36), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n665_), .A2(new_n671_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n669_), .B(KEYINPUT36), .ZN(new_n673_));
  NAND4_X1  g472(.A1(new_n661_), .A2(new_n663_), .A3(new_n664_), .A4(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n672_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT37), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT75), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n676_), .B1(new_n674_), .B2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n675_), .A2(new_n678_), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n672_), .B(new_n674_), .C1(new_n677_), .C2(new_n676_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n653_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT79), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n638_), .A2(new_n682_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n683_), .A2(new_n319_), .A3(new_n419_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT38), .ZN(new_n685_));
  INV_X1    g484(.A(new_n675_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n686_), .A2(new_n653_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n638_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n419_), .ZN(new_n689_));
  OAI21_X1  g488(.A(G1gat), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n685_), .A2(new_n690_), .ZN(G1324gat));
  INV_X1    g490(.A(KEYINPUT100), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n604_), .A2(new_n610_), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n638_), .A2(new_n693_), .A3(new_n687_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n692_), .B1(new_n694_), .B2(new_n320_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n693_), .ZN(new_n696_));
  OAI211_X1 g495(.A(KEYINPUT100), .B(G8gat), .C1(new_n688_), .C2(new_n696_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n695_), .A2(new_n697_), .A3(KEYINPUT39), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n683_), .A2(new_n320_), .A3(new_n693_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT39), .ZN(new_n700_));
  OAI211_X1 g499(.A(new_n692_), .B(new_n700_), .C1(new_n694_), .C2(new_n320_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n698_), .A2(new_n699_), .A3(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT40), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n702_), .B(new_n703_), .ZN(G1325gat));
  OAI21_X1  g503(.A(G15gat), .B1(new_n688_), .B2(new_n613_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  XOR2_X1   g505(.A(KEYINPUT101), .B(KEYINPUT41), .Z(new_n707_));
  OR2_X1    g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(G15gat), .ZN(new_n709_));
  INV_X1    g508(.A(new_n613_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n683_), .A2(new_n709_), .A3(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT102), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n706_), .A2(new_n707_), .ZN(new_n713_));
  OR2_X1    g512(.A1(new_n711_), .A2(KEYINPUT102), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n708_), .A2(new_n712_), .A3(new_n713_), .A4(new_n714_), .ZN(G1326gat));
  INV_X1    g514(.A(G22gat), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n683_), .A2(new_n716_), .A3(new_n612_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n638_), .A2(new_n612_), .A3(new_n687_), .ZN(new_n718_));
  XOR2_X1   g517(.A(KEYINPUT103), .B(KEYINPUT42), .Z(new_n719_));
  AND3_X1   g518(.A1(new_n718_), .A2(G22gat), .A3(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(new_n718_), .B2(G22gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n717_), .B1(new_n720_), .B2(new_n721_), .ZN(G1327gat));
  NAND2_X1  g521(.A1(new_n686_), .A2(new_n653_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT104), .ZN(new_n724_));
  NOR3_X1   g523(.A1(new_n351_), .A2(new_n637_), .A3(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(G29gat), .B1(new_n725_), .B2(new_n419_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n679_), .A2(new_n680_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n727_), .B1(new_n615_), .B2(new_n636_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(KEYINPUT43), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT43), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n727_), .B(new_n730_), .C1(new_n615_), .C2(new_n636_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n351_), .B1(new_n729_), .B2(new_n731_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n732_), .A2(KEYINPUT44), .A3(new_n653_), .ZN(new_n733_));
  AND3_X1   g532(.A1(new_n733_), .A2(G29gat), .A3(new_n419_), .ZN(new_n734_));
  AOI21_X1  g533(.A(KEYINPUT44), .B1(new_n732_), .B2(new_n653_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n726_), .B1(new_n734_), .B2(new_n736_), .ZN(G1328gat));
  NAND2_X1  g536(.A1(new_n733_), .A2(new_n693_), .ZN(new_n738_));
  OAI21_X1  g537(.A(G36gat), .B1(new_n738_), .B2(new_n735_), .ZN(new_n739_));
  INV_X1    g538(.A(G36gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n725_), .A2(new_n740_), .A3(new_n693_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT45), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT46), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(KEYINPUT105), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n739_), .A2(new_n742_), .A3(new_n744_), .ZN(new_n745_));
  OR2_X1    g544(.A1(new_n743_), .A2(KEYINPUT105), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n745_), .B(new_n746_), .ZN(G1329gat));
  NAND3_X1  g546(.A1(new_n736_), .A2(G43gat), .A3(new_n733_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n725_), .A2(new_n710_), .ZN(new_n749_));
  OAI22_X1  g548(.A1(new_n748_), .A2(new_n613_), .B1(G43gat), .B2(new_n749_), .ZN(new_n750_));
  XOR2_X1   g549(.A(KEYINPUT106), .B(KEYINPUT47), .Z(new_n751_));
  XNOR2_X1  g550(.A(new_n750_), .B(new_n751_), .ZN(G1330gat));
  AOI21_X1  g551(.A(G50gat), .B1(new_n725_), .B2(new_n612_), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n735_), .A2(new_n302_), .A3(new_n616_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n754_), .B2(new_n733_), .ZN(G1331gat));
  INV_X1    g554(.A(new_n350_), .ZN(new_n756_));
  OAI221_X1 g555(.A(new_n756_), .B1(new_n615_), .B2(new_n636_), .C1(new_n299_), .C2(new_n300_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(new_n682_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(G57gat), .B1(new_n760_), .B2(new_n419_), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n757_), .A2(new_n686_), .A3(new_n653_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n689_), .A2(new_n235_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n761_), .B1(new_n762_), .B2(new_n763_), .ZN(G1332gat));
  AOI21_X1  g563(.A(new_n236_), .B1(new_n762_), .B2(new_n693_), .ZN(new_n765_));
  XOR2_X1   g564(.A(new_n765_), .B(KEYINPUT48), .Z(new_n766_));
  NAND3_X1  g565(.A1(new_n760_), .A2(new_n236_), .A3(new_n693_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(G1333gat));
  INV_X1    g567(.A(G71gat), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n769_), .B1(new_n762_), .B2(new_n710_), .ZN(new_n770_));
  XOR2_X1   g569(.A(new_n770_), .B(KEYINPUT49), .Z(new_n771_));
  NAND2_X1  g570(.A1(new_n710_), .A2(new_n769_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT107), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n771_), .B1(new_n759_), .B2(new_n773_), .ZN(G1334gat));
  NAND2_X1  g573(.A1(new_n762_), .A2(new_n612_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(G78gat), .ZN(new_n776_));
  XNOR2_X1  g575(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n776_), .B(new_n777_), .ZN(new_n778_));
  OR2_X1    g577(.A1(new_n616_), .A2(G78gat), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n778_), .B1(new_n759_), .B2(new_n779_), .ZN(G1335gat));
  NOR2_X1   g579(.A1(new_n757_), .A2(new_n724_), .ZN(new_n781_));
  AOI21_X1  g580(.A(G85gat), .B1(new_n781_), .B2(new_n419_), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n756_), .B(new_n653_), .C1(new_n299_), .C2(new_n300_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT109), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT72), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n293_), .B1(new_n292_), .B2(new_n206_), .ZN(new_n787_));
  AOI211_X1 g586(.A(KEYINPUT71), .B(new_n287_), .C1(new_n291_), .C2(new_n283_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n297_), .B1(new_n789_), .B2(new_n288_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n298_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n786_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n296_), .A2(KEYINPUT72), .A3(new_n298_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n794_), .A2(KEYINPUT109), .A3(new_n756_), .A4(new_n653_), .ZN(new_n795_));
  AOI22_X1  g594(.A1(new_n785_), .A2(new_n795_), .B1(new_n729_), .B2(new_n731_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n419_), .A2(G85gat), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n797_), .B(KEYINPUT110), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n782_), .B1(new_n796_), .B2(new_n798_), .ZN(G1336gat));
  AOI21_X1  g598(.A(G92gat), .B1(new_n781_), .B2(new_n693_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n696_), .A2(new_n564_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n800_), .B1(new_n796_), .B2(new_n801_), .ZN(G1337gat));
  NOR2_X1   g601(.A1(new_n217_), .A2(new_n218_), .ZN(new_n803_));
  NOR4_X1   g602(.A1(new_n757_), .A2(new_n803_), .A3(new_n613_), .A4(new_n724_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT112), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT113), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(KEYINPUT51), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n796_), .A2(new_n710_), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n808_), .A2(KEYINPUT111), .A3(G99gat), .ZN(new_n809_));
  AOI21_X1  g608(.A(KEYINPUT111), .B1(new_n808_), .B2(G99gat), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n805_), .B(new_n807_), .C1(new_n809_), .C2(new_n810_), .ZN(new_n811_));
  OR2_X1    g610(.A1(new_n806_), .A2(KEYINPUT51), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n811_), .B(new_n812_), .ZN(G1338gat));
  AOI221_X4 g612(.A(new_n616_), .B1(new_n729_), .B2(new_n731_), .C1(new_n785_), .C2(new_n795_), .ZN(new_n814_));
  OAI21_X1  g613(.A(KEYINPUT115), .B1(new_n814_), .B2(new_n215_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n785_), .A2(new_n795_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n729_), .A2(new_n731_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n816_), .A2(new_n612_), .A3(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT115), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n818_), .A2(new_n819_), .A3(G106gat), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n815_), .A2(KEYINPUT52), .A3(new_n820_), .ZN(new_n821_));
  NOR4_X1   g620(.A1(new_n757_), .A2(G106gat), .A3(new_n616_), .A4(new_n724_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n822_), .B(KEYINPUT114), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n824_));
  OAI211_X1 g623(.A(KEYINPUT115), .B(new_n824_), .C1(new_n814_), .C2(new_n215_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n821_), .A2(new_n823_), .A3(new_n825_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n828_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n821_), .A2(new_n827_), .A3(new_n823_), .A4(new_n825_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n829_), .A2(new_n830_), .ZN(G1339gat));
  NOR2_X1   g630(.A1(new_n263_), .A2(new_n266_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n274_), .A2(new_n275_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n271_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n834_), .A2(KEYINPUT55), .A3(new_n277_), .ZN(new_n835_));
  OR2_X1    g634(.A1(new_n277_), .A2(KEYINPUT55), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n835_), .A2(new_n206_), .A3(new_n836_), .ZN(new_n837_));
  OR2_X1    g636(.A1(new_n837_), .A2(KEYINPUT56), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(KEYINPUT56), .ZN(new_n839_));
  AND3_X1   g638(.A1(new_n838_), .A2(new_n288_), .A3(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n333_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n332_), .A2(new_n338_), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n841_), .B(new_n347_), .C1(new_n842_), .C2(new_n333_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n843_), .A2(new_n349_), .ZN(new_n844_));
  AOI22_X1  g643(.A1(new_n840_), .A2(new_n350_), .B1(new_n295_), .B2(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n845_), .A2(new_n686_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(KEYINPUT57), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n838_), .A2(new_n288_), .A3(new_n844_), .A4(new_n839_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT58), .ZN(new_n849_));
  OR3_X1    g648(.A1(new_n848_), .A2(KEYINPUT119), .A3(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(KEYINPUT119), .B1(new_n848_), .B2(new_n849_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n848_), .A2(new_n849_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n850_), .A2(new_n851_), .A3(new_n727_), .A4(new_n852_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n854_), .B1(new_n845_), .B2(new_n686_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n847_), .A2(new_n853_), .A3(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n653_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n350_), .B1(new_n296_), .B2(new_n298_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n681_), .ZN(new_n859_));
  OAI21_X1  g658(.A(KEYINPUT117), .B1(new_n859_), .B2(KEYINPUT54), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(KEYINPUT54), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT117), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT54), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n858_), .A2(new_n862_), .A3(new_n681_), .A4(new_n863_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n860_), .A2(new_n861_), .A3(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n857_), .A2(new_n865_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n611_), .A2(new_n689_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(KEYINPUT120), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(G113gat), .B1(new_n870_), .B2(new_n350_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n865_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n853_), .A2(new_n855_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT122), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n853_), .A2(KEYINPUT122), .A3(new_n855_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n875_), .A2(new_n847_), .A3(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n872_), .B1(new_n877_), .B2(new_n653_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n868_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n869_), .A2(KEYINPUT59), .ZN(new_n882_));
  AND2_X1   g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n756_), .A2(new_n386_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n871_), .B1(new_n883_), .B2(new_n884_), .ZN(G1340gat));
  INV_X1    g684(.A(KEYINPUT60), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n886_), .B1(new_n301_), .B2(G120gat), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n870_), .B(new_n887_), .C1(new_n886_), .C2(G120gat), .ZN(new_n888_));
  AND3_X1   g687(.A1(new_n881_), .A2(new_n794_), .A3(new_n882_), .ZN(new_n889_));
  INV_X1    g688(.A(G120gat), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n888_), .B1(new_n889_), .B2(new_n890_), .ZN(G1341gat));
  INV_X1    g690(.A(new_n653_), .ZN(new_n892_));
  AOI21_X1  g691(.A(G127gat), .B1(new_n870_), .B2(new_n892_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n653_), .A2(new_n383_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n893_), .B1(new_n883_), .B2(new_n894_), .ZN(G1342gat));
  AOI21_X1  g694(.A(G134gat), .B1(new_n870_), .B2(new_n686_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n727_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n897_), .A2(new_n384_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n896_), .B1(new_n883_), .B2(new_n898_), .ZN(G1343gat));
  AOI21_X1  g698(.A(new_n693_), .B1(new_n857_), .B2(new_n865_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n616_), .A2(new_n710_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n902_), .A2(new_n689_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n900_), .A2(new_n903_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n904_), .A2(new_n756_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(new_n356_), .ZN(G1344gat));
  NOR2_X1   g705(.A1(new_n904_), .A2(new_n301_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(new_n357_), .ZN(G1345gat));
  NOR2_X1   g707(.A1(new_n904_), .A2(new_n653_), .ZN(new_n909_));
  XOR2_X1   g708(.A(KEYINPUT61), .B(G155gat), .Z(new_n910_));
  XNOR2_X1  g709(.A(new_n909_), .B(new_n910_), .ZN(G1346gat));
  NOR3_X1   g710(.A1(new_n904_), .A2(new_n668_), .A3(new_n897_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n904_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(new_n686_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n912_), .B1(new_n668_), .B2(new_n914_), .ZN(G1347gat));
  NAND3_X1  g714(.A1(new_n689_), .A2(new_n693_), .A3(new_n559_), .ZN(new_n916_));
  OR3_X1    g715(.A1(new_n878_), .A2(KEYINPUT123), .A3(new_n916_), .ZN(new_n917_));
  OAI21_X1  g716(.A(KEYINPUT123), .B1(new_n878_), .B2(new_n916_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(KEYINPUT22), .B(G169gat), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n350_), .A2(new_n919_), .ZN(new_n920_));
  XOR2_X1   g719(.A(new_n920_), .B(KEYINPUT124), .Z(new_n921_));
  NAND3_X1  g720(.A1(new_n917_), .A2(new_n918_), .A3(new_n921_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT62), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n878_), .A2(new_n916_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(new_n350_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n923_), .B1(new_n925_), .B2(G169gat), .ZN(new_n926_));
  AOI211_X1 g725(.A(KEYINPUT62), .B(new_n343_), .C1(new_n924_), .C2(new_n350_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n922_), .B1(new_n926_), .B2(new_n927_), .ZN(G1348gat));
  NAND3_X1  g727(.A1(new_n917_), .A2(new_n794_), .A3(new_n918_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n696_), .B1(new_n857_), .B2(new_n865_), .ZN(new_n930_));
  AND4_X1   g729(.A1(G176gat), .A2(new_n794_), .A3(new_n689_), .A4(new_n559_), .ZN(new_n931_));
  AOI22_X1  g730(.A1(new_n929_), .A2(new_n494_), .B1(new_n930_), .B2(new_n931_), .ZN(G1349gat));
  NOR2_X1   g731(.A1(new_n653_), .A2(new_n570_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n917_), .A2(new_n918_), .A3(new_n933_), .ZN(new_n934_));
  INV_X1    g733(.A(G183gat), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n872_), .A2(new_n892_), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n935_), .B1(new_n936_), .B2(new_n916_), .ZN(new_n937_));
  AND2_X1   g736(.A1(new_n934_), .A2(new_n937_), .ZN(G1350gat));
  NAND3_X1  g737(.A1(new_n917_), .A2(new_n727_), .A3(new_n918_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n939_), .A2(G190gat), .ZN(new_n940_));
  NAND4_X1  g739(.A1(new_n917_), .A2(new_n569_), .A3(new_n686_), .A4(new_n918_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n940_), .A2(new_n941_), .ZN(G1351gat));
  NAND3_X1  g741(.A1(new_n689_), .A2(new_n901_), .A3(KEYINPUT125), .ZN(new_n943_));
  INV_X1    g742(.A(KEYINPUT125), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n944_), .B1(new_n902_), .B2(new_n419_), .ZN(new_n945_));
  NAND4_X1  g744(.A1(new_n866_), .A2(new_n693_), .A3(new_n943_), .A4(new_n945_), .ZN(new_n946_));
  INV_X1    g745(.A(KEYINPUT126), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n946_), .A2(new_n947_), .ZN(new_n948_));
  NAND4_X1  g747(.A1(new_n930_), .A2(KEYINPUT126), .A3(new_n943_), .A4(new_n945_), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n756_), .B1(new_n948_), .B2(new_n949_), .ZN(new_n950_));
  XNOR2_X1  g749(.A(new_n950_), .B(new_n345_), .ZN(G1352gat));
  AOI21_X1  g750(.A(new_n301_), .B1(new_n948_), .B2(new_n949_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n953_));
  XNOR2_X1  g752(.A(new_n952_), .B(new_n953_), .ZN(G1353gat));
  XNOR2_X1  g753(.A(KEYINPUT63), .B(G211gat), .ZN(new_n955_));
  AOI211_X1 g754(.A(new_n653_), .B(new_n955_), .C1(new_n948_), .C2(new_n949_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n948_), .A2(new_n949_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n957_), .A2(new_n892_), .ZN(new_n958_));
  NOR2_X1   g757(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n959_));
  AOI21_X1  g758(.A(new_n956_), .B1(new_n958_), .B2(new_n959_), .ZN(G1354gat));
  AOI21_X1  g759(.A(G218gat), .B1(new_n957_), .B2(new_n686_), .ZN(new_n961_));
  AOI211_X1 g760(.A(new_n443_), .B(new_n897_), .C1(new_n948_), .C2(new_n949_), .ZN(new_n962_));
  NOR2_X1   g761(.A1(new_n961_), .A2(new_n962_), .ZN(G1355gat));
endmodule


