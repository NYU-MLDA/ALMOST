//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 1 0 0 0 1 1 1 1 0 1 0 0 0 0 0 1 1 0 0 1 1 0 1 1 0 0 0 0 0 1 0 1 1 0 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n742_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n802_,
    new_n803_, new_n805_, new_n806_, new_n807_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_, new_n902_, new_n903_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n910_, new_n911_, new_n912_,
    new_n913_, new_n915_, new_n916_, new_n917_, new_n918_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n948_, new_n949_, new_n950_, new_n952_, new_n953_, new_n954_,
    new_n955_, new_n956_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n963_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n972_, new_n973_, new_n974_;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT0), .ZN(new_n203_));
  INV_X1    g002(.A(G57gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G85gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G225gat), .A2(G233gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G155gat), .B(G162gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT3), .ZN(new_n210_));
  INV_X1    g009(.A(G141gat), .ZN(new_n211_));
  INV_X1    g010(.A(G148gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G141gat), .A2(G148gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT2), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n213_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT89), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n220_), .B(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n209_), .B1(new_n219_), .B2(new_n222_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n209_), .A2(KEYINPUT1), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n211_), .A2(new_n212_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(new_n214_), .A3(new_n226_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n224_), .A2(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT90), .B1(new_n223_), .B2(new_n228_), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n224_), .A2(new_n227_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n209_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n220_), .B(KEYINPUT89), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n231_), .B1(new_n232_), .B2(new_n218_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT90), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n230_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  XOR2_X1   g034(.A(G127gat), .B(G134gat), .Z(new_n236_));
  XOR2_X1   g035(.A(G113gat), .B(G120gat), .Z(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n229_), .A2(new_n235_), .A3(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n240_), .A2(KEYINPUT4), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n223_), .A2(new_n228_), .ZN(new_n242_));
  AOI21_X1  g041(.A(KEYINPUT96), .B1(new_n242_), .B2(new_n238_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n240_), .A2(new_n243_), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n229_), .A2(new_n235_), .A3(KEYINPUT96), .A4(new_n239_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  AOI211_X1 g045(.A(new_n208_), .B(new_n241_), .C1(new_n246_), .C2(KEYINPUT4), .ZN(new_n247_));
  INV_X1    g046(.A(new_n208_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n248_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n207_), .B1(new_n247_), .B2(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n241_), .B1(new_n246_), .B2(KEYINPUT4), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(new_n248_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n249_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n207_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n252_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n250_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G8gat), .B(G36gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G64gat), .B(G92gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G226gat), .A2(G233gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT19), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT93), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G197gat), .B(G204gat), .ZN(new_n268_));
  XOR2_X1   g067(.A(G211gat), .B(G218gat), .Z(new_n269_));
  INV_X1    g068(.A(KEYINPUT21), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n268_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G211gat), .B(G218gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(KEYINPUT21), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n272_), .A2(new_n268_), .A3(KEYINPUT21), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(G169gat), .ZN(new_n277_));
  INV_X1    g076(.A(G176gat), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n277_), .A2(new_n278_), .A3(KEYINPUT83), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT83), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n280_), .B1(G169gat), .B2(G176gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n279_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT24), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(KEYINPUT25), .B(G183gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT26), .B(G190gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G169gat), .A2(G176gat), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n279_), .A2(new_n281_), .A3(KEYINPUT24), .A4(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G183gat), .A2(G190gat), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT23), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n293_));
  AND2_X1   g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n284_), .A2(new_n287_), .A3(new_n289_), .A4(new_n294_), .ZN(new_n295_));
  OR2_X1    g094(.A1(G183gat), .A2(G190gat), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n292_), .A2(new_n296_), .A3(new_n293_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n277_), .A2(KEYINPUT22), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT22), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(G169gat), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n298_), .A2(new_n300_), .A3(new_n278_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n297_), .A2(new_n301_), .A3(new_n288_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n295_), .A2(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n267_), .B1(new_n276_), .B2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n276_), .A2(new_n303_), .A3(new_n267_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n301_), .A2(KEYINPUT84), .ZN(new_n308_));
  XNOR2_X1  g107(.A(KEYINPUT22), .B(G169gat), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT84), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n309_), .A2(new_n310_), .A3(new_n278_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n308_), .A2(new_n311_), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n292_), .A2(new_n296_), .A3(KEYINPUT85), .A4(new_n293_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT85), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n297_), .A2(new_n314_), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n312_), .A2(new_n288_), .A3(new_n313_), .A4(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(new_n295_), .ZN(new_n317_));
  OAI21_X1  g116(.A(KEYINPUT20), .B1(new_n317_), .B2(new_n276_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n266_), .B1(new_n307_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n276_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n303_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT94), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n321_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT94), .B1(new_n276_), .B2(new_n303_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n266_), .A2(KEYINPUT20), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n327_), .B1(new_n317_), .B2(new_n276_), .ZN(new_n328_));
  AND2_X1   g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n263_), .B1(new_n320_), .B2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n326_), .A2(new_n328_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n321_), .A2(new_n295_), .A3(new_n316_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n306_), .ZN(new_n333_));
  OAI211_X1 g132(.A(KEYINPUT20), .B(new_n332_), .C1(new_n333_), .C2(new_n304_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n262_), .B(new_n331_), .C1(new_n335_), .C2(new_n266_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n330_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT27), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n317_), .A2(new_n276_), .ZN(new_n340_));
  OAI21_X1  g139(.A(KEYINPUT20), .B1(new_n276_), .B2(new_n303_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n265_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n342_), .B1(new_n334_), .B2(new_n265_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(new_n263_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n336_), .A2(new_n344_), .A3(KEYINPUT27), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n257_), .A2(new_n339_), .A3(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n229_), .A2(new_n235_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT29), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G78gat), .B(G106gat), .ZN(new_n351_));
  XOR2_X1   g150(.A(new_n350_), .B(new_n351_), .Z(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G22gat), .B(G50gat), .ZN(new_n354_));
  XOR2_X1   g153(.A(new_n354_), .B(KEYINPUT28), .Z(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n229_), .A2(new_n235_), .A3(KEYINPUT29), .ZN(new_n357_));
  OR2_X1    g156(.A1(new_n357_), .A2(KEYINPUT91), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n321_), .B1(new_n357_), .B2(KEYINPUT91), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G228gat), .A2(G233gat), .ZN(new_n361_));
  XOR2_X1   g160(.A(new_n361_), .B(KEYINPUT92), .Z(new_n362_));
  NAND2_X1  g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n362_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n276_), .B(new_n364_), .C1(new_n242_), .C2(new_n349_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n356_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n364_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n365_), .ZN(new_n368_));
  NOR3_X1   g167(.A1(new_n367_), .A2(new_n368_), .A3(new_n355_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n353_), .B1(new_n366_), .B2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n363_), .A2(new_n365_), .A3(new_n356_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n355_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n371_), .A2(new_n352_), .A3(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n370_), .A2(new_n373_), .ZN(new_n374_));
  XOR2_X1   g173(.A(G71gat), .B(G99gat), .Z(new_n375_));
  XOR2_X1   g174(.A(G15gat), .B(G43gat), .Z(new_n376_));
  XOR2_X1   g175(.A(new_n375_), .B(new_n376_), .Z(new_n377_));
  NAND3_X1  g176(.A1(new_n316_), .A2(KEYINPUT30), .A3(new_n295_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(KEYINPUT30), .B1(new_n316_), .B2(new_n295_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n377_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G227gat), .A2(G233gat), .ZN(new_n382_));
  XOR2_X1   g181(.A(new_n382_), .B(KEYINPUT86), .Z(new_n383_));
  INV_X1    g182(.A(KEYINPUT30), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n317_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n377_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(new_n378_), .A3(new_n386_), .ZN(new_n387_));
  AND3_X1   g186(.A1(new_n381_), .A2(new_n383_), .A3(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n383_), .B1(new_n381_), .B2(new_n387_), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT87), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n383_), .ZN(new_n391_));
  NOR3_X1   g190(.A1(new_n379_), .A2(new_n380_), .A3(new_n377_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n386_), .B1(new_n385_), .B2(new_n378_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n391_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT87), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n381_), .A2(new_n383_), .A3(new_n387_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n394_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n238_), .B(KEYINPUT31), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n390_), .A2(new_n397_), .A3(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n398_), .ZN(new_n400_));
  OAI211_X1 g199(.A(KEYINPUT87), .B(new_n400_), .C1(new_n388_), .C2(new_n389_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT88), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n399_), .A2(KEYINPUT88), .A3(new_n401_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n374_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  NOR3_X1   g205(.A1(new_n366_), .A2(new_n369_), .A3(new_n353_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n352_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n409_), .A2(new_n402_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n347_), .B1(new_n406_), .B2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n404_), .A2(new_n405_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n249_), .B1(new_n251_), .B2(new_n248_), .ZN(new_n413_));
  AOI21_X1  g212(.A(KEYINPUT33), .B1(new_n413_), .B2(new_n254_), .ZN(new_n414_));
  AOI211_X1 g213(.A(new_n248_), .B(new_n241_), .C1(new_n246_), .C2(KEYINPUT4), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n246_), .A2(new_n248_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(new_n207_), .ZN(new_n417_));
  OAI211_X1 g216(.A(new_n330_), .B(new_n336_), .C1(new_n415_), .C2(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n414_), .A2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n413_), .A2(KEYINPUT33), .A3(new_n254_), .ZN(new_n420_));
  AND2_X1   g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n343_), .A2(KEYINPUT32), .A3(new_n262_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n262_), .A2(KEYINPUT32), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n423_), .B(new_n331_), .C1(new_n335_), .C2(new_n266_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n425_), .B1(new_n250_), .B2(new_n255_), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n412_), .B(new_n374_), .C1(new_n421_), .C2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n411_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT64), .ZN(new_n429_));
  AND2_X1   g228(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n430_));
  NOR2_X1   g229(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(G106gat), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n429_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NOR4_X1   g233(.A1(new_n430_), .A2(new_n431_), .A3(KEYINPUT64), .A4(G106gat), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G99gat), .A2(G106gat), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT6), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(G92gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n206_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G85gat), .A2(G92gat), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n443_), .A2(KEYINPUT9), .A3(new_n444_), .ZN(new_n445_));
  OR2_X1    g244(.A1(new_n444_), .A2(KEYINPUT9), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n441_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  NOR3_X1   g246(.A1(new_n436_), .A2(KEYINPUT65), .A3(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT65), .ZN(new_n449_));
  XNOR2_X1  g248(.A(KEYINPUT10), .B(G99gat), .ZN(new_n450_));
  OAI21_X1  g249(.A(KEYINPUT64), .B1(new_n450_), .B2(G106gat), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n432_), .A2(new_n429_), .A3(new_n433_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n445_), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n439_), .B(new_n440_), .C1(KEYINPUT9), .C2(new_n444_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n449_), .B1(new_n453_), .B2(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT69), .B1(new_n448_), .B2(new_n457_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(G99gat), .A2(G106gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(KEYINPUT7), .ZN(new_n460_));
  NAND2_X1  g259(.A1(KEYINPUT66), .A2(KEYINPUT6), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(KEYINPUT66), .A2(KEYINPUT6), .ZN(new_n463_));
  OAI211_X1 g262(.A(G99gat), .B(G106gat), .C1(new_n462_), .C2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n463_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n465_), .A2(new_n437_), .A3(new_n461_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n460_), .A2(new_n464_), .A3(new_n466_), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n443_), .A2(new_n444_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT8), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT8), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n468_), .A2(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n472_), .B1(new_n460_), .B2(new_n441_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n470_), .A2(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT65), .B1(new_n436_), .B2(new_n447_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT69), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n453_), .A2(new_n456_), .A3(new_n449_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n476_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n458_), .A2(new_n475_), .A3(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(G36gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(G29gat), .ZN(new_n482_));
  INV_X1    g281(.A(G29gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(G36gat), .ZN(new_n484_));
  INV_X1    g283(.A(G43gat), .ZN(new_n485_));
  AND3_X1   g284(.A1(new_n482_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n485_), .B1(new_n482_), .B2(new_n484_), .ZN(new_n487_));
  OAI21_X1  g286(.A(KEYINPUT72), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n483_), .A2(G36gat), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n481_), .A2(G29gat), .ZN(new_n490_));
  OAI21_X1  g289(.A(G43gat), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT72), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n482_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n491_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n488_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(G50gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n488_), .A2(new_n494_), .A3(G50gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(KEYINPUT73), .B(KEYINPUT15), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n497_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n499_), .ZN(new_n501_));
  AND3_X1   g300(.A1(new_n488_), .A2(new_n494_), .A3(G50gat), .ZN(new_n502_));
  AOI21_X1  g301(.A(G50gat), .B1(new_n488_), .B2(new_n494_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n501_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n480_), .A2(new_n500_), .A3(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n476_), .A2(new_n478_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n471_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n507_), .A2(new_n473_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n502_), .A2(new_n503_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT35), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G232gat), .A2(G233gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT34), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  AOI22_X1  g313(.A1(new_n509_), .A2(new_n510_), .B1(new_n511_), .B2(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n514_), .A2(new_n511_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n505_), .A2(new_n515_), .A3(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n517_), .B1(new_n505_), .B2(new_n515_), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT76), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n505_), .A2(new_n515_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(new_n516_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT76), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n523_), .A2(new_n524_), .A3(new_n518_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G190gat), .B(G218gat), .ZN(new_n526_));
  INV_X1    g325(.A(G134gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT74), .ZN(new_n529_));
  INV_X1    g328(.A(G162gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT36), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n521_), .A2(new_n525_), .A3(new_n534_), .ZN(new_n535_));
  AND2_X1   g334(.A1(new_n531_), .A2(new_n532_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n523_), .A2(new_n536_), .A3(new_n518_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n535_), .A2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G127gat), .B(G155gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G183gat), .B(G211gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n543_), .A2(KEYINPUT17), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(KEYINPUT17), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT79), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(KEYINPUT77), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT77), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n545_), .A2(new_n549_), .A3(new_n546_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G15gat), .B(G22gat), .ZN(new_n552_));
  INV_X1    g351(.A(G1gat), .ZN(new_n553_));
  INV_X1    g352(.A(G8gat), .ZN(new_n554_));
  OAI21_X1  g353(.A(KEYINPUT14), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n552_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G1gat), .B(G8gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n551_), .A2(new_n558_), .ZN(new_n559_));
  XOR2_X1   g358(.A(new_n556_), .B(new_n557_), .Z(new_n560_));
  NAND3_X1  g359(.A1(new_n548_), .A2(new_n560_), .A3(new_n550_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n559_), .A2(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G57gat), .B(G64gat), .ZN(new_n563_));
  AND2_X1   g362(.A1(new_n563_), .A2(KEYINPUT11), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n563_), .A2(KEYINPUT11), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G71gat), .B(G78gat), .ZN(new_n566_));
  OR3_X1    g365(.A1(new_n564_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n563_), .A2(new_n566_), .A3(KEYINPUT11), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  AND2_X1   g368(.A1(G231gat), .A2(G233gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n544_), .B1(new_n562_), .B2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n559_), .A2(new_n571_), .A3(new_n561_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n428_), .A2(new_n538_), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(G120gat), .B(G148gat), .Z(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(G204gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(KEYINPUT5), .B(G176gat), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n579_), .B(new_n580_), .Z(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT12), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n569_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n480_), .A2(new_n584_), .ZN(new_n585_));
  AND2_X1   g384(.A1(G230gat), .A2(G233gat), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n586_), .B1(new_n509_), .B2(new_n569_), .ZN(new_n587_));
  OAI211_X1 g386(.A(new_n476_), .B(new_n478_), .C1(new_n507_), .C2(new_n473_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n569_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(new_n583_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n585_), .A2(new_n587_), .A3(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(KEYINPUT67), .B1(new_n588_), .B2(new_n589_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n448_), .A2(new_n457_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT67), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n595_), .A2(new_n475_), .A3(new_n596_), .A4(new_n569_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n594_), .A2(new_n590_), .A3(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(new_n586_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(KEYINPUT68), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT68), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n598_), .A2(new_n601_), .A3(new_n586_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n593_), .B1(new_n600_), .B2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT70), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n582_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  AND3_X1   g404(.A1(new_n598_), .A2(new_n601_), .A3(new_n586_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n601_), .B1(new_n598_), .B2(new_n586_), .ZN(new_n607_));
  OAI211_X1 g406(.A(new_n604_), .B(new_n592_), .C1(new_n606_), .C2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(KEYINPUT71), .B1(new_n605_), .B2(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n592_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(KEYINPUT70), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT71), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n612_), .A2(new_n613_), .A3(new_n608_), .A4(new_n582_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n603_), .A2(new_n581_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n610_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT13), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n504_), .A2(new_n500_), .A3(new_n558_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(G229gat), .A2(G233gat), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n497_), .A2(new_n560_), .A3(new_n498_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n619_), .A2(new_n620_), .A3(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(KEYINPUT81), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT81), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n619_), .A2(new_n624_), .A3(new_n620_), .A4(new_n621_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n620_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n558_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n627_), .A2(new_n621_), .A3(KEYINPUT80), .ZN(new_n628_));
  AOI21_X1  g427(.A(KEYINPUT80), .B1(new_n627_), .B2(new_n621_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n626_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n623_), .A2(new_n625_), .A3(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(G113gat), .B(G141gat), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(G169gat), .ZN(new_n633_));
  INV_X1    g432(.A(G197gat), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n631_), .A2(new_n636_), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n623_), .A2(new_n630_), .A3(new_n625_), .A4(new_n635_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n638_), .A2(KEYINPUT82), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n638_), .A2(KEYINPUT82), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n637_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n612_), .A2(new_n608_), .A3(new_n582_), .ZN(new_n642_));
  AOI22_X1  g441(.A1(new_n642_), .A2(KEYINPUT71), .B1(new_n603_), .B2(new_n581_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n643_), .A2(KEYINPUT13), .A3(new_n614_), .ZN(new_n644_));
  AND3_X1   g443(.A1(new_n618_), .A2(new_n641_), .A3(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n577_), .A2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT99), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(new_n256_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(G1gat), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT38), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n638_), .A2(KEYINPUT82), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n638_), .A2(KEYINPUT82), .ZN(new_n652_));
  AOI22_X1  g451(.A1(new_n651_), .A2(new_n652_), .B1(new_n631_), .B2(new_n636_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n653_), .B1(new_n411_), .B2(new_n427_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT97), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n618_), .A2(new_n644_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n537_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n533_), .B1(new_n523_), .B2(new_n518_), .ZN(new_n659_));
  OAI21_X1  g458(.A(KEYINPUT37), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(KEYINPUT75), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT37), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n535_), .A2(new_n662_), .A3(new_n537_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT75), .ZN(new_n664_));
  OAI211_X1 g463(.A(new_n664_), .B(KEYINPUT37), .C1(new_n658_), .C2(new_n659_), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n661_), .A2(new_n663_), .A3(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n575_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n655_), .A2(new_n657_), .A3(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(KEYINPUT98), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT98), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n655_), .A2(new_n671_), .A3(new_n657_), .A4(new_n668_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n257_), .A2(G1gat), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n670_), .A2(new_n672_), .A3(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT100), .ZN(new_n675_));
  AND3_X1   g474(.A1(new_n674_), .A2(new_n675_), .A3(new_n650_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n674_), .B2(new_n650_), .ZN(new_n677_));
  OAI221_X1 g476(.A(new_n649_), .B1(new_n650_), .B2(new_n674_), .C1(new_n676_), .C2(new_n677_), .ZN(G1324gat));
  NAND2_X1  g477(.A1(new_n339_), .A2(new_n345_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(G8gat), .B1(new_n646_), .B2(new_n680_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT39), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n670_), .A2(new_n672_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n679_), .A2(new_n554_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n682_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT40), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  OAI211_X1 g486(.A(new_n682_), .B(KEYINPUT40), .C1(new_n683_), .C2(new_n684_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1325gat));
  OR3_X1    g488(.A1(new_n683_), .A2(G15gat), .A3(new_n412_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n412_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n647_), .A2(new_n691_), .ZN(new_n692_));
  AND3_X1   g491(.A1(new_n692_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n693_));
  AOI21_X1  g492(.A(KEYINPUT41), .B1(new_n692_), .B2(G15gat), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n690_), .B1(new_n693_), .B2(new_n694_), .ZN(G1326gat));
  NAND2_X1  g494(.A1(new_n647_), .A2(new_n409_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT42), .ZN(new_n697_));
  AND3_X1   g496(.A1(new_n696_), .A2(new_n697_), .A3(G22gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n697_), .B1(new_n696_), .B2(G22gat), .ZN(new_n699_));
  OR2_X1    g498(.A1(new_n374_), .A2(G22gat), .ZN(new_n700_));
  OAI22_X1  g499(.A1(new_n698_), .A2(new_n699_), .B1(new_n683_), .B2(new_n700_), .ZN(G1327gat));
  INV_X1    g500(.A(KEYINPUT43), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n702_), .B1(new_n428_), .B2(new_n666_), .ZN(new_n703_));
  AND3_X1   g502(.A1(new_n399_), .A2(KEYINPUT88), .A3(new_n401_), .ZN(new_n704_));
  AOI21_X1  g503(.A(KEYINPUT88), .B1(new_n399_), .B2(new_n401_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n409_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n402_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(new_n374_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n346_), .B1(new_n706_), .B2(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n374_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n426_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  OAI211_X1 g511(.A(new_n702_), .B(new_n666_), .C1(new_n709_), .C2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n667_), .B(new_n645_), .C1(new_n703_), .C2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n666_), .B1(new_n709_), .B2(new_n712_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(KEYINPUT43), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n575_), .B1(new_n719_), .B2(new_n713_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n720_), .A2(KEYINPUT44), .A3(new_n645_), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n717_), .A2(new_n721_), .A3(G29gat), .A4(new_n256_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n538_), .A2(new_n575_), .ZN(new_n723_));
  AND4_X1   g522(.A1(new_n256_), .A2(new_n655_), .A3(new_n657_), .A4(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n722_), .B1(G29gat), .B2(new_n724_), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n725_), .B(KEYINPUT101), .Z(G1328gat));
  NAND3_X1  g525(.A1(new_n717_), .A2(new_n679_), .A3(new_n721_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(KEYINPUT102), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT102), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n717_), .A2(new_n721_), .A3(new_n729_), .A4(new_n679_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n728_), .A2(G36gat), .A3(new_n730_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n680_), .A2(G36gat), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n655_), .A2(new_n657_), .A3(new_n723_), .A4(new_n732_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT45), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n731_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT46), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n731_), .A2(new_n734_), .A3(KEYINPUT46), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(G1329gat));
  NAND4_X1  g538(.A1(new_n717_), .A2(new_n721_), .A3(G43gat), .A4(new_n707_), .ZN(new_n740_));
  AND4_X1   g539(.A1(new_n691_), .A2(new_n655_), .A3(new_n657_), .A4(new_n723_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n740_), .B1(G43gat), .B2(new_n741_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g542(.A1(new_n374_), .A2(G50gat), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n655_), .A2(new_n657_), .A3(new_n723_), .A4(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n717_), .A2(new_n409_), .A3(new_n721_), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n746_), .A2(KEYINPUT103), .A3(G50gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(KEYINPUT103), .B1(new_n746_), .B2(G50gat), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n745_), .B1(new_n747_), .B2(new_n748_), .ZN(G1331gat));
  AOI21_X1  g548(.A(new_n641_), .B1(new_n618_), .B2(new_n644_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n666_), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n750_), .A2(new_n428_), .A3(new_n751_), .A4(new_n575_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT104), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n753_), .A2(new_n204_), .A3(new_n256_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n577_), .A2(new_n750_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT105), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n577_), .A2(KEYINPUT105), .A3(new_n750_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n757_), .A2(new_n256_), .A3(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(G57gat), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n754_), .A2(new_n760_), .ZN(G1332gat));
  NOR2_X1   g560(.A1(new_n680_), .A2(G64gat), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT107), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n753_), .A2(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n757_), .A2(new_n679_), .A3(new_n758_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(G64gat), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT106), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT106), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n765_), .A2(new_n768_), .A3(G64gat), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n767_), .A2(KEYINPUT48), .A3(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(KEYINPUT48), .B1(new_n767_), .B2(new_n769_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n764_), .B1(new_n770_), .B2(new_n771_), .ZN(G1333gat));
  NOR2_X1   g571(.A1(new_n412_), .A2(G71gat), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT109), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n753_), .A2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n757_), .A2(new_n691_), .A3(new_n758_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(G71gat), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT108), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT108), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n776_), .A2(new_n779_), .A3(G71gat), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n778_), .A2(KEYINPUT49), .A3(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(KEYINPUT49), .B1(new_n778_), .B2(new_n780_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n775_), .B1(new_n781_), .B2(new_n782_), .ZN(G1334gat));
  INV_X1    g582(.A(G78gat), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n753_), .A2(new_n784_), .A3(new_n409_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n757_), .A2(new_n409_), .A3(new_n758_), .ZN(new_n786_));
  XOR2_X1   g585(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n787_));
  AND3_X1   g586(.A1(new_n786_), .A2(G78gat), .A3(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n787_), .B1(new_n786_), .B2(G78gat), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n785_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT111), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n785_), .B(KEYINPUT111), .C1(new_n788_), .C2(new_n789_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(G1335gat));
  NAND2_X1  g593(.A1(new_n720_), .A2(new_n750_), .ZN(new_n795_));
  XOR2_X1   g594(.A(new_n795_), .B(KEYINPUT112), .Z(new_n796_));
  OAI21_X1  g595(.A(G85gat), .B1(new_n796_), .B2(new_n257_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n750_), .A2(new_n428_), .A3(new_n723_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n799_), .A2(new_n206_), .A3(new_n256_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n797_), .A2(new_n800_), .ZN(G1336gat));
  OAI21_X1  g600(.A(G92gat), .B1(new_n796_), .B2(new_n680_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n799_), .A2(new_n442_), .A3(new_n679_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(G1337gat));
  OAI21_X1  g603(.A(G99gat), .B1(new_n795_), .B2(new_n412_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n799_), .A2(new_n707_), .A3(new_n432_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n807_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g607(.A1(new_n799_), .A2(new_n433_), .A3(new_n409_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n720_), .A2(new_n409_), .A3(new_n750_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT113), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n433_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT52), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n720_), .A2(KEYINPUT113), .A3(new_n409_), .A4(new_n750_), .ZN(new_n814_));
  AND3_X1   g613(.A1(new_n812_), .A2(new_n813_), .A3(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n813_), .B1(new_n812_), .B2(new_n814_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n809_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(KEYINPUT53), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT53), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n819_), .B(new_n809_), .C1(new_n815_), .C2(new_n816_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n820_), .ZN(G1339gat));
  INV_X1    g620(.A(KEYINPUT114), .ZN(new_n822_));
  AND3_X1   g621(.A1(new_n653_), .A2(new_n575_), .A3(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n822_), .B1(new_n653_), .B2(new_n575_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n618_), .A2(new_n644_), .A3(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(KEYINPUT115), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT115), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n618_), .A2(new_n825_), .A3(new_n644_), .A4(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT117), .ZN(new_n830_));
  XOR2_X1   g629(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n666_), .B1(new_n830_), .B2(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n827_), .A2(new_n829_), .A3(new_n833_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n832_), .A2(new_n830_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n835_), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n827_), .A2(new_n837_), .A3(new_n829_), .A4(new_n833_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT57), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n585_), .A2(new_n591_), .A3(new_n594_), .A4(new_n597_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n586_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT55), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n592_), .A2(new_n842_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n585_), .A2(new_n587_), .A3(new_n591_), .A4(KEYINPUT55), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n841_), .A2(new_n843_), .A3(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n582_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(KEYINPUT56), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT56), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n845_), .A2(new_n848_), .A3(new_n582_), .ZN(new_n849_));
  AND4_X1   g648(.A1(new_n641_), .A2(new_n847_), .A3(new_n615_), .A4(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n620_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n619_), .A2(new_n626_), .A3(new_n621_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n851_), .A2(new_n636_), .A3(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n853_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(KEYINPUT118), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT118), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n856_), .B(new_n853_), .C1(new_n639_), .C2(new_n640_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n850_), .B1(new_n616_), .B2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n538_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n839_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  AOI22_X1  g660(.A1(new_n643_), .A2(new_n614_), .B1(new_n857_), .B2(new_n855_), .ZN(new_n862_));
  OAI211_X1 g661(.A(KEYINPUT57), .B(new_n538_), .C1(new_n862_), .C2(new_n850_), .ZN(new_n863_));
  AND3_X1   g662(.A1(new_n847_), .A2(new_n615_), .A3(new_n849_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n858_), .A2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT58), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n858_), .A2(new_n864_), .A3(KEYINPUT58), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n867_), .A2(new_n666_), .A3(new_n868_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n861_), .A2(new_n863_), .A3(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n667_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n836_), .A2(new_n838_), .A3(new_n871_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n708_), .A2(new_n257_), .A3(new_n679_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(G113gat), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n874_), .A2(new_n875_), .A3(new_n641_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT59), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n873_), .A2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT119), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n871_), .A2(new_n879_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n870_), .A2(KEYINPUT119), .A3(new_n667_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  AND2_X1   g681(.A1(new_n836_), .A2(new_n838_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n878_), .B1(new_n882_), .B2(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n877_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n884_), .A2(new_n885_), .A3(new_n653_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n876_), .B1(new_n886_), .B2(new_n875_), .ZN(G1340gat));
  INV_X1    g686(.A(G120gat), .ZN(new_n888_));
  AOI21_X1  g687(.A(KEYINPUT60), .B1(new_n656_), .B2(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n889_), .B1(KEYINPUT60), .B2(new_n888_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n872_), .A2(new_n873_), .A3(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT120), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n891_), .B(new_n892_), .ZN(new_n893_));
  NOR3_X1   g692(.A1(new_n884_), .A2(new_n885_), .A3(new_n657_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n894_), .B2(new_n888_), .ZN(G1341gat));
  INV_X1    g694(.A(G127gat), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n874_), .A2(new_n896_), .A3(new_n575_), .ZN(new_n897_));
  NOR3_X1   g696(.A1(new_n884_), .A2(new_n885_), .A3(new_n667_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n898_), .B2(new_n896_), .ZN(G1342gat));
  AOI21_X1  g698(.A(G134gat), .B1(new_n874_), .B2(new_n860_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n884_), .A2(new_n885_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n666_), .A2(G134gat), .ZN(new_n902_));
  XOR2_X1   g701(.A(new_n902_), .B(KEYINPUT121), .Z(new_n903_));
  AOI21_X1  g702(.A(new_n900_), .B1(new_n901_), .B2(new_n903_), .ZN(G1343gat));
  AND2_X1   g703(.A1(new_n872_), .A2(new_n406_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n257_), .A2(new_n679_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n905_), .A2(new_n641_), .A3(new_n906_), .ZN(new_n907_));
  XOR2_X1   g706(.A(KEYINPUT122), .B(G141gat), .Z(new_n908_));
  XNOR2_X1  g707(.A(new_n907_), .B(new_n908_), .ZN(G1344gat));
  NAND2_X1  g708(.A1(new_n905_), .A2(new_n906_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n911_), .A2(new_n212_), .A3(new_n656_), .ZN(new_n912_));
  OAI21_X1  g711(.A(G148gat), .B1(new_n910_), .B2(new_n657_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(G1345gat));
  XNOR2_X1  g713(.A(KEYINPUT61), .B(G155gat), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n911_), .A2(new_n575_), .A3(new_n916_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n915_), .B1(new_n910_), .B2(new_n667_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(G1346gat));
  NAND4_X1  g718(.A1(new_n872_), .A2(new_n406_), .A3(new_n860_), .A4(new_n906_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(new_n530_), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT123), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n920_), .A2(KEYINPUT123), .A3(new_n530_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n666_), .A2(G162gat), .ZN(new_n925_));
  XOR2_X1   g724(.A(new_n925_), .B(KEYINPUT124), .Z(new_n926_));
  AOI22_X1  g725(.A1(new_n923_), .A2(new_n924_), .B1(new_n911_), .B2(new_n926_), .ZN(G1347gat));
  NOR2_X1   g726(.A1(new_n680_), .A2(new_n256_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n691_), .A2(new_n928_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n929_), .A2(new_n409_), .ZN(new_n930_));
  AND3_X1   g729(.A1(new_n870_), .A2(KEYINPUT119), .A3(new_n667_), .ZN(new_n931_));
  AOI21_X1  g730(.A(KEYINPUT119), .B1(new_n870_), .B2(new_n667_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n931_), .A2(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n836_), .A2(new_n838_), .ZN(new_n934_));
  OAI211_X1 g733(.A(new_n641_), .B(new_n930_), .C1(new_n933_), .C2(new_n934_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(G169gat), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT62), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n936_), .A2(new_n937_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n935_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n882_), .A2(new_n883_), .ZN(new_n940_));
  NAND4_X1  g739(.A1(new_n940_), .A2(new_n641_), .A3(new_n309_), .A4(new_n930_), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n938_), .A2(new_n939_), .A3(new_n941_), .ZN(G1348gat));
  NAND2_X1  g741(.A1(new_n872_), .A2(new_n374_), .ZN(new_n943_));
  NOR4_X1   g742(.A1(new_n943_), .A2(new_n278_), .A3(new_n657_), .A4(new_n929_), .ZN(new_n944_));
  AND2_X1   g743(.A1(new_n940_), .A2(new_n930_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n945_), .A2(new_n656_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n944_), .B1(new_n946_), .B2(new_n278_), .ZN(G1349gat));
  INV_X1    g746(.A(G183gat), .ZN(new_n948_));
  OR3_X1    g747(.A1(new_n943_), .A2(new_n667_), .A3(new_n929_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n667_), .A2(new_n285_), .ZN(new_n950_));
  AOI22_X1  g749(.A1(new_n948_), .A2(new_n949_), .B1(new_n945_), .B2(new_n950_), .ZN(G1350gat));
  NAND4_X1  g750(.A1(new_n940_), .A2(new_n286_), .A3(new_n860_), .A4(new_n930_), .ZN(new_n952_));
  OAI211_X1 g751(.A(new_n666_), .B(new_n930_), .C1(new_n933_), .C2(new_n934_), .ZN(new_n953_));
  INV_X1    g752(.A(KEYINPUT125), .ZN(new_n954_));
  AND3_X1   g753(.A1(new_n953_), .A2(new_n954_), .A3(G190gat), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n954_), .B1(new_n953_), .B2(G190gat), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n952_), .B1(new_n955_), .B2(new_n956_), .ZN(G1351gat));
  NAND4_X1  g756(.A1(new_n872_), .A2(new_n641_), .A3(new_n406_), .A4(new_n928_), .ZN(new_n958_));
  AND3_X1   g757(.A1(new_n958_), .A2(KEYINPUT126), .A3(new_n634_), .ZN(new_n959_));
  AOI21_X1  g758(.A(KEYINPUT126), .B1(new_n958_), .B2(new_n634_), .ZN(new_n960_));
  NOR2_X1   g759(.A1(new_n958_), .A2(new_n634_), .ZN(new_n961_));
  NOR3_X1   g760(.A1(new_n959_), .A2(new_n960_), .A3(new_n961_), .ZN(G1352gat));
  NAND3_X1  g761(.A1(new_n905_), .A2(new_n656_), .A3(new_n928_), .ZN(new_n963_));
  XNOR2_X1  g762(.A(new_n963_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g763(.A(new_n667_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n965_));
  NAND4_X1  g764(.A1(new_n872_), .A2(new_n406_), .A3(new_n928_), .A4(new_n965_), .ZN(new_n966_));
  NOR2_X1   g765(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n967_));
  AND3_X1   g766(.A1(new_n966_), .A2(KEYINPUT127), .A3(new_n967_), .ZN(new_n968_));
  AOI21_X1  g767(.A(KEYINPUT127), .B1(new_n966_), .B2(new_n967_), .ZN(new_n969_));
  NOR2_X1   g768(.A1(new_n966_), .A2(new_n967_), .ZN(new_n970_));
  NOR3_X1   g769(.A1(new_n968_), .A2(new_n969_), .A3(new_n970_), .ZN(G1354gat));
  NAND2_X1  g770(.A1(new_n905_), .A2(new_n928_), .ZN(new_n972_));
  OAI21_X1  g771(.A(G218gat), .B1(new_n972_), .B2(new_n751_), .ZN(new_n973_));
  OR2_X1    g772(.A1(new_n538_), .A2(G218gat), .ZN(new_n974_));
  OAI21_X1  g773(.A(new_n973_), .B1(new_n972_), .B2(new_n974_), .ZN(G1355gat));
endmodule


