//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 0 0 1 1 1 0 1 0 0 1 1 0 0 1 0 1 0 0 1 1 0 0 0 0 1 0 0 1 0 1 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 0 0 1 0 0 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n700_,
    new_n701_, new_n702_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n872_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n904_, new_n905_, new_n906_,
    new_n907_, new_n908_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n921_, new_n922_, new_n923_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n930_, new_n931_;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202_));
  INV_X1    g001(.A(G1gat), .ZN(new_n203_));
  INV_X1    g002(.A(G8gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT14), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n202_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G1gat), .B(G8gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G29gat), .B(G36gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G43gat), .B(G50gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n209_), .B(new_n210_), .ZN(new_n211_));
  XOR2_X1   g010(.A(new_n208_), .B(new_n211_), .Z(new_n212_));
  NAND2_X1  g011(.A1(G229gat), .A2(G233gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT74), .B(KEYINPUT15), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n211_), .B(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(new_n208_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n208_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(new_n211_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n218_), .A2(new_n220_), .A3(new_n213_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n215_), .A2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G113gat), .B(G141gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G169gat), .B(G197gat), .ZN(new_n224_));
  XOR2_X1   g023(.A(new_n223_), .B(new_n224_), .Z(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT80), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n222_), .B(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G57gat), .B(G64gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT11), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(KEYINPUT68), .ZN(new_n231_));
  XOR2_X1   g030(.A(KEYINPUT67), .B(G71gat), .Z(new_n232_));
  INV_X1    g031(.A(G78gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT67), .B(G71gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(G78gat), .ZN(new_n236_));
  OAI211_X1 g035(.A(new_n234_), .B(new_n236_), .C1(KEYINPUT11), .C2(new_n229_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n231_), .B(new_n237_), .ZN(new_n238_));
  XOR2_X1   g037(.A(KEYINPUT10), .B(G99gat), .Z(new_n239_));
  XOR2_X1   g038(.A(KEYINPUT64), .B(G106gat), .Z(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  XOR2_X1   g040(.A(G85gat), .B(G92gat), .Z(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT9), .ZN(new_n243_));
  INV_X1    g042(.A(G85gat), .ZN(new_n244_));
  INV_X1    g043(.A(G92gat), .ZN(new_n245_));
  OR3_X1    g044(.A1(new_n244_), .A2(new_n245_), .A3(KEYINPUT9), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G99gat), .A2(G106gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(KEYINPUT6), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT6), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n249_), .A2(G99gat), .A3(G106gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n241_), .A2(new_n243_), .A3(new_n246_), .A4(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(G99gat), .ZN(new_n253_));
  INV_X1    g052(.A(G106gat), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n253_), .A2(new_n254_), .A3(KEYINPUT65), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT7), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT7), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n257_), .A2(new_n253_), .A3(new_n254_), .A4(KEYINPUT65), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n256_), .A2(new_n251_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT8), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n260_), .A2(KEYINPUT66), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  AND3_X1   g061(.A1(new_n259_), .A2(new_n242_), .A3(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n262_), .B1(new_n259_), .B2(new_n242_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n252_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT12), .B1(new_n238_), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n238_), .A2(new_n265_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G230gat), .A2(G233gat), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT69), .B1(new_n263_), .B2(new_n264_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n259_), .A2(new_n242_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(new_n261_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT69), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n259_), .A2(new_n242_), .A3(new_n262_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n272_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n270_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(new_n252_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n277_), .A2(KEYINPUT12), .A3(new_n238_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n268_), .A2(new_n269_), .A3(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n267_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n238_), .A2(new_n265_), .ZN(new_n281_));
  OAI211_X1 g080(.A(G230gat), .B(G233gat), .C1(new_n280_), .C2(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(KEYINPUT70), .B(KEYINPUT5), .Z(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT71), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G120gat), .B(G148gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G176gat), .B(G204gat), .ZN(new_n287_));
  XOR2_X1   g086(.A(new_n286_), .B(new_n287_), .Z(new_n288_));
  NAND3_X1  g087(.A1(new_n279_), .A2(new_n282_), .A3(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT72), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT72), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n279_), .A2(new_n282_), .A3(new_n291_), .A4(new_n288_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n288_), .B1(new_n279_), .B2(new_n282_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(KEYINPUT13), .B1(new_n293_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT13), .ZN(new_n298_));
  AOI211_X1 g097(.A(new_n298_), .B(new_n294_), .C1(new_n290_), .C2(new_n292_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n297_), .A2(new_n300_), .A3(KEYINPUT73), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT73), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n302_), .B1(new_n296_), .B2(new_n299_), .ZN(new_n303_));
  AND2_X1   g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(G134gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(G127gat), .ZN(new_n306_));
  INV_X1    g105(.A(G127gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(G134gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(G120gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(G113gat), .ZN(new_n311_));
  INV_X1    g110(.A(G113gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(G120gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n311_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n309_), .A2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G127gat), .B(G134gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G113gat), .B(G120gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n315_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT31), .ZN(new_n320_));
  OAI21_X1  g119(.A(KEYINPUT85), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n321_), .B1(new_n320_), .B2(new_n319_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G71gat), .B(G99gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(G43gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n322_), .B(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G227gat), .A2(G233gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(G15gat), .ZN(new_n327_));
  XOR2_X1   g126(.A(new_n327_), .B(KEYINPUT30), .Z(new_n328_));
  XNOR2_X1  g127(.A(new_n325_), .B(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G183gat), .A2(G190gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT23), .ZN(new_n331_));
  INV_X1    g130(.A(G190gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT81), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT81), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(G190gat), .ZN(new_n335_));
  INV_X1    g134(.A(G183gat), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n333_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n331_), .A2(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(G169gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(G169gat), .A2(G176gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(KEYINPUT83), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT83), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n345_), .B1(G169gat), .B2(G176gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT24), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n349_), .A2(KEYINPUT84), .A3(new_n331_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G169gat), .A2(G176gat), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n344_), .A2(KEYINPUT24), .A3(new_n346_), .A4(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT84), .ZN(new_n353_));
  AOI21_X1  g152(.A(KEYINPUT24), .B1(new_n344_), .B2(new_n346_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT23), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n330_), .B(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n353_), .B1(new_n354_), .B2(new_n356_), .ZN(new_n357_));
  AND3_X1   g156(.A1(new_n350_), .A2(new_n352_), .A3(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n336_), .A2(KEYINPUT25), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT25), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(G183gat), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT26), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n363_), .B1(new_n333_), .B2(new_n335_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n362_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT82), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  OAI211_X1 g167(.A(KEYINPUT82), .B(new_n362_), .C1(new_n364_), .C2(new_n365_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n342_), .B1(new_n358_), .B2(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT86), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  OR2_X1    g172(.A1(new_n329_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n329_), .A2(new_n373_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  XOR2_X1   g175(.A(G8gat), .B(G36gat), .Z(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT18), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G64gat), .B(G92gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G226gat), .A2(G233gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT19), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  XOR2_X1   g183(.A(G211gat), .B(G218gat), .Z(new_n385_));
  NOR2_X1   g184(.A1(G197gat), .A2(G204gat), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G197gat), .A2(G204gat), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n385_), .A2(KEYINPUT21), .A3(new_n387_), .A4(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n387_), .A2(KEYINPUT21), .A3(new_n388_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT21), .ZN(new_n391_));
  AND2_X1   g190(.A1(G197gat), .A2(G204gat), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n391_), .B1(new_n392_), .B2(new_n386_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G211gat), .B(G218gat), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n390_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n389_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT89), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n389_), .A2(new_n395_), .A3(KEYINPUT89), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n370_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n350_), .A2(new_n352_), .A3(new_n357_), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n400_), .B(new_n341_), .C1(new_n401_), .C2(new_n402_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(G183gat), .A2(G190gat), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n340_), .B1(new_n356_), .B2(new_n404_), .ZN(new_n405_));
  AND3_X1   g204(.A1(new_n351_), .A2(KEYINPUT91), .A3(KEYINPUT24), .ZN(new_n406_));
  AOI21_X1  g205(.A(KEYINPUT91), .B1(new_n351_), .B2(KEYINPUT24), .ZN(new_n407_));
  NOR3_X1   g206(.A1(new_n347_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n408_));
  AND2_X1   g207(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n359_), .B(new_n361_), .C1(new_n409_), .C2(new_n365_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n343_), .A2(new_n348_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n331_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n405_), .B1(new_n408_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(new_n396_), .ZN(new_n414_));
  AND2_X1   g213(.A1(new_n414_), .A2(KEYINPUT20), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n384_), .B1(new_n403_), .B2(new_n415_), .ZN(new_n416_));
  OAI211_X1 g215(.A(KEYINPUT20), .B(new_n384_), .C1(new_n413_), .C2(new_n396_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n341_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n400_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n417_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n381_), .B1(new_n416_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n417_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n422_), .B1(new_n371_), .B2(new_n400_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n414_), .A2(KEYINPUT20), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n424_), .B1(new_n371_), .B2(new_n400_), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n423_), .B(new_n380_), .C1(new_n425_), .C2(new_n384_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n421_), .A2(new_n426_), .ZN(new_n427_));
  OR2_X1    g226(.A1(new_n427_), .A2(KEYINPUT27), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G78gat), .B(G106gat), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT88), .ZN(new_n431_));
  INV_X1    g230(.A(G155gat), .ZN(new_n432_));
  INV_X1    g231(.A(G162gat), .ZN(new_n433_));
  AOI21_X1  g232(.A(KEYINPUT1), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G155gat), .A2(G162gat), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n431_), .B1(new_n434_), .B2(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(G155gat), .A2(G162gat), .ZN(new_n438_));
  OAI211_X1 g237(.A(KEYINPUT88), .B(new_n435_), .C1(new_n438_), .C2(KEYINPUT1), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n435_), .A2(KEYINPUT1), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n437_), .A2(new_n439_), .A3(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G141gat), .A2(G148gat), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT87), .ZN(new_n444_));
  NOR3_X1   g243(.A1(new_n444_), .A2(G141gat), .A3(G148gat), .ZN(new_n445_));
  INV_X1    g244(.A(G141gat), .ZN(new_n446_));
  INV_X1    g245(.A(G148gat), .ZN(new_n447_));
  AOI21_X1  g246(.A(KEYINPUT87), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n443_), .B1(new_n445_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n442_), .A2(new_n450_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(G141gat), .A2(G148gat), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT3), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT2), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n443_), .A2(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n454_), .A2(new_n456_), .A3(new_n457_), .A4(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n436_), .A2(new_n438_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n451_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT29), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n396_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n464_), .A2(G228gat), .A3(G233gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G228gat), .A2(G233gat), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n419_), .A2(new_n463_), .A3(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n430_), .B1(new_n465_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n465_), .A2(new_n430_), .A3(new_n467_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n462_), .A2(KEYINPUT29), .ZN(new_n472_));
  XOR2_X1   g271(.A(G22gat), .B(G50gat), .Z(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT28), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n472_), .B(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT90), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n475_), .B1(new_n468_), .B2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n471_), .A2(new_n477_), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n469_), .A2(new_n476_), .A3(new_n470_), .A4(new_n475_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT20), .B1(new_n413_), .B2(new_n396_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT98), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n481_), .B(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n371_), .A2(new_n400_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n383_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n425_), .A2(new_n384_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(new_n381_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n488_), .A2(KEYINPUT27), .A3(new_n426_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT92), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n435_), .B1(new_n438_), .B2(KEYINPUT1), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n440_), .B1(new_n491_), .B2(new_n431_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n449_), .B1(new_n492_), .B2(new_n439_), .ZN(new_n493_));
  AND2_X1   g292(.A1(new_n459_), .A2(new_n460_), .ZN(new_n494_));
  OAI211_X1 g293(.A(new_n490_), .B(new_n319_), .C1(new_n493_), .C2(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n309_), .A2(new_n314_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n316_), .A2(new_n317_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n490_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n315_), .A2(new_n318_), .A3(KEYINPUT92), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n451_), .A2(new_n498_), .A3(new_n499_), .A4(new_n461_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n495_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G225gat), .A2(G233gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G1gat), .B(G29gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G57gat), .B(G85gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n503_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n502_), .B(KEYINPUT93), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  AOI22_X1  g311(.A1(new_n442_), .A2(new_n450_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT4), .ZN(new_n514_));
  AND3_X1   g313(.A1(new_n315_), .A2(new_n318_), .A3(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(KEYINPUT94), .B1(new_n513_), .B2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT94), .ZN(new_n518_));
  OAI211_X1 g317(.A(new_n518_), .B(new_n515_), .C1(new_n493_), .C2(new_n494_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n512_), .B1(new_n517_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n501_), .A2(KEYINPUT4), .ZN(new_n521_));
  AND3_X1   g320(.A1(new_n520_), .A2(new_n521_), .A3(KEYINPUT95), .ZN(new_n522_));
  AOI21_X1  g321(.A(KEYINPUT95), .B1(new_n520_), .B2(new_n521_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n510_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n503_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT95), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n518_), .B1(new_n462_), .B2(new_n515_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n519_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n511_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n514_), .B1(new_n495_), .B2(new_n500_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n526_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n520_), .A2(new_n521_), .A3(KEYINPUT95), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n525_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n524_), .B1(new_n533_), .B2(new_n508_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n428_), .A2(new_n480_), .A3(new_n489_), .A4(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT97), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n509_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n537_), .B1(new_n538_), .B2(KEYINPUT33), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT33), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n524_), .A2(KEYINPUT97), .A3(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n538_), .A2(KEYINPUT33), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n508_), .B1(new_n501_), .B2(new_n511_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n502_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n543_), .B1(new_n544_), .B2(new_n530_), .ZN(new_n545_));
  AND3_X1   g344(.A1(new_n421_), .A2(new_n426_), .A3(new_n545_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n539_), .A2(new_n541_), .A3(new_n542_), .A4(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n487_), .A2(KEYINPUT32), .A3(new_n380_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n380_), .A2(KEYINPUT32), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n423_), .B(new_n549_), .C1(new_n425_), .C2(new_n384_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n534_), .A2(new_n548_), .A3(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n480_), .B1(new_n547_), .B2(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n536_), .B1(new_n552_), .B2(KEYINPUT99), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT99), .ZN(new_n554_));
  AOI211_X1 g353(.A(new_n554_), .B(new_n480_), .C1(new_n547_), .C2(new_n551_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n376_), .B1(new_n553_), .B2(new_n555_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n428_), .A2(new_n489_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n480_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n376_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(new_n535_), .ZN(new_n561_));
  OR2_X1    g360(.A1(new_n559_), .A2(new_n561_), .ZN(new_n562_));
  AOI211_X1 g361(.A(new_n228_), .B(new_n304_), .C1(new_n556_), .C2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G190gat), .B(G218gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G134gat), .B(G162gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n566_), .A2(KEYINPUT36), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n277_), .A2(new_n217_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT75), .ZN(new_n569_));
  INV_X1    g368(.A(new_n252_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n570_), .B1(new_n274_), .B2(new_n272_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(new_n211_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n573_));
  NAND2_X1  g372(.A1(G232gat), .A2(G233gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n568_), .A2(new_n569_), .A3(new_n572_), .A4(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(KEYINPUT35), .B1(new_n568_), .B2(new_n572_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n570_), .B1(new_n270_), .B2(new_n275_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n217_), .ZN(new_n580_));
  OAI211_X1 g379(.A(new_n569_), .B(new_n572_), .C1(new_n579_), .C2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(new_n575_), .ZN(new_n582_));
  OAI211_X1 g381(.A(new_n567_), .B(new_n577_), .C1(new_n578_), .C2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(KEYINPUT76), .ZN(new_n584_));
  AOI22_X1  g383(.A1(new_n277_), .A2(new_n217_), .B1(new_n211_), .B2(new_n571_), .ZN(new_n585_));
  OAI211_X1 g384(.A(new_n581_), .B(new_n575_), .C1(new_n585_), .C2(KEYINPUT35), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT76), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n586_), .A2(new_n587_), .A3(new_n567_), .A4(new_n577_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n586_), .A2(new_n577_), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n566_), .B(KEYINPUT36), .Z(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT77), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  AOI22_X1  g391(.A1(new_n584_), .A2(new_n588_), .B1(new_n589_), .B2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT78), .ZN(new_n594_));
  AND3_X1   g393(.A1(new_n593_), .A2(new_n594_), .A3(KEYINPUT37), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n594_), .A2(KEYINPUT37), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n594_), .A2(KEYINPUT37), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NOR3_X1   g397(.A1(new_n593_), .A2(new_n596_), .A3(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n595_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G231gat), .A2(G233gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n208_), .B(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n238_), .B(new_n602_), .ZN(new_n603_));
  XOR2_X1   g402(.A(G127gat), .B(G155gat), .Z(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT16), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G183gat), .B(G211gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT17), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n607_), .A2(new_n608_), .ZN(new_n610_));
  OR3_X1    g409(.A1(new_n603_), .A2(new_n609_), .A3(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n603_), .A2(new_n609_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n600_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT79), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n563_), .A2(new_n203_), .A3(new_n616_), .A4(new_n534_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT38), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n556_), .A2(new_n562_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n584_), .A2(new_n588_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n589_), .A2(new_n592_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  AND3_X1   g421(.A1(new_n619_), .A2(KEYINPUT100), .A3(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(KEYINPUT100), .B1(new_n619_), .B2(new_n622_), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n613_), .ZN(new_n626_));
  NOR3_X1   g425(.A1(new_n304_), .A2(new_n228_), .A3(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n625_), .A2(new_n534_), .A3(new_n627_), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n628_), .A2(KEYINPUT101), .A3(G1gat), .ZN(new_n629_));
  AOI21_X1  g428(.A(KEYINPUT101), .B1(new_n628_), .B2(G1gat), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n618_), .B1(new_n629_), .B2(new_n630_), .ZN(G1324gat));
  INV_X1    g430(.A(new_n557_), .ZN(new_n632_));
  OAI211_X1 g431(.A(new_n632_), .B(new_n627_), .C1(new_n623_), .C2(new_n624_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT39), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n633_), .A2(new_n634_), .A3(G8gat), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n634_), .B1(new_n633_), .B2(G8gat), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n563_), .A2(new_n616_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n632_), .A2(new_n204_), .ZN(new_n638_));
  OAI22_X1  g437(.A1(new_n635_), .A2(new_n636_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT40), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  OAI221_X1 g440(.A(KEYINPUT40), .B1(new_n637_), .B2(new_n638_), .C1(new_n635_), .C2(new_n636_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(G1325gat));
  OR3_X1    g442(.A1(new_n637_), .A2(G15gat), .A3(new_n376_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n625_), .A2(new_n560_), .A3(new_n627_), .ZN(new_n645_));
  AND3_X1   g444(.A1(new_n645_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n646_));
  AOI21_X1  g445(.A(KEYINPUT41), .B1(new_n645_), .B2(G15gat), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n644_), .B1(new_n646_), .B2(new_n647_), .ZN(G1326gat));
  OR3_X1    g447(.A1(new_n637_), .A2(G22gat), .A3(new_n558_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n625_), .A2(new_n480_), .A3(new_n627_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(G22gat), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n651_), .A2(KEYINPUT42), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n651_), .A2(KEYINPUT42), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n649_), .B1(new_n652_), .B2(new_n653_), .ZN(G1327gat));
  NOR3_X1   g453(.A1(new_n304_), .A2(new_n228_), .A3(new_n613_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT43), .ZN(new_n656_));
  INV_X1    g455(.A(new_n600_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n656_), .B1(new_n619_), .B2(new_n657_), .ZN(new_n658_));
  AOI211_X1 g457(.A(KEYINPUT43), .B(new_n600_), .C1(new_n556_), .C2(new_n562_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n655_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT44), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  OAI211_X1 g461(.A(KEYINPUT44), .B(new_n655_), .C1(new_n658_), .C2(new_n659_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n662_), .A2(new_n534_), .A3(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(G29gat), .ZN(new_n665_));
  INV_X1    g464(.A(new_n619_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n301_), .A2(new_n303_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n228_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n622_), .A2(new_n613_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n667_), .A2(new_n668_), .A3(new_n669_), .ZN(new_n670_));
  OAI21_X1  g469(.A(KEYINPUT102), .B1(new_n666_), .B2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n670_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT102), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n672_), .A2(new_n673_), .A3(new_n619_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n671_), .A2(new_n674_), .ZN(new_n675_));
  OR3_X1    g474(.A1(new_n675_), .A2(G29gat), .A3(new_n535_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n665_), .A2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(KEYINPUT103), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT103), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n665_), .A2(new_n679_), .A3(new_n676_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(G1328gat));
  NAND3_X1  g480(.A1(new_n662_), .A2(new_n632_), .A3(new_n663_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(G36gat), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n557_), .A2(G36gat), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n671_), .A2(new_n674_), .A3(new_n684_), .ZN(new_n685_));
  XOR2_X1   g484(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT105), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n685_), .B(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n683_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT46), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n683_), .A2(KEYINPUT46), .A3(new_n688_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(G1329gat));
  NAND4_X1  g492(.A1(new_n662_), .A2(G43gat), .A3(new_n560_), .A4(new_n663_), .ZN(new_n694_));
  INV_X1    g493(.A(G43gat), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n695_), .B1(new_n675_), .B2(new_n376_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n696_), .ZN(new_n697_));
  XOR2_X1   g496(.A(KEYINPUT106), .B(KEYINPUT47), .Z(new_n698_));
  XNOR2_X1  g497(.A(new_n697_), .B(new_n698_), .ZN(G1330gat));
  NAND4_X1  g498(.A1(new_n662_), .A2(G50gat), .A3(new_n480_), .A4(new_n663_), .ZN(new_n700_));
  INV_X1    g499(.A(G50gat), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n701_), .B1(new_n675_), .B2(new_n558_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n700_), .A2(new_n702_), .ZN(G1331gat));
  NAND2_X1  g502(.A1(new_n613_), .A2(new_n228_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n667_), .A2(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n625_), .A2(new_n534_), .A3(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(G57gat), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n616_), .A2(new_n304_), .ZN(new_n708_));
  AOI21_X1  g507(.A(KEYINPUT107), .B1(new_n619_), .B2(new_n228_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT107), .ZN(new_n710_));
  AOI211_X1 g509(.A(new_n710_), .B(new_n668_), .C1(new_n556_), .C2(new_n562_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n709_), .A2(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(KEYINPUT108), .B1(new_n708_), .B2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n619_), .A2(new_n228_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(new_n710_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n619_), .A2(KEYINPUT107), .A3(new_n228_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT108), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n717_), .A2(new_n616_), .A3(new_n718_), .A4(new_n304_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n713_), .A2(new_n719_), .ZN(new_n720_));
  OR2_X1    g519(.A1(new_n535_), .A2(G57gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n707_), .B1(new_n720_), .B2(new_n721_), .ZN(G1332gat));
  NOR2_X1   g521(.A1(new_n557_), .A2(G64gat), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n713_), .A2(new_n719_), .A3(new_n723_), .ZN(new_n724_));
  OAI211_X1 g523(.A(new_n632_), .B(new_n705_), .C1(new_n623_), .C2(new_n624_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n725_), .A2(KEYINPUT48), .A3(G64gat), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(G64gat), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT48), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n724_), .A2(new_n726_), .A3(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT109), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n724_), .A2(new_n729_), .A3(KEYINPUT109), .A4(new_n726_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1333gat));
  NAND3_X1  g533(.A1(new_n625_), .A2(new_n560_), .A3(new_n705_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(G71gat), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n736_), .A2(KEYINPUT49), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n736_), .A2(KEYINPUT49), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n376_), .A2(G71gat), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT110), .Z(new_n740_));
  OAI22_X1  g539(.A1(new_n737_), .A2(new_n738_), .B1(new_n720_), .B2(new_n740_), .ZN(G1334gat));
  NAND3_X1  g540(.A1(new_n625_), .A2(new_n480_), .A3(new_n705_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(G78gat), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n743_), .A2(KEYINPUT50), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n743_), .A2(KEYINPUT50), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n480_), .A2(new_n233_), .ZN(new_n746_));
  OAI22_X1  g545(.A1(new_n744_), .A2(new_n745_), .B1(new_n720_), .B2(new_n746_), .ZN(G1335gat));
  OR2_X1    g546(.A1(new_n658_), .A2(new_n659_), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n301_), .A2(new_n303_), .A3(new_n228_), .A4(new_n626_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT111), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n748_), .A2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n534_), .A2(G85gat), .ZN(new_n752_));
  XOR2_X1   g551(.A(new_n752_), .B(KEYINPUT112), .Z(new_n753_));
  NOR3_X1   g552(.A1(new_n667_), .A2(new_n622_), .A3(new_n613_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n717_), .A2(new_n534_), .A3(new_n754_), .ZN(new_n755_));
  AOI22_X1  g554(.A1(new_n751_), .A2(new_n753_), .B1(new_n244_), .B2(new_n755_), .ZN(G1336gat));
  NAND4_X1  g555(.A1(new_n748_), .A2(G92gat), .A3(new_n632_), .A4(new_n750_), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n632_), .B(new_n754_), .C1(new_n709_), .C2(new_n711_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT113), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n758_), .A2(new_n759_), .A3(new_n245_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n758_), .B2(new_n245_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n757_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT114), .ZN(G1337gat));
  AND2_X1   g562(.A1(new_n560_), .A2(new_n239_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n717_), .A2(KEYINPUT116), .A3(new_n754_), .A4(new_n764_), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n754_), .B(new_n764_), .C1(new_n709_), .C2(new_n711_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT116), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n765_), .A2(new_n768_), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n750_), .B(new_n560_), .C1(new_n658_), .C2(new_n659_), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n770_), .A2(KEYINPUT115), .A3(G99gat), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT115), .B1(new_n770_), .B2(G99gat), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n769_), .B(KEYINPUT117), .C1(new_n771_), .C2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT51), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT117), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n775_), .B1(new_n765_), .B2(new_n768_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n776_), .B(new_n777_), .C1(new_n772_), .C2(new_n771_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n774_), .A2(new_n778_), .ZN(G1338gat));
  NAND4_X1  g578(.A1(new_n717_), .A2(new_n480_), .A3(new_n240_), .A4(new_n754_), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n750_), .B(new_n480_), .C1(new_n658_), .C2(new_n659_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n782_));
  AND3_X1   g581(.A1(new_n781_), .A2(new_n782_), .A3(G106gat), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n782_), .B1(new_n781_), .B2(G106gat), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n780_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT53), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT53), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n780_), .B(new_n787_), .C1(new_n783_), .C2(new_n784_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n788_), .ZN(G1339gat));
  NAND2_X1  g588(.A1(new_n560_), .A2(new_n534_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n559_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n269_), .B1(new_n268_), .B2(new_n278_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n279_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n268_), .A2(new_n278_), .A3(KEYINPUT55), .A4(new_n269_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n288_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT56), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n797_), .A2(KEYINPUT56), .A3(new_n798_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n212_), .A2(new_n213_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n218_), .A2(new_n220_), .A3(new_n214_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n804_), .A2(new_n805_), .A3(new_n226_), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n806_), .B(KEYINPUT118), .ZN(new_n807_));
  INV_X1    g606(.A(new_n222_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n807_), .B1(new_n225_), .B2(new_n808_), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n809_), .A2(new_n293_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n803_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT58), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT56), .B1(new_n797_), .B2(new_n798_), .ZN(new_n814_));
  AOI211_X1 g613(.A(new_n800_), .B(new_n288_), .C1(new_n795_), .C2(new_n796_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n810_), .B(KEYINPUT58), .C1(new_n814_), .C2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT120), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n803_), .A2(KEYINPUT120), .A3(KEYINPUT58), .A4(new_n810_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n657_), .A2(new_n813_), .A3(new_n818_), .A4(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n293_), .A2(new_n668_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n821_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n293_), .A2(new_n295_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n809_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n622_), .B1(new_n822_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT57), .ZN(new_n827_));
  NOR3_X1   g626(.A1(new_n826_), .A2(KEYINPUT121), .A3(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT121), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n668_), .B(new_n293_), .C1(new_n814_), .C2(new_n815_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n593_), .B1(new_n830_), .B2(new_n824_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n829_), .B1(new_n831_), .B2(KEYINPUT57), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n820_), .B1(new_n828_), .B2(new_n832_), .ZN(new_n833_));
  OR3_X1    g632(.A1(new_n831_), .A2(KEYINPUT119), .A3(KEYINPUT57), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n826_), .A2(new_n827_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT119), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n626_), .B1(new_n833_), .B2(new_n837_), .ZN(new_n838_));
  NOR3_X1   g637(.A1(new_n296_), .A2(new_n299_), .A3(new_n704_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n600_), .A2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT54), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n840_), .B(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n792_), .B1(new_n838_), .B2(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n844_), .A2(new_n312_), .A3(new_n668_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(KEYINPUT59), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT59), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n820_), .B(new_n835_), .C1(new_n828_), .C2(new_n832_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n842_), .B1(new_n848_), .B2(new_n626_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n791_), .B(KEYINPUT122), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n847_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n228_), .B1(new_n846_), .B2(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n845_), .B1(new_n852_), .B2(new_n312_), .ZN(G1340gat));
  AOI21_X1  g652(.A(new_n667_), .B1(new_n846_), .B2(new_n851_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n667_), .A2(KEYINPUT60), .ZN(new_n855_));
  MUX2_X1   g654(.A(KEYINPUT60), .B(new_n855_), .S(new_n310_), .Z(new_n856_));
  AND3_X1   g655(.A1(new_n844_), .A2(KEYINPUT123), .A3(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(KEYINPUT123), .B1(new_n844_), .B2(new_n856_), .ZN(new_n858_));
  OAI22_X1  g657(.A1(new_n854_), .A2(new_n310_), .B1(new_n857_), .B2(new_n858_), .ZN(G1341gat));
  NAND3_X1  g658(.A1(new_n844_), .A2(new_n307_), .A3(new_n613_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n626_), .B1(new_n846_), .B2(new_n851_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(new_n861_), .B2(new_n307_), .ZN(G1342gat));
  NAND3_X1  g661(.A1(new_n844_), .A2(new_n305_), .A3(new_n593_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n600_), .B1(new_n846_), .B2(new_n851_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n864_), .B2(new_n305_), .ZN(G1343gat));
  NAND2_X1  g664(.A1(new_n838_), .A2(new_n843_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n632_), .A2(new_n558_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n867_), .A2(new_n534_), .A3(new_n376_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n866_), .A2(new_n668_), .A3(new_n869_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g670(.A1(new_n866_), .A2(new_n304_), .A3(new_n869_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g672(.A1(new_n866_), .A2(new_n613_), .A3(new_n869_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(KEYINPUT61), .B(G155gat), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n874_), .B(new_n875_), .ZN(G1346gat));
  NAND2_X1  g675(.A1(new_n866_), .A2(new_n869_), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n877_), .A2(new_n433_), .A3(new_n600_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT124), .ZN(new_n879_));
  AOI211_X1 g678(.A(new_n622_), .B(new_n868_), .C1(new_n838_), .C2(new_n843_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n879_), .B1(new_n880_), .B2(G162gat), .ZN(new_n881_));
  OAI211_X1 g680(.A(KEYINPUT124), .B(new_n433_), .C1(new_n877_), .C2(new_n622_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n878_), .B1(new_n881_), .B2(new_n882_), .ZN(G1347gat));
  INV_X1    g682(.A(new_n849_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT62), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n561_), .A2(new_n557_), .A3(new_n480_), .ZN(new_n886_));
  NAND4_X1  g685(.A1(new_n884_), .A2(new_n885_), .A3(new_n668_), .A4(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n886_), .ZN(new_n888_));
  NOR4_X1   g687(.A1(new_n849_), .A2(KEYINPUT22), .A3(new_n228_), .A4(new_n888_), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n887_), .B(G169gat), .C1(new_n889_), .C2(new_n885_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n849_), .A2(new_n888_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT22), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n891_), .A2(new_n892_), .A3(new_n668_), .ZN(new_n893_));
  INV_X1    g692(.A(G169gat), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n893_), .A2(KEYINPUT62), .A3(new_n894_), .ZN(new_n895_));
  AND2_X1   g694(.A1(new_n890_), .A2(new_n895_), .ZN(G1348gat));
  AOI21_X1  g695(.A(G176gat), .B1(new_n891_), .B2(new_n304_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n888_), .B1(new_n838_), .B2(new_n843_), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n304_), .A2(G176gat), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n897_), .B1(new_n898_), .B2(new_n899_), .ZN(G1349gat));
  AOI21_X1  g699(.A(G183gat), .B1(new_n898_), .B2(new_n613_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n626_), .A2(new_n362_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n901_), .B1(new_n891_), .B2(new_n902_), .ZN(G1350gat));
  OAI211_X1 g702(.A(new_n891_), .B(new_n593_), .C1(new_n365_), .C2(new_n409_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT125), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n891_), .A2(new_n657_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n905_), .B1(new_n906_), .B2(G190gat), .ZN(new_n907_));
  AOI211_X1 g706(.A(KEYINPUT125), .B(new_n332_), .C1(new_n891_), .C2(new_n657_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n904_), .B1(new_n907_), .B2(new_n908_), .ZN(G1351gat));
  NOR3_X1   g708(.A1(new_n560_), .A2(new_n534_), .A3(new_n558_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT126), .ZN(new_n911_));
  AND2_X1   g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n910_), .A2(new_n911_), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n912_), .A2(new_n913_), .A3(new_n557_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n866_), .A2(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  AOI21_X1  g715(.A(G197gat), .B1(new_n916_), .B2(new_n668_), .ZN(new_n917_));
  INV_X1    g716(.A(G197gat), .ZN(new_n918_));
  NOR3_X1   g717(.A1(new_n915_), .A2(new_n918_), .A3(new_n228_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n917_), .A2(new_n919_), .ZN(G1352gat));
  XNOR2_X1  g719(.A(KEYINPUT127), .B(G204gat), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n921_), .B1(new_n916_), .B2(new_n304_), .ZN(new_n922_));
  AND4_X1   g721(.A1(new_n304_), .A2(new_n866_), .A3(new_n914_), .A4(new_n921_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n922_), .A2(new_n923_), .ZN(G1353gat));
  XNOR2_X1  g723(.A(KEYINPUT63), .B(G211gat), .ZN(new_n925_));
  NOR3_X1   g724(.A1(new_n915_), .A2(new_n626_), .A3(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n916_), .A2(new_n613_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n926_), .B1(new_n927_), .B2(new_n928_), .ZN(G1354gat));
  OR3_X1    g728(.A1(new_n915_), .A2(G218gat), .A3(new_n622_), .ZN(new_n930_));
  OAI21_X1  g729(.A(G218gat), .B1(new_n915_), .B2(new_n600_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(G1355gat));
endmodule


