//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 1 0 1 0 1 1 0 1 1 0 1 0 0 1 0 1 0 1 0 0 1 1 0 1 0 1 0 1 1 1 1 1 1 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 1 1 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n636_, new_n637_, new_n638_, new_n640_,
    new_n641_, new_n642_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n657_, new_n658_, new_n659_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n683_, new_n684_, new_n685_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n834_, new_n835_, new_n836_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n843_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n882_, new_n883_, new_n885_, new_n886_, new_n888_, new_n889_,
    new_n890_, new_n892_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_;
  INV_X1    g000(.A(KEYINPUT6), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT65), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT65), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT6), .ZN(new_n205_));
  AND2_X1   g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  AND3_X1   g005(.A1(new_n203_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n206_), .B1(new_n203_), .B2(new_n205_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT7), .ZN(new_n209_));
  INV_X1    g008(.A(G99gat), .ZN(new_n210_));
  INV_X1    g009(.A(G106gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n209_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NOR3_X1   g013(.A1(new_n207_), .A2(new_n208_), .A3(new_n214_), .ZN(new_n215_));
  XOR2_X1   g014(.A(G85gat), .B(G92gat), .Z(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT67), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT8), .B1(new_n215_), .B2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n206_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n204_), .A2(KEYINPUT6), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n202_), .A2(KEYINPUT65), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n219_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n203_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n222_), .A2(new_n223_), .A3(new_n213_), .A4(new_n212_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n217_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT8), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n224_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n218_), .A2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT64), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT64), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n231_), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(KEYINPUT9), .A2(G85gat), .ZN(new_n233_));
  INV_X1    g032(.A(G92gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  OR2_X1    g034(.A1(KEYINPUT9), .A2(G85gat), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n230_), .A2(new_n232_), .A3(new_n235_), .A4(new_n236_), .ZN(new_n237_));
  OR2_X1    g036(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n238_), .A2(new_n211_), .A3(new_n239_), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n237_), .A2(new_n222_), .A3(new_n223_), .A4(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT66), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n207_), .A2(new_n208_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n243_), .A2(new_n244_), .A3(new_n237_), .A4(new_n240_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n242_), .A2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G57gat), .B(G64gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(KEYINPUT11), .ZN(new_n248_));
  XOR2_X1   g047(.A(G71gat), .B(G78gat), .Z(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n247_), .A2(KEYINPUT11), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  OR2_X1    g051(.A1(new_n248_), .A2(new_n249_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n228_), .A2(new_n246_), .A3(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT12), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n224_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n226_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n241_), .B(new_n244_), .ZN(new_n260_));
  OAI211_X1 g059(.A(new_n253_), .B(new_n252_), .C1(new_n259_), .C2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n256_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT68), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n263_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n228_), .A2(KEYINPUT68), .A3(new_n246_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n252_), .A2(KEYINPUT12), .A3(new_n253_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n264_), .A2(new_n265_), .A3(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G230gat), .A2(G233gat), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n262_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n261_), .A2(new_n255_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n269_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n270_), .A2(new_n273_), .ZN(new_n274_));
  XOR2_X1   g073(.A(G120gat), .B(G148gat), .Z(new_n275_));
  XNOR2_X1  g074(.A(G176gat), .B(G204gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n278_));
  XOR2_X1   g077(.A(new_n277_), .B(new_n278_), .Z(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT70), .B1(new_n274_), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n270_), .A2(new_n282_), .A3(new_n273_), .A4(new_n279_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n281_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n274_), .A2(new_n280_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT13), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n284_), .A2(KEYINPUT13), .A3(new_n285_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G29gat), .B(G36gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G43gat), .B(G50gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT72), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G15gat), .B(G22gat), .ZN(new_n296_));
  INV_X1    g095(.A(G1gat), .ZN(new_n297_));
  INV_X1    g096(.A(G8gat), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT14), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n296_), .A2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G1gat), .B(G8gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  OR2_X1    g101(.A1(new_n295_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G229gat), .A2(G233gat), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  XOR2_X1   g104(.A(KEYINPUT71), .B(KEYINPUT15), .Z(new_n306_));
  XNOR2_X1  g105(.A(new_n293_), .B(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(new_n302_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n295_), .B(new_n302_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n304_), .ZN(new_n310_));
  AOI22_X1  g109(.A1(new_n305_), .A2(new_n308_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G113gat), .B(G141gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G169gat), .B(G197gat), .ZN(new_n313_));
  XOR2_X1   g112(.A(new_n312_), .B(new_n313_), .Z(new_n314_));
  OR2_X1    g113(.A1(new_n311_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n311_), .A2(new_n314_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n290_), .A2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n254_), .B(new_n302_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G231gat), .A2(G233gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT17), .ZN(new_n323_));
  XOR2_X1   g122(.A(G127gat), .B(G155gat), .Z(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT16), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G183gat), .B(G211gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  OR3_X1    g126(.A1(new_n322_), .A2(new_n323_), .A3(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(KEYINPUT17), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n322_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n319_), .A2(new_n332_), .ZN(new_n333_));
  OR2_X1    g132(.A1(new_n333_), .A2(KEYINPUT91), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G190gat), .B(G218gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G134gat), .B(G162gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  XOR2_X1   g136(.A(new_n337_), .B(KEYINPUT36), .Z(new_n338_));
  NOR2_X1   g137(.A1(new_n259_), .A2(new_n260_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT35), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G232gat), .A2(G233gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT34), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  AOI22_X1  g142(.A1(new_n339_), .A2(new_n293_), .B1(new_n340_), .B2(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n264_), .A2(new_n307_), .A3(new_n265_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n343_), .A2(new_n340_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n346_), .A2(new_n347_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n338_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n350_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n337_), .A2(KEYINPUT36), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n352_), .A2(new_n353_), .A3(new_n348_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n351_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G71gat), .B(G99gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(G43gat), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n360_), .B1(G169gat), .B2(G176gat), .ZN(new_n361_));
  OR2_X1    g160(.A1(new_n361_), .A2(KEYINPUT74), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G183gat), .A2(G190gat), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT23), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  NOR3_X1   g164(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT25), .B(G183gat), .ZN(new_n368_));
  INV_X1    g167(.A(G190gat), .ZN(new_n369_));
  OAI21_X1  g168(.A(KEYINPUT26), .B1(new_n369_), .B2(KEYINPUT73), .ZN(new_n370_));
  OR2_X1    g169(.A1(new_n369_), .A2(KEYINPUT26), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n368_), .B(new_n370_), .C1(new_n371_), .C2(KEYINPUT73), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n361_), .A2(KEYINPUT74), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n362_), .A2(new_n367_), .A3(new_n372_), .A4(new_n373_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(G183gat), .A2(G190gat), .ZN(new_n375_));
  OR2_X1    g174(.A1(new_n365_), .A2(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(G169gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n374_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G227gat), .A2(G233gat), .ZN(new_n381_));
  XOR2_X1   g180(.A(new_n381_), .B(G15gat), .Z(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT30), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n380_), .B(new_n383_), .ZN(new_n384_));
  XOR2_X1   g183(.A(G127gat), .B(G134gat), .Z(new_n385_));
  XOR2_X1   g184(.A(G113gat), .B(G120gat), .Z(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  OR2_X1    g187(.A1(new_n388_), .A2(KEYINPUT31), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(KEYINPUT31), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n389_), .A2(KEYINPUT75), .A3(new_n390_), .ZN(new_n391_));
  AND2_X1   g190(.A1(new_n384_), .A2(new_n391_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n384_), .A2(new_n391_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n359_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  OR2_X1    g193(.A1(new_n384_), .A2(new_n391_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n384_), .A2(new_n391_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n395_), .A2(new_n358_), .A3(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n394_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(G197gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(G204gat), .ZN(new_n401_));
  INV_X1    g200(.A(G204gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(G197gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n404_), .A2(KEYINPUT21), .ZN(new_n405_));
  XOR2_X1   g204(.A(G211gat), .B(G218gat), .Z(new_n406_));
  NOR2_X1   g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n404_), .A2(KEYINPUT79), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT79), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT21), .B1(new_n401_), .B2(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n407_), .B1(new_n408_), .B2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n406_), .A2(KEYINPUT21), .A3(new_n404_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  OR2_X1    g212(.A1(G141gat), .A2(G148gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G141gat), .A2(G148gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(G155gat), .A2(G162gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G155gat), .A2(G162gat), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n417_), .B1(KEYINPUT1), .B2(new_n418_), .ZN(new_n419_));
  OR2_X1    g218(.A1(new_n418_), .A2(KEYINPUT1), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n416_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT76), .ZN(new_n422_));
  AOI21_X1  g221(.A(KEYINPUT3), .B1(new_n414_), .B2(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n423_), .B1(new_n422_), .B2(new_n414_), .ZN(new_n424_));
  OAI21_X1  g223(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT77), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n415_), .B(KEYINPUT2), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n424_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n418_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n429_), .A2(new_n417_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n421_), .B1(new_n428_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT29), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n413_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n433_), .A2(G228gat), .A3(G233gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G228gat), .A2(G233gat), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n413_), .B(new_n435_), .C1(new_n431_), .C2(new_n432_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G78gat), .B(G106gat), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n434_), .A2(new_n436_), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT80), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n431_), .A2(new_n432_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(KEYINPUT78), .B(KEYINPUT28), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G22gat), .B(G50gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n442_), .B(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n441_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n434_), .A2(new_n436_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(new_n437_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(new_n439_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n447_), .A2(new_n450_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n449_), .A2(KEYINPUT80), .A3(new_n439_), .A4(new_n446_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n380_), .A2(new_n413_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT82), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n380_), .A2(new_n413_), .A3(KEYINPUT82), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(KEYINPUT26), .B(G190gat), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n361_), .B1(new_n368_), .B2(new_n459_), .ZN(new_n460_));
  AOI22_X1  g259(.A1(new_n376_), .A2(new_n378_), .B1(new_n460_), .B2(new_n367_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n461_), .A2(KEYINPUT83), .A3(new_n411_), .A4(new_n412_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(KEYINPUT81), .B(KEYINPUT19), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G226gat), .A2(G233gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT20), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n461_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT83), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n466_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n458_), .A2(new_n462_), .A3(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G64gat), .B(G92gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT85), .ZN(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT84), .B(KEYINPUT18), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G8gat), .B(G36gat), .ZN(new_n475_));
  XOR2_X1   g274(.A(new_n474_), .B(new_n475_), .Z(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  OR2_X1    g276(.A1(new_n380_), .A2(new_n413_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT20), .ZN(new_n479_));
  INV_X1    g278(.A(new_n461_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n479_), .B1(new_n480_), .B2(new_n413_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n478_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n465_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  AND3_X1   g283(.A1(new_n470_), .A2(new_n477_), .A3(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n477_), .B1(new_n470_), .B2(new_n484_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G225gat), .A2(G233gat), .ZN(new_n488_));
  XOR2_X1   g287(.A(new_n488_), .B(KEYINPUT87), .Z(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n388_), .A2(KEYINPUT86), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT86), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n387_), .A2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n491_), .A2(new_n431_), .A3(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NOR3_X1   g294(.A1(new_n431_), .A2(KEYINPUT86), .A3(new_n388_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n490_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G1gat), .B(G29gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G57gat), .B(G85gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(KEYINPUT88), .B(KEYINPUT0), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT4), .ZN(new_n503_));
  INV_X1    g302(.A(new_n431_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n504_), .A2(new_n492_), .A3(new_n387_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n503_), .B1(new_n505_), .B2(new_n494_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n504_), .A2(new_n503_), .A3(new_n388_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(new_n489_), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n497_), .B(new_n502_), .C1(new_n506_), .C2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT33), .ZN(new_n510_));
  OR2_X1    g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n509_), .A2(new_n510_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n489_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n502_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n507_), .A2(new_n490_), .ZN(new_n515_));
  OAI211_X1 g314(.A(new_n513_), .B(new_n514_), .C1(new_n506_), .C2(new_n515_), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n487_), .A2(new_n511_), .A3(new_n512_), .A4(new_n516_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n497_), .B1(new_n506_), .B2(new_n508_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(new_n514_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(new_n509_), .ZN(new_n520_));
  AND2_X1   g319(.A1(new_n477_), .A2(KEYINPUT32), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n478_), .A2(new_n481_), .A3(new_n465_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT89), .B(KEYINPUT20), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n467_), .A2(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n525_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n522_), .B1(new_n526_), .B2(new_n465_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n521_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n470_), .A2(new_n484_), .ZN(new_n529_));
  OAI211_X1 g328(.A(new_n520_), .B(new_n528_), .C1(new_n521_), .C2(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n453_), .B1(new_n517_), .B2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n520_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT27), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n533_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n527_), .A2(new_n476_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n470_), .A2(new_n477_), .A3(new_n484_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n535_), .A2(KEYINPUT27), .A3(new_n536_), .ZN(new_n537_));
  AND4_X1   g336(.A1(new_n532_), .A2(new_n453_), .A3(new_n534_), .A4(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n399_), .B1(new_n531_), .B2(new_n538_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n534_), .A2(new_n452_), .A3(new_n537_), .A4(new_n451_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n532_), .A2(new_n398_), .ZN(new_n541_));
  OAI21_X1  g340(.A(KEYINPUT90), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n529_), .A2(new_n476_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(new_n536_), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n469_), .A2(new_n462_), .ZN(new_n545_));
  AOI22_X1  g344(.A1(new_n545_), .A2(new_n458_), .B1(new_n483_), .B2(new_n482_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n533_), .B1(new_n546_), .B2(new_n477_), .ZN(new_n547_));
  AOI22_X1  g346(.A1(new_n544_), .A2(new_n533_), .B1(new_n547_), .B2(new_n535_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT90), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n399_), .A2(new_n520_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n453_), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n548_), .A2(new_n549_), .A3(new_n550_), .A4(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n542_), .A2(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n356_), .B1(new_n539_), .B2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n333_), .A2(KEYINPUT91), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n334_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT92), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  OAI21_X1  g357(.A(G1gat), .B1(new_n558_), .B2(new_n532_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n539_), .A2(new_n553_), .ZN(new_n560_));
  AND2_X1   g359(.A1(new_n560_), .A2(new_n319_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n355_), .A2(KEYINPUT37), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT37), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n351_), .A2(new_n354_), .A3(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n566_), .A2(new_n331_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n561_), .A2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n568_), .A2(new_n297_), .A3(new_n520_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT38), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n559_), .A2(new_n570_), .ZN(G1324gat));
  INV_X1    g370(.A(new_n568_), .ZN(new_n572_));
  NOR3_X1   g371(.A1(new_n572_), .A2(G8gat), .A3(new_n548_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n548_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n334_), .A2(new_n574_), .A3(new_n554_), .A4(new_n555_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT93), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(G8gat), .B1(new_n575_), .B2(new_n576_), .ZN(new_n579_));
  OAI21_X1  g378(.A(KEYINPUT39), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n575_), .A2(new_n576_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT39), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n581_), .A2(new_n582_), .A3(G8gat), .A4(new_n577_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n573_), .B1(new_n580_), .B2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(KEYINPUT94), .B(KEYINPUT40), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n585_), .ZN(new_n587_));
  AOI211_X1 g386(.A(new_n573_), .B(new_n587_), .C1(new_n580_), .C2(new_n583_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n586_), .A2(new_n588_), .ZN(G1325gat));
  OR3_X1    g388(.A1(new_n572_), .A2(G15gat), .A3(new_n399_), .ZN(new_n590_));
  OAI21_X1  g389(.A(G15gat), .B1(new_n558_), .B2(new_n399_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT41), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n591_), .A2(new_n592_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n590_), .B1(new_n593_), .B2(new_n594_), .ZN(G1326gat));
  OAI21_X1  g394(.A(G22gat), .B1(new_n558_), .B2(new_n551_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n596_), .A2(KEYINPUT42), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(KEYINPUT42), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n551_), .A2(G22gat), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n599_), .B(KEYINPUT95), .Z(new_n600_));
  OAI22_X1  g399(.A1(new_n597_), .A2(new_n598_), .B1(new_n572_), .B2(new_n600_), .ZN(G1327gat));
  NOR3_X1   g400(.A1(new_n290_), .A2(new_n318_), .A3(new_n332_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT96), .ZN(new_n603_));
  AOI221_X4 g402(.A(new_n565_), .B1(new_n603_), .B2(KEYINPUT43), .C1(new_n539_), .C2(new_n553_), .ZN(new_n604_));
  OAI21_X1  g403(.A(KEYINPUT43), .B1(new_n565_), .B2(new_n603_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n605_), .B1(new_n560_), .B2(new_n566_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n602_), .B1(new_n604_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT44), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  OAI211_X1 g408(.A(new_n602_), .B(KEYINPUT44), .C1(new_n604_), .C2(new_n606_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  OAI21_X1  g410(.A(G29gat), .B1(new_n611_), .B2(new_n532_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n332_), .A2(new_n355_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT97), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n561_), .A2(new_n614_), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n532_), .A2(G29gat), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n612_), .B1(new_n615_), .B2(new_n616_), .ZN(G1328gat));
  XNOR2_X1  g416(.A(new_n574_), .B(KEYINPUT99), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n619_), .A2(G36gat), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  OR3_X1    g420(.A1(new_n615_), .A2(new_n621_), .A3(KEYINPUT100), .ZN(new_n622_));
  OAI21_X1  g421(.A(KEYINPUT100), .B1(new_n615_), .B2(new_n621_), .ZN(new_n623_));
  AND3_X1   g422(.A1(new_n622_), .A2(KEYINPUT45), .A3(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(KEYINPUT45), .B1(new_n622_), .B2(new_n623_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n609_), .A2(new_n574_), .A3(new_n610_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT98), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  OAI21_X1  g428(.A(G36gat), .B1(new_n627_), .B2(new_n628_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n626_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT46), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  OAI211_X1 g432(.A(new_n626_), .B(KEYINPUT46), .C1(new_n629_), .C2(new_n630_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(G1329gat));
  NAND2_X1  g434(.A1(new_n398_), .A2(G43gat), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n615_), .A2(new_n399_), .ZN(new_n637_));
  OAI22_X1  g436(.A1(new_n611_), .A2(new_n636_), .B1(G43gat), .B2(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g438(.A(G50gat), .B1(new_n611_), .B2(new_n551_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n551_), .A2(G50gat), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n641_), .B(KEYINPUT101), .Z(new_n642_));
  OAI21_X1  g441(.A(new_n640_), .B1(new_n615_), .B2(new_n642_), .ZN(G1331gat));
  INV_X1    g442(.A(G57gat), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n567_), .A2(new_n290_), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n645_), .A2(KEYINPUT102), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n317_), .B1(new_n539_), .B2(new_n553_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(KEYINPUT102), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n646_), .A2(new_n647_), .A3(new_n648_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n644_), .B1(new_n649_), .B2(new_n532_), .ZN(new_n650_));
  XOR2_X1   g449(.A(new_n650_), .B(KEYINPUT103), .Z(new_n651_));
  NOR2_X1   g450(.A1(new_n331_), .A2(new_n317_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n290_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n554_), .A2(new_n653_), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n654_), .A2(new_n644_), .A3(new_n532_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n651_), .A2(new_n655_), .ZN(G1332gat));
  OAI21_X1  g455(.A(G64gat), .B1(new_n654_), .B2(new_n619_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT48), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n619_), .A2(G64gat), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n658_), .B1(new_n649_), .B2(new_n659_), .ZN(G1333gat));
  OAI21_X1  g459(.A(G71gat), .B1(new_n654_), .B2(new_n399_), .ZN(new_n661_));
  XOR2_X1   g460(.A(KEYINPUT104), .B(KEYINPUT49), .Z(new_n662_));
  XNOR2_X1  g461(.A(new_n661_), .B(new_n662_), .ZN(new_n663_));
  OR2_X1    g462(.A1(new_n399_), .A2(G71gat), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n663_), .B1(new_n649_), .B2(new_n664_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT105), .ZN(G1334gat));
  OAI21_X1  g465(.A(G78gat), .B1(new_n654_), .B2(new_n551_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(KEYINPUT106), .B(KEYINPUT50), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n667_), .B(new_n668_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n551_), .A2(G78gat), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT107), .Z(new_n671_));
  OAI21_X1  g470(.A(new_n669_), .B1(new_n649_), .B2(new_n671_), .ZN(G1335gat));
  AND2_X1   g471(.A1(new_n614_), .A2(new_n290_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(new_n647_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n674_), .A2(G85gat), .A3(new_n532_), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n604_), .A2(new_n606_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n290_), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n677_), .A2(new_n317_), .A3(new_n332_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n676_), .A2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(new_n520_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n675_), .B1(new_n680_), .B2(G85gat), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT108), .ZN(G1336gat));
  OAI21_X1  g481(.A(new_n234_), .B1(new_n674_), .B2(new_n548_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT109), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n619_), .A2(new_n234_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n679_), .B2(new_n685_), .ZN(G1337gat));
  INV_X1    g485(.A(KEYINPUT113), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n398_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n674_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT112), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT51), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n691_), .A2(new_n692_), .A3(KEYINPUT111), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n398_), .B(new_n678_), .C1(new_n604_), .C2(new_n606_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT110), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n694_), .A2(new_n695_), .A3(G99gat), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n695_), .B1(new_n694_), .B2(G99gat), .ZN(new_n698_));
  OAI211_X1 g497(.A(new_n690_), .B(new_n693_), .C1(new_n697_), .C2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n694_), .A2(G99gat), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(KEYINPUT110), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n689_), .B1(new_n701_), .B2(new_n696_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT111), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n699_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(KEYINPUT51), .B1(new_n702_), .B2(KEYINPUT112), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n687_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n690_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n692_), .B1(new_n707_), .B2(new_n691_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(KEYINPUT111), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n708_), .A2(KEYINPUT113), .A3(new_n699_), .A4(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n706_), .A2(new_n710_), .ZN(G1338gat));
  NAND4_X1  g510(.A1(new_n673_), .A2(new_n211_), .A3(new_n453_), .A4(new_n647_), .ZN(new_n712_));
  OAI211_X1 g511(.A(new_n453_), .B(new_n678_), .C1(new_n604_), .C2(new_n606_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(G106gat), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(KEYINPUT114), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT52), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT114), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n713_), .A2(new_n717_), .A3(G106gat), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n715_), .A2(new_n716_), .A3(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n716_), .B1(new_n715_), .B2(new_n718_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n712_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(KEYINPUT53), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT53), .ZN(new_n723_));
  OAI211_X1 g522(.A(new_n723_), .B(new_n712_), .C1(new_n719_), .C2(new_n720_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n722_), .A2(new_n724_), .ZN(G1339gat));
  NAND3_X1  g524(.A1(new_n288_), .A2(new_n289_), .A3(new_n652_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT115), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n565_), .B1(new_n726_), .B2(KEYINPUT115), .ZN(new_n729_));
  OAI21_X1  g528(.A(KEYINPUT54), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  OR2_X1    g529(.A1(new_n726_), .A2(KEYINPUT115), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT54), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n731_), .A2(new_n732_), .A3(new_n565_), .A4(new_n727_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n730_), .A2(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n314_), .B1(new_n309_), .B2(new_n304_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n303_), .A2(new_n308_), .A3(new_n310_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT118), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n735_), .A2(KEYINPUT118), .A3(new_n736_), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n739_), .A2(new_n316_), .A3(new_n740_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n741_), .A2(new_n284_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT116), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n270_), .A2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT55), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT55), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n270_), .A2(new_n743_), .A3(new_n746_), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n228_), .A2(KEYINPUT68), .A3(new_n246_), .ZN(new_n748_));
  AOI21_X1  g547(.A(KEYINPUT68), .B1(new_n228_), .B2(new_n246_), .ZN(new_n749_));
  NOR3_X1   g548(.A1(new_n748_), .A2(new_n749_), .A3(new_n266_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n254_), .B1(new_n228_), .B2(new_n246_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(KEYINPUT12), .B2(new_n255_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n272_), .B1(new_n750_), .B2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(KEYINPUT117), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT117), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n755_), .B(new_n272_), .C1(new_n750_), .C2(new_n752_), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n745_), .A2(new_n747_), .A3(new_n754_), .A4(new_n756_), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n757_), .A2(KEYINPUT56), .A3(new_n280_), .ZN(new_n758_));
  AOI21_X1  g557(.A(KEYINPUT56), .B1(new_n757_), .B2(new_n280_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n742_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT58), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n565_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n757_), .A2(new_n280_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT56), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n757_), .A2(KEYINPUT56), .A3(new_n280_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n767_), .A2(KEYINPUT119), .A3(KEYINPUT58), .A4(new_n742_), .ZN(new_n768_));
  OAI211_X1 g567(.A(KEYINPUT58), .B(new_n742_), .C1(new_n758_), .C2(new_n759_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT119), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n762_), .A2(new_n768_), .A3(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n284_), .A2(new_n317_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n773_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n286_), .A2(new_n741_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n355_), .B1(new_n774_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT57), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n773_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n780_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(new_n775_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n782_), .A2(KEYINPUT57), .A3(new_n355_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n772_), .A2(new_n779_), .A3(new_n783_), .ZN(new_n784_));
  AND3_X1   g583(.A1(new_n784_), .A2(KEYINPUT120), .A3(new_n331_), .ZN(new_n785_));
  AOI21_X1  g584(.A(KEYINPUT120), .B1(new_n784_), .B2(new_n331_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n734_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n540_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n532_), .A2(new_n399_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n790_), .A2(KEYINPUT59), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n787_), .A2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n790_), .ZN(new_n793_));
  AOI21_X1  g592(.A(KEYINPUT57), .B1(new_n782_), .B2(new_n355_), .ZN(new_n794_));
  AOI211_X1 g593(.A(new_n778_), .B(new_n356_), .C1(new_n781_), .C2(new_n775_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n332_), .B1(new_n796_), .B2(new_n772_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n734_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n793_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT59), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n792_), .A2(new_n317_), .A3(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(G113gat), .ZN(new_n802_));
  OR2_X1    g601(.A1(new_n318_), .A2(G113gat), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n802_), .B1(new_n799_), .B2(new_n803_), .ZN(G1340gat));
  XOR2_X1   g603(.A(KEYINPUT121), .B(G120gat), .Z(new_n805_));
  AOI21_X1  g604(.A(new_n677_), .B1(new_n799_), .B2(KEYINPUT59), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n805_), .B1(new_n792_), .B2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n784_), .A2(new_n331_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n790_), .B1(new_n808_), .B2(new_n734_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n677_), .A2(KEYINPUT60), .ZN(new_n810_));
  MUX2_X1   g609(.A(KEYINPUT60), .B(new_n810_), .S(new_n805_), .Z(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(KEYINPUT122), .B1(new_n807_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n805_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n791_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT120), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n808_), .A2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n784_), .A2(KEYINPUT120), .A3(new_n331_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n816_), .B1(new_n820_), .B2(new_n734_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT59), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n290_), .B1(new_n809_), .B2(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n815_), .B1(new_n821_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT122), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n824_), .A2(new_n825_), .A3(new_n812_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n814_), .A2(new_n826_), .ZN(G1341gat));
  AOI21_X1  g626(.A(G127gat), .B1(new_n809_), .B2(new_n332_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT123), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n828_), .B(new_n829_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n792_), .A2(new_n800_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n332_), .A2(G127gat), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n830_), .B1(new_n831_), .B2(new_n832_), .ZN(G1342gat));
  NAND3_X1  g632(.A1(new_n792_), .A2(new_n566_), .A3(new_n800_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(G134gat), .ZN(new_n835_));
  OR2_X1    g634(.A1(new_n355_), .A2(G134gat), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n835_), .B1(new_n799_), .B2(new_n836_), .ZN(G1343gat));
  NOR2_X1   g636(.A1(new_n797_), .A2(new_n798_), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n619_), .A2(new_n520_), .A3(new_n453_), .A4(new_n399_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n317_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g641(.A1(new_n840_), .A2(new_n290_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n843_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g643(.A(KEYINPUT124), .B(KEYINPUT125), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  XOR2_X1   g645(.A(KEYINPUT61), .B(G155gat), .Z(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n840_), .A2(new_n332_), .A3(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n848_), .B1(new_n840_), .B2(new_n332_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n846_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n851_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n853_), .A2(new_n845_), .A3(new_n849_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n852_), .A2(new_n854_), .ZN(G1346gat));
  AOI21_X1  g654(.A(G162gat), .B1(new_n840_), .B2(new_n356_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n566_), .A2(G162gat), .ZN(new_n857_));
  XOR2_X1   g656(.A(new_n857_), .B(KEYINPUT126), .Z(new_n858_));
  AOI21_X1  g657(.A(new_n856_), .B1(new_n840_), .B2(new_n858_), .ZN(G1347gat));
  INV_X1    g658(.A(KEYINPUT22), .ZN(new_n860_));
  NOR3_X1   g659(.A1(new_n619_), .A2(new_n453_), .A3(new_n541_), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n787_), .A2(new_n860_), .A3(new_n317_), .A4(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(G169gat), .ZN(new_n863_));
  AND3_X1   g662(.A1(new_n862_), .A2(KEYINPUT62), .A3(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n862_), .A2(KEYINPUT62), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT62), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n787_), .A2(new_n866_), .A3(new_n317_), .A4(new_n861_), .ZN(new_n867_));
  AND2_X1   g666(.A1(new_n867_), .A2(G169gat), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n864_), .B1(new_n865_), .B2(new_n868_), .ZN(G1348gat));
  INV_X1    g668(.A(new_n861_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n870_), .B1(new_n820_), .B2(new_n734_), .ZN(new_n871_));
  AOI21_X1  g670(.A(G176gat), .B1(new_n871_), .B2(new_n290_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n838_), .A2(new_n870_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n873_), .A2(G176gat), .A3(new_n290_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(KEYINPUT127), .B1(new_n872_), .B2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT127), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n787_), .A2(new_n861_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n878_), .A2(new_n677_), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n877_), .B(new_n874_), .C1(new_n879_), .C2(G176gat), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n876_), .A2(new_n880_), .ZN(G1349gat));
  AOI21_X1  g680(.A(G183gat), .B1(new_n873_), .B2(new_n332_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n331_), .A2(new_n368_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n882_), .B1(new_n871_), .B2(new_n883_), .ZN(G1350gat));
  OAI21_X1  g683(.A(G190gat), .B1(new_n878_), .B2(new_n565_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n871_), .A2(new_n356_), .A3(new_n459_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(G1351gat));
  NAND3_X1  g686(.A1(new_n453_), .A2(new_n532_), .A3(new_n399_), .ZN(new_n888_));
  NOR3_X1   g687(.A1(new_n838_), .A2(new_n619_), .A3(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(new_n317_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n290_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g692(.A1(new_n889_), .A2(new_n332_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(KEYINPUT63), .B(G211gat), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n896_), .B1(new_n894_), .B2(new_n897_), .ZN(G1354gat));
  INV_X1    g697(.A(G218gat), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n889_), .A2(new_n899_), .A3(new_n356_), .ZN(new_n900_));
  AND2_X1   g699(.A1(new_n889_), .A2(new_n566_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(new_n899_), .ZN(G1355gat));
endmodule


