//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 0 1 0 0 0 1 1 0 1 1 1 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 0 1 0 1 0 0 1 1 0 0 1 0 0 1 1 1 0 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n665_,
    new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n750_, new_n751_, new_n752_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n776_, new_n777_, new_n778_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n864_, new_n865_, new_n866_, new_n867_, new_n869_,
    new_n870_, new_n871_, new_n873_, new_n874_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n910_, new_n912_,
    new_n913_, new_n914_, new_n915_, new_n917_, new_n918_, new_n919_,
    new_n921_, new_n923_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_, new_n930_;
  NAND2_X1  g000(.A1(G99gat), .A2(G106gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT6), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT6), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n204_), .A2(G99gat), .A3(G106gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT7), .ZN(new_n208_));
  INV_X1    g007(.A(G99gat), .ZN(new_n209_));
  INV_X1    g008(.A(G106gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n208_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n206_), .A2(new_n207_), .A3(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT66), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(G85gat), .ZN(new_n215_));
  INV_X1    g014(.A(G92gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G85gat), .A2(G92gat), .ZN(new_n218_));
  AND2_X1   g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n206_), .A2(KEYINPUT66), .A3(new_n207_), .A4(new_n211_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT67), .B(KEYINPUT8), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n214_), .A2(new_n219_), .A3(new_n220_), .A4(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT68), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT8), .ZN(new_n224_));
  AOI211_X1 g023(.A(new_n223_), .B(new_n224_), .C1(new_n212_), .C2(new_n219_), .ZN(new_n225_));
  AND2_X1   g024(.A1(new_n203_), .A2(new_n205_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n211_), .A2(new_n207_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n219_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(KEYINPUT68), .B1(new_n228_), .B2(KEYINPUT8), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n222_), .B1(new_n225_), .B2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G29gat), .B(G36gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G43gat), .B(G50gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n231_), .B(new_n232_), .ZN(new_n233_));
  AND2_X1   g032(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n234_));
  NOR2_X1   g033(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n235_));
  NOR3_X1   g034(.A1(new_n234_), .A2(new_n235_), .A3(KEYINPUT64), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT64), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT10), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(new_n209_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n237_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n210_), .B1(new_n236_), .B2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n217_), .A2(KEYINPUT9), .A3(new_n218_), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n218_), .A2(KEYINPUT9), .ZN(new_n244_));
  AND3_X1   g043(.A1(new_n206_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(KEYINPUT65), .B1(new_n242_), .B2(new_n245_), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT64), .B1(new_n234_), .B2(new_n235_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n239_), .A2(new_n237_), .A3(new_n240_), .ZN(new_n248_));
  AOI21_X1  g047(.A(G106gat), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n206_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT65), .ZN(new_n251_));
  NOR3_X1   g050(.A1(new_n249_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n246_), .A2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n230_), .A2(new_n233_), .A3(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n242_), .A2(new_n245_), .A3(KEYINPUT65), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n251_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n255_), .A2(KEYINPUT69), .A3(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(KEYINPUT69), .B1(new_n255_), .B2(new_n256_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n230_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT70), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n230_), .B(KEYINPUT70), .C1(new_n257_), .C2(new_n258_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n233_), .B(KEYINPUT15), .ZN(new_n264_));
  AOI21_X1  g063(.A(KEYINPUT73), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT73), .ZN(new_n266_));
  INV_X1    g065(.A(new_n264_), .ZN(new_n267_));
  AOI211_X1 g066(.A(new_n266_), .B(new_n267_), .C1(new_n261_), .C2(new_n262_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n254_), .B1(new_n265_), .B2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G232gat), .A2(G233gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT34), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT35), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n269_), .A2(new_n273_), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n271_), .A2(KEYINPUT35), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n275_), .B1(new_n272_), .B2(KEYINPUT74), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n276_), .B1(KEYINPUT74), .B2(new_n272_), .ZN(new_n277_));
  AND2_X1   g076(.A1(new_n254_), .A2(new_n277_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n278_), .B1(new_n265_), .B2(new_n268_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n274_), .A2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G190gat), .B(G218gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G134gat), .B(G162gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  XOR2_X1   g082(.A(new_n283_), .B(KEYINPUT36), .Z(new_n284_));
  NAND2_X1  g083(.A1(new_n280_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n262_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT69), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n287_), .B1(new_n246_), .B2(new_n252_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n255_), .A2(new_n256_), .A3(KEYINPUT69), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(KEYINPUT70), .B1(new_n290_), .B2(new_n230_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n264_), .B1(new_n286_), .B2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(new_n266_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n263_), .A2(KEYINPUT73), .A3(new_n264_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n272_), .B1(new_n295_), .B2(new_n254_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n283_), .A2(KEYINPUT36), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n279_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT75), .ZN(new_n299_));
  NOR3_X1   g098(.A1(new_n296_), .A2(new_n298_), .A3(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n297_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n301_), .B1(new_n295_), .B2(new_n278_), .ZN(new_n302_));
  AOI21_X1  g101(.A(KEYINPUT75), .B1(new_n302_), .B2(new_n274_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n285_), .B1(new_n300_), .B2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT37), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n299_), .B1(new_n296_), .B2(new_n298_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n302_), .A2(new_n274_), .A3(KEYINPUT75), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n309_), .A2(KEYINPUT37), .A3(new_n285_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n306_), .A2(new_n310_), .ZN(new_n311_));
  XOR2_X1   g110(.A(G127gat), .B(G155gat), .Z(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT16), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G183gat), .B(G211gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT78), .B(KEYINPUT17), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G231gat), .A2(G233gat), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n317_), .B(KEYINPUT77), .Z(new_n318_));
  XOR2_X1   g117(.A(new_n318_), .B(KEYINPUT76), .Z(new_n319_));
  XNOR2_X1  g118(.A(G15gat), .B(G22gat), .ZN(new_n320_));
  INV_X1    g119(.A(G1gat), .ZN(new_n321_));
  INV_X1    g120(.A(G8gat), .ZN(new_n322_));
  OAI21_X1  g121(.A(KEYINPUT14), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n320_), .A2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G1gat), .B(G8gat), .ZN(new_n325_));
  XOR2_X1   g124(.A(new_n324_), .B(new_n325_), .Z(new_n326_));
  XNOR2_X1  g125(.A(new_n319_), .B(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G57gat), .B(G64gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT11), .ZN(new_n329_));
  XOR2_X1   g128(.A(G71gat), .B(G78gat), .Z(new_n330_));
  AND2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n331_), .B1(KEYINPUT11), .B2(new_n328_), .ZN(new_n332_));
  OR2_X1    g131(.A1(new_n329_), .A2(new_n330_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n327_), .B(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  AOI211_X1 g136(.A(new_n315_), .B(new_n316_), .C1(new_n337_), .C2(KEYINPUT71), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n338_), .B1(KEYINPUT71), .B2(new_n337_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n315_), .B(KEYINPUT17), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n336_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n311_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT71), .ZN(new_n344_));
  OAI21_X1  g143(.A(KEYINPUT12), .B1(new_n334_), .B2(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n345_), .B1(new_n344_), .B2(new_n334_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n263_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G230gat), .A2(G233gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n230_), .A2(new_n253_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n349_), .A2(new_n335_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT12), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n349_), .A2(new_n335_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n350_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n347_), .A2(new_n348_), .A3(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n348_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n352_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n355_), .B1(new_n356_), .B2(new_n350_), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n354_), .A2(new_n357_), .ZN(new_n358_));
  XOR2_X1   g157(.A(G120gat), .B(G148gat), .Z(new_n359_));
  XNOR2_X1  g158(.A(G176gat), .B(G204gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n362_));
  XOR2_X1   g161(.A(new_n361_), .B(new_n362_), .Z(new_n363_));
  OR2_X1    g162(.A1(new_n358_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n358_), .A2(new_n363_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT13), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n343_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(G169gat), .ZN(new_n370_));
  INV_X1    g169(.A(G176gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G169gat), .A2(G176gat), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n372_), .A2(KEYINPUT24), .A3(new_n373_), .ZN(new_n374_));
  XOR2_X1   g173(.A(new_n374_), .B(KEYINPUT85), .Z(new_n375_));
  INV_X1    g174(.A(KEYINPUT23), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n376_), .A2(G183gat), .A3(G190gat), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G183gat), .A2(G190gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT23), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT86), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT86), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n379_), .A2(new_n382_), .A3(KEYINPUT23), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n378_), .B1(new_n381_), .B2(new_n383_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n372_), .A2(KEYINPUT24), .ZN(new_n385_));
  OAI21_X1  g184(.A(KEYINPUT87), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n383_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n382_), .B1(new_n379_), .B2(KEYINPUT23), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n377_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT87), .ZN(new_n390_));
  INV_X1    g189(.A(new_n385_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n389_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT25), .B(G183gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT26), .B(G190gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(KEYINPUT84), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT84), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n393_), .A2(new_n394_), .A3(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n396_), .A2(new_n398_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n375_), .A2(new_n386_), .A3(new_n392_), .A4(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(G169gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n380_), .A2(new_n377_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(G183gat), .A2(G190gat), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n402_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n400_), .A2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(KEYINPUT30), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G227gat), .A2(G233gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(G15gat), .ZN(new_n410_));
  INV_X1    g209(.A(G43gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n410_), .B(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G71gat), .B(G99gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n412_), .B(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n408_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT88), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n415_), .B(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n408_), .A2(new_n414_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT89), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G127gat), .B(G134gat), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT90), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G113gat), .B(G120gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT31), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n417_), .A2(new_n420_), .A3(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n426_), .B1(new_n417_), .B2(new_n420_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G78gat), .B(G106gat), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G228gat), .A2(G233gat), .ZN(new_n433_));
  OR2_X1    g232(.A1(G197gat), .A2(G204gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G197gat), .A2(G204gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT21), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT95), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n434_), .A2(KEYINPUT21), .A3(new_n435_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G211gat), .B(G218gat), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n438_), .A2(new_n439_), .A3(new_n440_), .A4(new_n441_), .ZN(new_n442_));
  AND3_X1   g241(.A1(new_n438_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT95), .B1(new_n440_), .B2(new_n441_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n442_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G155gat), .A2(G162gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(KEYINPUT91), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT91), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n448_), .A2(G155gat), .A3(G162gat), .ZN(new_n449_));
  INV_X1    g248(.A(G155gat), .ZN(new_n450_));
  INV_X1    g249(.A(G162gat), .ZN(new_n451_));
  AOI22_X1  g250(.A1(new_n447_), .A2(new_n449_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G141gat), .A2(G148gat), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT93), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT2), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n453_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT3), .ZN(new_n457_));
  INV_X1    g256(.A(G141gat), .ZN(new_n458_));
  INV_X1    g257(.A(G148gat), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n457_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n456_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n455_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n452_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT94), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT94), .ZN(new_n466_));
  OAI211_X1 g265(.A(new_n452_), .B(new_n466_), .C1(new_n462_), .C2(new_n463_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n465_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n447_), .A2(new_n449_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT1), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT1), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n447_), .A2(new_n449_), .A3(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n450_), .A2(new_n451_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n470_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT92), .ZN(new_n475_));
  XOR2_X1   g274(.A(G141gat), .B(G148gat), .Z(new_n476_));
  AND3_X1   g275(.A1(new_n474_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n475_), .B1(new_n474_), .B2(new_n476_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n468_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT29), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT97), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n445_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n479_), .A2(KEYINPUT97), .A3(KEYINPUT29), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n433_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT96), .ZN(new_n485_));
  OAI211_X1 g284(.A(new_n442_), .B(new_n433_), .C1(new_n443_), .C2(new_n444_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n485_), .B1(new_n480_), .B2(new_n487_), .ZN(new_n488_));
  AOI211_X1 g287(.A(KEYINPUT96), .B(new_n486_), .C1(new_n479_), .C2(KEYINPUT29), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  OAI211_X1 g289(.A(KEYINPUT98), .B(new_n432_), .C1(new_n484_), .C2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G22gat), .B(G50gat), .ZN(new_n492_));
  OR3_X1    g291(.A1(new_n479_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT28), .B1(new_n479_), .B2(KEYINPUT29), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n492_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n493_), .A2(new_n494_), .A3(new_n492_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n484_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n490_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  XOR2_X1   g300(.A(new_n431_), .B(KEYINPUT98), .Z(new_n502_));
  OAI211_X1 g301(.A(new_n491_), .B(new_n498_), .C1(new_n501_), .C2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n431_), .A2(KEYINPUT99), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n499_), .A2(new_n500_), .A3(new_n504_), .ZN(new_n505_));
  OAI211_X1 g304(.A(KEYINPUT99), .B(new_n431_), .C1(new_n484_), .C2(new_n490_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n497_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n507_), .A2(new_n495_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n505_), .A2(new_n506_), .A3(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n503_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G8gat), .B(G36gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT18), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G64gat), .B(G92gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT32), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G226gat), .A2(G233gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT19), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT20), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT100), .ZN(new_n521_));
  AND3_X1   g320(.A1(new_n395_), .A2(new_n521_), .A3(new_n374_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n521_), .B1(new_n395_), .B2(new_n374_), .ZN(new_n523_));
  OAI211_X1 g322(.A(new_n391_), .B(new_n403_), .C1(new_n522_), .C2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(KEYINPUT22), .B(G169gat), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT101), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  AND2_X1   g326(.A1(new_n370_), .A2(KEYINPUT22), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n370_), .A2(KEYINPUT22), .ZN(new_n529_));
  NOR3_X1   g328(.A1(new_n528_), .A2(new_n529_), .A3(KEYINPUT101), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n371_), .B1(new_n527_), .B2(new_n530_), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n531_), .B(new_n373_), .C1(new_n384_), .C2(new_n405_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n524_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n445_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n520_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n400_), .A2(new_n406_), .A3(new_n445_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n519_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n524_), .A2(new_n532_), .A3(new_n445_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT20), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n445_), .B1(new_n400_), .B2(new_n406_), .ZN(new_n540_));
  NOR3_X1   g339(.A1(new_n539_), .A2(new_n540_), .A3(new_n518_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n516_), .B1(new_n537_), .B2(new_n541_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n518_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n535_), .A2(new_n519_), .A3(new_n536_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n542_), .B1(new_n516_), .B2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G1gat), .B(G29gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(G85gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(KEYINPUT0), .B(G57gat), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n548_), .B(new_n549_), .Z(new_n550_));
  NAND2_X1  g349(.A1(G225gat), .A2(G233gat), .ZN(new_n551_));
  XOR2_X1   g350(.A(new_n423_), .B(new_n424_), .Z(new_n552_));
  NAND3_X1  g351(.A1(new_n479_), .A2(new_n552_), .A3(KEYINPUT102), .ZN(new_n553_));
  OAI211_X1 g352(.A(new_n425_), .B(new_n468_), .C1(new_n478_), .C2(new_n477_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n553_), .A2(KEYINPUT4), .A3(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT4), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n479_), .A2(new_n552_), .A3(KEYINPUT102), .A4(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n551_), .B1(new_n555_), .B2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n551_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n479_), .A2(new_n552_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n559_), .B1(new_n560_), .B2(new_n554_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n550_), .B1(new_n558_), .B2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT105), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n555_), .A2(new_n557_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(new_n559_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n561_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n550_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n566_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT106), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT106), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n566_), .A2(new_n567_), .A3(new_n571_), .A4(new_n568_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n546_), .B1(new_n564_), .B2(new_n573_), .ZN(new_n574_));
  NOR3_X1   g373(.A1(new_n537_), .A2(new_n541_), .A3(new_n514_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n533_), .A2(new_n534_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n576_), .A2(new_n536_), .A3(KEYINPUT20), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(new_n518_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n540_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n579_), .A2(KEYINPUT20), .A3(new_n519_), .A4(new_n538_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n515_), .B1(new_n578_), .B2(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n575_), .A2(new_n581_), .ZN(new_n582_));
  OAI211_X1 g381(.A(KEYINPUT33), .B(new_n550_), .C1(new_n558_), .C2(new_n561_), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT33), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n562_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT103), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n560_), .A2(new_n554_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n550_), .B1(new_n589_), .B2(new_n559_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n590_), .B1(new_n559_), .B2(new_n565_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT104), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n590_), .B(KEYINPUT104), .C1(new_n559_), .C2(new_n565_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n562_), .A2(KEYINPUT103), .A3(new_n585_), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n584_), .A2(new_n588_), .A3(new_n595_), .A4(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n510_), .B1(new_n574_), .B2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n562_), .B(KEYINPUT105), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT27), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n600_), .B1(new_n575_), .B2(new_n581_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n545_), .A2(new_n514_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n578_), .A2(new_n580_), .A3(new_n515_), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n602_), .A2(new_n603_), .A3(KEYINPUT107), .A4(KEYINPUT27), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n601_), .A2(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n537_), .A2(new_n541_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n600_), .B1(new_n606_), .B2(new_n515_), .ZN(new_n607_));
  AOI21_X1  g406(.A(KEYINPUT107), .B1(new_n607_), .B2(new_n602_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n605_), .A2(new_n608_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n570_), .A2(new_n572_), .ZN(new_n610_));
  AND4_X1   g409(.A1(new_n599_), .A2(new_n609_), .A3(new_n510_), .A4(new_n610_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n430_), .B1(new_n598_), .B2(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n564_), .A2(new_n573_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n429_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n510_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(new_n609_), .ZN(new_n616_));
  OR2_X1    g415(.A1(new_n614_), .A2(new_n616_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n612_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n326_), .A2(new_n233_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT79), .ZN(new_n620_));
  OR2_X1    g419(.A1(new_n326_), .A2(new_n233_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(KEYINPUT80), .ZN(new_n623_));
  NAND2_X1  g422(.A1(G229gat), .A2(G233gat), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT80), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n620_), .A2(new_n626_), .A3(new_n621_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n623_), .A2(new_n625_), .A3(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n620_), .B1(new_n326_), .B2(new_n267_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(new_n624_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(G113gat), .B(G141gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(G169gat), .B(G197gat), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(KEYINPUT81), .B(KEYINPUT82), .ZN(new_n634_));
  XOR2_X1   g433(.A(new_n633_), .B(new_n634_), .Z(new_n635_));
  NAND3_X1  g434(.A1(new_n628_), .A2(new_n630_), .A3(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n628_), .A2(new_n630_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n635_), .ZN(new_n638_));
  AOI21_X1  g437(.A(KEYINPUT83), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT83), .ZN(new_n640_));
  AOI211_X1 g439(.A(new_n640_), .B(new_n635_), .C1(new_n628_), .C2(new_n630_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n636_), .B1(new_n639_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n618_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n369_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n613_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n646_), .A2(new_n321_), .A3(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT38), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n304_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n618_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n367_), .ZN(new_n653_));
  NOR3_X1   g452(.A1(new_n653_), .A2(new_n643_), .A3(new_n342_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n652_), .A2(new_n654_), .ZN(new_n655_));
  OAI21_X1  g454(.A(G1gat), .B1(new_n655_), .B2(new_n613_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n648_), .A2(new_n649_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n650_), .A2(new_n656_), .A3(new_n657_), .ZN(G1324gat));
  OAI21_X1  g457(.A(G8gat), .B1(new_n655_), .B2(new_n609_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT39), .ZN(new_n660_));
  INV_X1    g459(.A(new_n609_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n646_), .A2(new_n322_), .A3(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n662_), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g463(.A(G15gat), .B1(new_n655_), .B2(new_n430_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT41), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n645_), .A2(G15gat), .A3(new_n430_), .ZN(new_n667_));
  OR2_X1    g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1326gat));
  OAI21_X1  g467(.A(G22gat), .B1(new_n655_), .B2(new_n615_), .ZN(new_n669_));
  XOR2_X1   g468(.A(KEYINPUT108), .B(KEYINPUT42), .Z(new_n670_));
  XNOR2_X1  g469(.A(new_n669_), .B(new_n670_), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n615_), .A2(G22gat), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n671_), .B1(new_n645_), .B2(new_n672_), .ZN(G1327gat));
  NAND2_X1  g472(.A1(new_n612_), .A2(new_n617_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT43), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n674_), .A2(new_n675_), .A3(new_n311_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT109), .ZN(new_n677_));
  AOI221_X4 g476(.A(new_n305_), .B1(new_n280_), .B2(new_n284_), .C1(new_n307_), .C2(new_n308_), .ZN(new_n678_));
  AOI21_X1  g477(.A(KEYINPUT37), .B1(new_n309_), .B2(new_n285_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n677_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n306_), .A2(KEYINPUT109), .A3(new_n310_), .ZN(new_n681_));
  AOI22_X1  g480(.A1(new_n680_), .A2(new_n681_), .B1(new_n612_), .B2(new_n617_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n676_), .B1(new_n682_), .B2(new_n675_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n342_), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n653_), .A2(new_n643_), .A3(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n683_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT110), .ZN(new_n687_));
  AOI21_X1  g486(.A(KEYINPUT44), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n683_), .A2(KEYINPUT110), .A3(new_n685_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n686_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(KEYINPUT44), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n690_), .A2(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(G29gat), .B1(new_n693_), .B2(new_n613_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT111), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n304_), .A2(new_n684_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n367_), .A2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n644_), .A2(new_n697_), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n698_), .A2(G29gat), .A3(new_n613_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n694_), .A2(new_n695_), .A3(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(G29gat), .ZN(new_n702_));
  AOI22_X1  g501(.A1(new_n688_), .A2(new_n689_), .B1(KEYINPUT44), .B2(new_n691_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n702_), .B1(new_n703_), .B2(new_n647_), .ZN(new_n704_));
  OAI21_X1  g503(.A(KEYINPUT111), .B1(new_n704_), .B2(new_n699_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n701_), .A2(new_n705_), .ZN(G1328gat));
  OAI21_X1  g505(.A(G36gat), .B1(new_n693_), .B2(new_n609_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(KEYINPUT113), .A2(KEYINPUT46), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n698_), .ZN(new_n710_));
  INV_X1    g509(.A(G36gat), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n710_), .A2(new_n711_), .A3(new_n661_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(KEYINPUT112), .B(KEYINPUT45), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n712_), .B(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n707_), .A2(new_n709_), .A3(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n711_), .B1(new_n703_), .B2(new_n661_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n708_), .B1(new_n717_), .B2(new_n714_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(G1329gat));
  OAI21_X1  g518(.A(new_n411_), .B1(new_n698_), .B2(new_n430_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n429_), .A2(G43gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n720_), .B1(new_n693_), .B2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(KEYINPUT47), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT47), .ZN(new_n724_));
  OAI211_X1 g523(.A(new_n724_), .B(new_n720_), .C1(new_n693_), .C2(new_n721_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(G1330gat));
  AOI21_X1  g525(.A(G50gat), .B1(new_n710_), .B2(new_n510_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n510_), .A2(G50gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n727_), .B1(new_n703_), .B2(new_n728_), .ZN(G1331gat));
  NAND3_X1  g528(.A1(new_n674_), .A2(new_n643_), .A3(new_n653_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(new_n343_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(G57gat), .B1(new_n733_), .B2(new_n647_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n367_), .A2(new_n642_), .A3(new_n342_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n652_), .A2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(G57gat), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n738_), .B1(new_n647_), .B2(KEYINPUT114), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n739_), .B1(KEYINPUT114), .B2(new_n738_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n734_), .B1(new_n737_), .B2(new_n740_), .ZN(G1332gat));
  OAI21_X1  g540(.A(G64gat), .B1(new_n736_), .B2(new_n609_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT48), .ZN(new_n743_));
  OR2_X1    g542(.A1(new_n609_), .A2(G64gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n743_), .B1(new_n732_), .B2(new_n744_), .ZN(G1333gat));
  OAI21_X1  g544(.A(G71gat), .B1(new_n736_), .B2(new_n430_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT49), .ZN(new_n747_));
  OR2_X1    g546(.A1(new_n430_), .A2(G71gat), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n747_), .B1(new_n732_), .B2(new_n748_), .ZN(G1334gat));
  OAI21_X1  g548(.A(G78gat), .B1(new_n736_), .B2(new_n615_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT50), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n615_), .A2(G78gat), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n751_), .B1(new_n732_), .B2(new_n752_), .ZN(G1335gat));
  NAND2_X1  g552(.A1(new_n731_), .A2(new_n696_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n755_), .A2(new_n215_), .A3(new_n647_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT116), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT115), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n367_), .A2(new_n642_), .A3(new_n684_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n683_), .A2(new_n758_), .A3(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n758_), .B1(new_n683_), .B2(new_n759_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n757_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n683_), .A2(new_n759_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(KEYINPUT115), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n765_), .A2(KEYINPUT116), .A3(new_n760_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n613_), .B1(new_n763_), .B2(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n756_), .B1(new_n767_), .B2(new_n215_), .ZN(G1336gat));
  NAND3_X1  g567(.A1(new_n755_), .A2(new_n216_), .A3(new_n661_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n609_), .B1(new_n763_), .B2(new_n766_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n769_), .B1(new_n770_), .B2(new_n216_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT117), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT117), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n773_), .B(new_n769_), .C1(new_n770_), .C2(new_n216_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(G1337gat));
  OAI211_X1 g574(.A(new_n755_), .B(new_n429_), .C1(new_n236_), .C2(new_n241_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n430_), .B1(new_n765_), .B2(new_n760_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n776_), .B1(new_n777_), .B2(new_n209_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND2_X1  g578(.A1(new_n680_), .A2(new_n681_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n675_), .B1(new_n780_), .B2(new_n674_), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n674_), .A2(new_n675_), .A3(new_n311_), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n510_), .B(new_n759_), .C1(new_n781_), .C2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT118), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n683_), .A2(KEYINPUT118), .A3(new_n510_), .A4(new_n759_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(G106gat), .ZN(new_n787_));
  OAI21_X1  g586(.A(KEYINPUT119), .B1(new_n785_), .B2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n783_), .A2(new_n784_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT119), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n789_), .A2(new_n790_), .A3(G106gat), .A4(new_n786_), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n788_), .A2(KEYINPUT52), .A3(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n793_));
  OAI211_X1 g592(.A(KEYINPUT119), .B(new_n793_), .C1(new_n785_), .C2(new_n787_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n755_), .A2(new_n210_), .A3(new_n510_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(KEYINPUT53), .B1(new_n792_), .B2(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n788_), .A2(KEYINPUT52), .A3(new_n791_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT53), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n798_), .A2(new_n799_), .A3(new_n794_), .A4(new_n795_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n797_), .A2(new_n800_), .ZN(G1339gat));
  INV_X1    g600(.A(KEYINPUT56), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT121), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n354_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(KEYINPUT120), .ZN(new_n807_));
  OR2_X1    g606(.A1(new_n354_), .A2(new_n805_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT120), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n354_), .A2(new_n809_), .A3(new_n805_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n347_), .A2(new_n353_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n355_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n807_), .A2(new_n808_), .A3(new_n810_), .A4(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n363_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n804_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n642_), .A2(new_n365_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n813_), .A2(new_n814_), .A3(new_n804_), .ZN(new_n818_));
  AND2_X1   g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n625_), .B1(new_n623_), .B2(new_n627_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n635_), .B1(new_n629_), .B2(new_n624_), .ZN(new_n821_));
  OAI22_X1  g620(.A1(new_n639_), .A2(new_n641_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n822_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n823_));
  OAI211_X1 g622(.A(KEYINPUT57), .B(new_n304_), .C1(new_n819_), .C2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT57), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n823_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n825_), .B1(new_n826_), .B2(new_n651_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(KEYINPUT122), .A2(KEYINPUT56), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n813_), .A2(new_n814_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(KEYINPUT122), .A2(KEYINPUT56), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n829_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n832_), .B1(new_n831_), .B2(new_n830_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n822_), .B1(new_n358_), .B2(new_n363_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n833_), .A2(KEYINPUT58), .A3(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n311_), .ZN(new_n836_));
  AOI21_X1  g635(.A(KEYINPUT58), .B1(new_n833_), .B2(new_n834_), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n824_), .B(new_n827_), .C1(new_n836_), .C2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n342_), .ZN(new_n839_));
  OAI21_X1  g638(.A(KEYINPUT54), .B1(new_n368_), .B2(new_n642_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT54), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n343_), .A2(new_n841_), .A3(new_n643_), .A4(new_n367_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n840_), .A2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n839_), .A2(new_n843_), .ZN(new_n844_));
  NOR3_X1   g643(.A1(new_n430_), .A2(new_n616_), .A3(new_n613_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(G113gat), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n847_), .A2(new_n848_), .A3(new_n642_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n847_), .A2(KEYINPUT59), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT59), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n846_), .A2(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n643_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n849_), .B1(new_n853_), .B2(new_n848_), .ZN(G1340gat));
  INV_X1    g653(.A(G120gat), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n855_), .B1(new_n367_), .B2(KEYINPUT60), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n847_), .B(new_n856_), .C1(KEYINPUT60), .C2(new_n855_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n367_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n858_), .B2(new_n855_), .ZN(G1341gat));
  INV_X1    g658(.A(G127gat), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n847_), .A2(new_n860_), .A3(new_n684_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n342_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(new_n862_), .B2(new_n860_), .ZN(G1342gat));
  AOI21_X1  g662(.A(G134gat), .B1(new_n847_), .B2(new_n651_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n850_), .A2(new_n852_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n311_), .A2(G134gat), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(KEYINPUT123), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n864_), .B1(new_n865_), .B2(new_n867_), .ZN(G1343gat));
  NOR4_X1   g667(.A1(new_n661_), .A2(new_n429_), .A3(new_n613_), .A4(new_n615_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n844_), .A2(new_n869_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n870_), .A2(new_n643_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(new_n458_), .ZN(G1344gat));
  NOR2_X1   g671(.A1(new_n870_), .A2(new_n367_), .ZN(new_n873_));
  XOR2_X1   g672(.A(KEYINPUT124), .B(G148gat), .Z(new_n874_));
  XNOR2_X1  g673(.A(new_n873_), .B(new_n874_), .ZN(G1345gat));
  INV_X1    g674(.A(new_n870_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT125), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n876_), .A2(new_n877_), .A3(new_n684_), .ZN(new_n878_));
  OAI21_X1  g677(.A(KEYINPUT125), .B1(new_n870_), .B2(new_n342_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(KEYINPUT61), .B(G155gat), .ZN(new_n880_));
  AND3_X1   g679(.A1(new_n878_), .A2(new_n879_), .A3(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n880_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n881_), .A2(new_n882_), .ZN(G1346gat));
  AOI21_X1  g682(.A(G162gat), .B1(new_n876_), .B2(new_n651_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n451_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n884_), .B1(new_n876_), .B2(new_n885_), .ZN(G1347gat));
  INV_X1    g685(.A(KEYINPUT127), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT126), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n370_), .B1(new_n888_), .B2(KEYINPUT62), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n614_), .A2(new_n510_), .A3(new_n609_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n892_), .B1(new_n839_), .B2(new_n843_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n890_), .B1(new_n893_), .B2(new_n642_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n888_), .A2(KEYINPUT62), .ZN(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n893_), .A2(new_n642_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n527_), .A2(new_n530_), .ZN(new_n898_));
  OAI22_X1  g697(.A1(new_n894_), .A2(new_n896_), .B1(new_n897_), .B2(new_n898_), .ZN(new_n899_));
  AOI211_X1 g698(.A(new_n895_), .B(new_n890_), .C1(new_n893_), .C2(new_n642_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n887_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n897_), .A2(new_n889_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(new_n895_), .ZN(new_n903_));
  OR2_X1    g702(.A1(new_n897_), .A2(new_n898_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n894_), .A2(new_n896_), .ZN(new_n905_));
  NAND4_X1  g704(.A1(new_n903_), .A2(new_n904_), .A3(KEYINPUT127), .A4(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n901_), .A2(new_n906_), .ZN(G1348gat));
  NAND2_X1  g706(.A1(new_n893_), .A2(new_n653_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g708(.A1(new_n893_), .A2(new_n684_), .ZN(new_n910_));
  MUX2_X1   g709(.A(new_n393_), .B(G183gat), .S(new_n910_), .Z(G1350gat));
  INV_X1    g710(.A(new_n893_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n311_), .ZN(new_n913_));
  OAI21_X1  g712(.A(G190gat), .B1(new_n912_), .B2(new_n913_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n893_), .A2(new_n394_), .A3(new_n651_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(G1351gat));
  NAND4_X1  g715(.A1(new_n430_), .A2(new_n613_), .A3(new_n510_), .A4(new_n661_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n917_), .B1(new_n839_), .B2(new_n843_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(new_n642_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g719(.A1(new_n918_), .A2(new_n653_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g721(.A1(new_n918_), .A2(new_n684_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n924_));
  AND2_X1   g723(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n925_));
  NOR3_X1   g724(.A1(new_n923_), .A2(new_n924_), .A3(new_n925_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n926_), .B1(new_n923_), .B2(new_n924_), .ZN(G1354gat));
  INV_X1    g726(.A(G218gat), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n918_), .A2(new_n928_), .A3(new_n651_), .ZN(new_n929_));
  AND2_X1   g728(.A1(new_n918_), .A2(new_n311_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n929_), .B1(new_n930_), .B2(new_n928_), .ZN(G1355gat));
endmodule


