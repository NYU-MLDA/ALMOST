//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 1 1 0 1 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 0 0 1 1 1 0 1 1 1 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n797_, new_n798_, new_n799_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n839_, new_n840_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_,
    new_n859_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_, new_n944_, new_n945_, new_n947_, new_n949_,
    new_n950_, new_n952_, new_n953_, new_n954_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n976_,
    new_n977_, new_n979_, new_n980_, new_n982_, new_n983_, new_n984_,
    new_n985_, new_n986_, new_n987_, new_n988_, new_n989_, new_n990_,
    new_n991_, new_n993_, new_n994_, new_n995_, new_n997_, new_n998_,
    new_n999_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1006_,
    new_n1007_;
  INV_X1    g000(.A(KEYINPUT27), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT98), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G169gat), .A2(G176gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT24), .ZN(new_n205_));
  INV_X1    g004(.A(G169gat), .ZN(new_n206_));
  INV_X1    g005(.A(G176gat), .ZN(new_n207_));
  AOI22_X1  g006(.A1(new_n205_), .A2(KEYINPUT95), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n208_), .B1(KEYINPUT95), .B2(new_n205_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n206_), .A2(new_n207_), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n212_), .B(new_n213_), .C1(new_n214_), .C2(KEYINPUT24), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n209_), .A2(new_n216_), .ZN(new_n217_));
  XOR2_X1   g016(.A(KEYINPUT25), .B(G183gat), .Z(new_n218_));
  XOR2_X1   g017(.A(KEYINPUT26), .B(G190gat), .Z(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT94), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT26), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(G190gat), .ZN(new_n222_));
  OR2_X1    g021(.A1(new_n221_), .A2(G190gat), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT94), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n218_), .B1(new_n220_), .B2(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n217_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n213_), .ZN(new_n228_));
  AOI21_X1  g027(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n229_));
  NOR2_X1   g028(.A1(G183gat), .A2(G190gat), .ZN(new_n230_));
  NOR3_X1   g029(.A1(new_n228_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  OR2_X1    g031(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n234_));
  AOI21_X1  g033(.A(G176gat), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT96), .ZN(new_n236_));
  INV_X1    g035(.A(new_n204_), .ZN(new_n237_));
  NOR3_X1   g036(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n234_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n207_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(KEYINPUT96), .B1(new_n241_), .B2(new_n204_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n232_), .B1(new_n238_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT97), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n236_), .B1(new_n235_), .B2(new_n237_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n241_), .A2(KEYINPUT96), .A3(new_n204_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n248_), .A2(KEYINPUT97), .A3(new_n232_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n227_), .B1(new_n245_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT21), .ZN(new_n251_));
  INV_X1    g050(.A(G197gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(G204gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT90), .B(G204gat), .ZN(new_n254_));
  OAI211_X1 g053(.A(new_n251_), .B(new_n253_), .C1(new_n254_), .C2(new_n252_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT91), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(G204gat), .ZN(new_n258_));
  AND2_X1   g057(.A1(new_n258_), .A2(KEYINPUT90), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n258_), .A2(KEYINPUT90), .ZN(new_n260_));
  OAI21_X1  g059(.A(G197gat), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n261_), .A2(KEYINPUT91), .A3(new_n251_), .A4(new_n253_), .ZN(new_n262_));
  XOR2_X1   g061(.A(G211gat), .B(G218gat), .Z(new_n263_));
  OAI21_X1  g062(.A(new_n252_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n251_), .B1(G197gat), .B2(G204gat), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n263_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n257_), .A2(new_n262_), .A3(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n261_), .A2(new_n253_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n268_), .A2(KEYINPUT21), .A3(new_n263_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n203_), .B1(new_n250_), .B2(new_n271_), .ZN(new_n272_));
  AND2_X1   g071(.A1(new_n220_), .A2(new_n225_), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n216_), .B(new_n209_), .C1(new_n273_), .C2(new_n218_), .ZN(new_n274_));
  AOI21_X1  g073(.A(KEYINPUT97), .B1(new_n248_), .B2(new_n232_), .ZN(new_n275_));
  AOI211_X1 g074(.A(new_n244_), .B(new_n231_), .C1(new_n246_), .C2(new_n247_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n274_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n277_), .A2(KEYINPUT98), .A3(new_n270_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n270_), .A2(KEYINPUT92), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT92), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n267_), .A2(new_n280_), .A3(new_n269_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n214_), .A2(KEYINPUT24), .A3(new_n204_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n283_), .A2(new_n215_), .ZN(new_n284_));
  AND2_X1   g083(.A1(KEYINPUT79), .A2(G190gat), .ZN(new_n285_));
  NOR2_X1   g084(.A1(KEYINPUT79), .A2(G190gat), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT26), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT80), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT80), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n289_), .B(KEYINPUT26), .C1(new_n285_), .C2(new_n286_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n288_), .A2(new_n290_), .ZN(new_n291_));
  AND2_X1   g090(.A1(KEYINPUT78), .A2(G183gat), .ZN(new_n292_));
  NOR2_X1   g091(.A1(KEYINPUT78), .A2(G183gat), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT25), .ZN(new_n294_));
  NOR3_X1   g093(.A1(new_n292_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n222_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n284_), .B1(new_n291_), .B2(new_n297_), .ZN(new_n298_));
  OR2_X1    g097(.A1(KEYINPUT78), .A2(G183gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(KEYINPUT78), .A2(G183gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT79), .B(G190gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n228_), .A2(new_n229_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n235_), .A2(new_n237_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n298_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n279_), .A2(new_n281_), .A3(new_n309_), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n272_), .A2(KEYINPUT20), .A3(new_n278_), .A4(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G226gat), .A2(G233gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT19), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n311_), .A2(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G8gat), .B(G36gat), .ZN(new_n315_));
  INV_X1    g114(.A(G92gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(KEYINPUT18), .B(G64gat), .ZN(new_n318_));
  XOR2_X1   g117(.A(new_n317_), .B(new_n318_), .Z(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT20), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n279_), .A2(new_n281_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n321_), .B1(new_n322_), .B2(new_n308_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n313_), .B1(new_n250_), .B2(new_n271_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  AND3_X1   g124(.A1(new_n314_), .A2(new_n320_), .A3(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n320_), .B1(new_n314_), .B2(new_n325_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n202_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  AND3_X1   g127(.A1(new_n267_), .A2(new_n280_), .A3(new_n269_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n280_), .B1(new_n267_), .B2(new_n269_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n321_), .B1(new_n331_), .B2(new_n309_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n313_), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n332_), .A2(new_n333_), .A3(new_n272_), .A4(new_n278_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n308_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n271_), .A2(new_n274_), .A3(new_n243_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n335_), .A2(KEYINPUT20), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT101), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n337_), .A2(new_n338_), .A3(new_n313_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n334_), .A2(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n338_), .B1(new_n337_), .B2(new_n313_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n319_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  AOI22_X1  g141(.A1(new_n311_), .A2(new_n313_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n202_), .B1(new_n343_), .B2(new_n320_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n342_), .A2(new_n344_), .ZN(new_n345_));
  AND2_X1   g144(.A1(new_n328_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G225gat), .A2(G233gat), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT4), .ZN(new_n349_));
  INV_X1    g148(.A(G127gat), .ZN(new_n350_));
  INV_X1    g149(.A(G134gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G127gat), .A2(G134gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G113gat), .B(G120gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT82), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(G113gat), .ZN(new_n359_));
  INV_X1    g158(.A(G120gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G113gat), .A2(G120gat), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n352_), .A2(new_n361_), .A3(new_n353_), .A4(new_n362_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n363_), .A2(KEYINPUT83), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT83), .ZN(new_n365_));
  INV_X1    g164(.A(new_n353_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(G127gat), .A2(G134gat), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  AND2_X1   g167(.A1(G113gat), .A2(G120gat), .ZN(new_n369_));
  NOR2_X1   g168(.A1(G113gat), .A2(G120gat), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n365_), .B1(new_n368_), .B2(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n358_), .B1(new_n364_), .B2(new_n372_), .ZN(new_n373_));
  OR2_X1    g172(.A1(G155gat), .A2(G162gat), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT88), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G155gat), .A2(G162gat), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n374_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  AND2_X1   g176(.A1(G155gat), .A2(G162gat), .ZN(new_n378_));
  NOR2_X1   g177(.A1(G155gat), .A2(G162gat), .ZN(new_n379_));
  OAI21_X1  g178(.A(KEYINPUT88), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n377_), .A2(new_n380_), .ZN(new_n381_));
  OR3_X1    g180(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G141gat), .A2(G148gat), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT2), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n386_));
  NAND3_X1  g185(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n382_), .A2(new_n385_), .A3(new_n386_), .A4(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n381_), .A2(new_n388_), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT87), .B1(new_n376_), .B2(KEYINPUT1), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT87), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT1), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n391_), .A2(new_n392_), .A3(G155gat), .A4(G162gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n376_), .A2(KEYINPUT1), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n390_), .A2(new_n393_), .A3(new_n374_), .A4(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(KEYINPUT86), .B1(G141gat), .B2(G148gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(new_n383_), .ZN(new_n397_));
  NOR3_X1   g196(.A1(KEYINPUT86), .A2(G141gat), .A3(G148gat), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n395_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n389_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n363_), .A2(KEYINPUT83), .ZN(new_n402_));
  AOI21_X1  g201(.A(KEYINPUT82), .B1(new_n354_), .B2(new_n355_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n368_), .A2(new_n371_), .A3(new_n365_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n402_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n373_), .A2(new_n401_), .A3(new_n405_), .ZN(new_n406_));
  AOI22_X1  g205(.A1(new_n388_), .A2(new_n381_), .B1(new_n395_), .B2(new_n399_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n356_), .A2(new_n363_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n349_), .B1(new_n406_), .B2(new_n409_), .ZN(new_n410_));
  AND3_X1   g209(.A1(new_n402_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n403_), .B1(new_n402_), .B2(new_n404_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(KEYINPUT4), .B1(new_n413_), .B2(new_n401_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n348_), .B1(new_n410_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT99), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  OAI211_X1 g216(.A(KEYINPUT99), .B(new_n348_), .C1(new_n410_), .C2(new_n414_), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n406_), .A2(new_n409_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(new_n347_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n417_), .A2(new_n418_), .A3(new_n420_), .ZN(new_n421_));
  XOR2_X1   g220(.A(G1gat), .B(G29gat), .Z(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT100), .B(G85gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(KEYINPUT0), .B(G57gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n421_), .A2(new_n427_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n417_), .A2(new_n426_), .A3(new_n418_), .A4(new_n420_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(G228gat), .ZN(new_n431_));
  INV_X1    g230(.A(G233gat), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n434_), .A2(KEYINPUT89), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n331_), .A2(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(KEYINPUT89), .B1(new_n401_), .B2(KEYINPUT29), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT29), .ZN(new_n438_));
  OAI221_X1 g237(.A(new_n270_), .B1(new_n280_), .B2(new_n435_), .C1(new_n438_), .C2(new_n407_), .ZN(new_n439_));
  AOI22_X1  g238(.A1(new_n436_), .A2(new_n437_), .B1(new_n433_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(G50gat), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n389_), .A2(new_n400_), .A3(new_n438_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT28), .ZN(new_n443_));
  INV_X1    g242(.A(G22gat), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT28), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n389_), .A2(new_n400_), .A3(new_n445_), .A4(new_n438_), .ZN(new_n446_));
  AND3_X1   g245(.A1(new_n443_), .A2(new_n444_), .A3(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n444_), .B1(new_n443_), .B2(new_n446_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n441_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  XOR2_X1   g248(.A(G78gat), .B(G106gat), .Z(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT93), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n445_), .B1(new_n407_), .B2(new_n438_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n446_), .ZN(new_n454_));
  OAI21_X1  g253(.A(G22gat), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n443_), .A2(new_n444_), .A3(new_n446_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(G50gat), .A3(new_n456_), .ZN(new_n457_));
  AND3_X1   g256(.A1(new_n449_), .A2(new_n452_), .A3(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n450_), .B1(new_n449_), .B2(new_n457_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n440_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  NOR3_X1   g259(.A1(new_n447_), .A2(new_n448_), .A3(new_n441_), .ZN(new_n461_));
  AOI21_X1  g260(.A(G50gat), .B1(new_n455_), .B2(new_n456_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n451_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n322_), .B(new_n437_), .C1(KEYINPUT89), .C2(new_n434_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n439_), .A2(new_n433_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n449_), .A2(new_n452_), .A3(new_n457_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n463_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n460_), .A2(new_n468_), .ZN(new_n469_));
  XOR2_X1   g268(.A(new_n413_), .B(KEYINPUT31), .Z(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G227gat), .A2(G233gat), .ZN(new_n472_));
  INV_X1    g271(.A(G15gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(G43gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n472_), .B(G15gat), .ZN(new_n476_));
  INV_X1    g275(.A(G43gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n475_), .A2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(KEYINPUT81), .B(KEYINPUT30), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  XOR2_X1   g280(.A(G71gat), .B(G99gat), .Z(new_n482_));
  NAND3_X1  g281(.A1(new_n299_), .A2(KEYINPUT25), .A3(new_n300_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n296_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n485_), .A2(new_n288_), .A3(new_n222_), .A4(new_n290_), .ZN(new_n486_));
  AOI221_X4 g285(.A(new_n482_), .B1(new_n305_), .B2(new_n306_), .C1(new_n486_), .C2(new_n284_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n482_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n488_), .B1(new_n298_), .B2(new_n307_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n481_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n304_), .B(new_n282_), .C1(KEYINPUT24), .C2(new_n214_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n289_), .B1(new_n302_), .B2(KEYINPUT26), .ZN(new_n492_));
  INV_X1    g291(.A(new_n290_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  AOI22_X1  g293(.A1(new_n483_), .A2(new_n484_), .B1(new_n221_), .B2(G190gat), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n491_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n307_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n482_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n298_), .A2(new_n307_), .A3(new_n488_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n479_), .A2(new_n480_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n480_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n501_), .B1(new_n475_), .B2(new_n478_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n500_), .A2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n498_), .A2(new_n499_), .A3(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n490_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT84), .ZN(new_n506_));
  AOI21_X1  g305(.A(KEYINPUT85), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT85), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n508_), .B1(new_n490_), .B2(new_n504_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n471_), .B1(new_n507_), .B2(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(KEYINPUT84), .B1(new_n490_), .B2(new_n504_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n470_), .B1(new_n511_), .B2(KEYINPUT85), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n510_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n469_), .A2(new_n513_), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n460_), .A2(new_n510_), .A3(new_n468_), .A4(new_n512_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n430_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n320_), .A2(KEYINPUT32), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n518_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n343_), .A2(new_n517_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n519_), .A2(new_n430_), .A3(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n314_), .A2(new_n325_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(new_n319_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n419_), .A2(new_n348_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(new_n427_), .ZN(new_n525_));
  OR2_X1    g324(.A1(new_n410_), .A2(new_n414_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n525_), .B1(new_n347_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT33), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n527_), .B1(new_n429_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n343_), .A2(new_n320_), .ZN(new_n530_));
  AOI22_X1  g329(.A1(new_n415_), .A2(new_n416_), .B1(new_n347_), .B2(new_n419_), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n531_), .A2(KEYINPUT33), .A3(new_n426_), .A4(new_n418_), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n523_), .A2(new_n529_), .A3(new_n530_), .A4(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n521_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n513_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(new_n469_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  AOI22_X1  g336(.A1(new_n346_), .A2(new_n516_), .B1(new_n534_), .B2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n441_), .A2(G43gat), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n477_), .A2(G50gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(KEYINPUT70), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G43gat), .B(G50gat), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT70), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n542_), .A2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G29gat), .B(G36gat), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n546_), .A2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n542_), .A2(new_n545_), .A3(new_n547_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G15gat), .B(G22gat), .ZN(new_n553_));
  INV_X1    g352(.A(G1gat), .ZN(new_n554_));
  INV_X1    g353(.A(G8gat), .ZN(new_n555_));
  OAI21_X1  g354(.A(KEYINPUT14), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n553_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G1gat), .B(G8gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n552_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT15), .ZN(new_n561_));
  INV_X1    g360(.A(new_n550_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n547_), .B1(new_n542_), .B2(new_n545_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n561_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n549_), .A2(KEYINPUT15), .A3(new_n550_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n560_), .B1(new_n567_), .B2(new_n559_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G229gat), .A2(G233gat), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(new_n551_), .B(new_n559_), .Z(new_n571_));
  INV_X1    g370(.A(new_n569_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n570_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT77), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G113gat), .B(G141gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G169gat), .B(G197gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n574_), .A2(new_n575_), .A3(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n578_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G99gat), .A2(G106gat), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT6), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n586_));
  NAND2_X1  g385(.A1(G85gat), .A2(G92gat), .ZN(new_n587_));
  OAI211_X1 g386(.A(new_n585_), .B(new_n586_), .C1(KEYINPUT9), .C2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(G85gat), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(new_n316_), .ZN(new_n590_));
  AND3_X1   g389(.A1(new_n590_), .A2(KEYINPUT9), .A3(new_n587_), .ZN(new_n591_));
  INV_X1    g390(.A(G99gat), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(KEYINPUT10), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT10), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(G99gat), .ZN(new_n595_));
  AOI21_X1  g394(.A(G106gat), .B1(new_n593_), .B2(new_n595_), .ZN(new_n596_));
  OR3_X1    g395(.A1(new_n588_), .A2(new_n591_), .A3(new_n596_), .ZN(new_n597_));
  AND2_X1   g396(.A1(G85gat), .A2(G92gat), .ZN(new_n598_));
  NOR2_X1   g397(.A1(G85gat), .A2(G92gat), .ZN(new_n599_));
  OAI21_X1  g398(.A(KEYINPUT64), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT64), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n590_), .A2(new_n601_), .A3(new_n587_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT8), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT7), .ZN(new_n605_));
  INV_X1    g404(.A(G106gat), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n605_), .A2(new_n592_), .A3(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n607_), .A2(new_n585_), .A3(new_n586_), .A4(new_n608_), .ZN(new_n609_));
  AND3_X1   g408(.A1(new_n603_), .A2(new_n604_), .A3(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n604_), .B1(new_n603_), .B2(new_n609_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n597_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT65), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  OAI211_X1 g413(.A(KEYINPUT65), .B(new_n597_), .C1(new_n610_), .C2(new_n611_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(new_n567_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(G232gat), .A2(G233gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT34), .ZN(new_n619_));
  OAI22_X1  g418(.A1(new_n552_), .A2(new_n612_), .B1(KEYINPUT35), .B2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(KEYINPUT35), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT69), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n617_), .A2(new_n621_), .A3(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n566_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n623_), .B1(new_n626_), .B2(new_n620_), .ZN(new_n627_));
  XOR2_X1   g426(.A(G190gat), .B(G218gat), .Z(new_n628_));
  XNOR2_X1  g427(.A(G134gat), .B(G162gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n628_), .B(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT36), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT71), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n625_), .A2(new_n627_), .A3(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT37), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n625_), .A2(new_n627_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n630_), .B(KEYINPUT36), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n637_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(KEYINPUT72), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT72), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n638_), .A2(new_n643_), .A3(new_n639_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n635_), .B1(new_n642_), .B2(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n641_), .B1(new_n645_), .B2(KEYINPUT37), .ZN(new_n646_));
  XNOR2_X1  g445(.A(G57gat), .B(G64gat), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n647_), .A2(KEYINPUT11), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(KEYINPUT11), .ZN(new_n649_));
  XOR2_X1   g448(.A(G71gat), .B(G78gat), .Z(new_n650_));
  NAND3_X1  g449(.A1(new_n648_), .A2(new_n649_), .A3(new_n650_), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n649_), .A2(new_n650_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT12), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n651_), .A2(new_n652_), .ZN(new_n656_));
  AOI21_X1  g455(.A(KEYINPUT12), .B1(new_n612_), .B2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT66), .ZN(new_n658_));
  AOI22_X1  g457(.A1(new_n616_), .A2(new_n655_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(G230gat), .A2(G233gat), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n588_), .A2(new_n591_), .A3(new_n596_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n598_), .A2(new_n599_), .A3(KEYINPUT64), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n601_), .B1(new_n590_), .B2(new_n587_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n609_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(KEYINPUT8), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n603_), .A2(new_n604_), .A3(new_n609_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n661_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n654_), .B1(new_n667_), .B2(new_n653_), .ZN(new_n668_));
  AOI22_X1  g467(.A1(new_n668_), .A2(KEYINPUT66), .B1(new_n667_), .B2(new_n653_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n659_), .A2(new_n660_), .A3(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n667_), .A2(new_n653_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n612_), .A2(new_n656_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n660_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n670_), .A2(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(G120gat), .B(G148gat), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT68), .ZN(new_n678_));
  XOR2_X1   g477(.A(new_n678_), .B(KEYINPUT67), .Z(new_n679_));
  XOR2_X1   g478(.A(G176gat), .B(G204gat), .Z(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT5), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n679_), .B(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n676_), .A2(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n670_), .A2(new_n675_), .A3(new_n682_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT13), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n684_), .A2(KEYINPUT13), .A3(new_n685_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n646_), .A2(new_n690_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(G183gat), .B(G211gat), .ZN(new_n692_));
  XNOR2_X1  g491(.A(G127gat), .B(G155gat), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n692_), .B(new_n693_), .Z(new_n694_));
  NAND2_X1  g493(.A1(G231gat), .A2(G233gat), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT73), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n559_), .B(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(new_n656_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT75), .ZN(new_n699_));
  XNOR2_X1  g498(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n698_), .A2(new_n699_), .A3(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n701_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n694_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n704_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n694_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n706_), .A2(new_n702_), .A3(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n705_), .A2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(KEYINPUT17), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT17), .ZN(new_n711_));
  NAND4_X1  g510(.A1(new_n705_), .A2(new_n708_), .A3(new_n711_), .A4(new_n698_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n691_), .A2(new_n714_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n582_), .B1(new_n715_), .B2(KEYINPUT76), .ZN(new_n716_));
  AOI211_X1 g515(.A(new_n538_), .B(new_n716_), .C1(KEYINPUT76), .C2(new_n715_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n717_), .A2(new_n554_), .A3(new_n430_), .ZN(new_n718_));
  XOR2_X1   g517(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n718_), .A2(new_n720_), .ZN(new_n721_));
  OR2_X1    g520(.A1(new_n721_), .A2(KEYINPUT103), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(KEYINPUT103), .ZN(new_n723_));
  INV_X1    g522(.A(new_n690_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(new_n582_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n538_), .A2(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n645_), .B(KEYINPUT104), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n727_), .A2(new_n713_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n726_), .A2(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n554_), .B1(new_n729_), .B2(new_n430_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n730_), .B1(new_n718_), .B2(new_n720_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n722_), .A2(new_n723_), .A3(new_n731_), .ZN(G1324gat));
  NAND2_X1  g531(.A1(new_n328_), .A2(new_n345_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n555_), .B1(new_n729_), .B2(new_n733_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT39), .Z(new_n735_));
  NAND3_X1  g534(.A1(new_n717_), .A2(new_n555_), .A3(new_n733_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n737_), .B(KEYINPUT40), .Z(G1325gat));
  NAND2_X1  g537(.A1(new_n729_), .A2(new_n513_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(G15gat), .ZN(new_n740_));
  OR2_X1    g539(.A1(new_n740_), .A2(KEYINPUT41), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(KEYINPUT41), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n717_), .A2(new_n473_), .A3(new_n513_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n741_), .A2(new_n742_), .A3(new_n743_), .ZN(new_n744_));
  XOR2_X1   g543(.A(new_n744_), .B(KEYINPUT105), .Z(G1326gat));
  INV_X1    g544(.A(new_n469_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n444_), .B1(new_n729_), .B2(new_n746_), .ZN(new_n747_));
  XOR2_X1   g546(.A(new_n747_), .B(KEYINPUT42), .Z(new_n748_));
  NAND3_X1  g547(.A1(new_n717_), .A2(new_n444_), .A3(new_n746_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(G1327gat));
  NOR2_X1   g549(.A1(new_n725_), .A2(new_n714_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT43), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n752_), .B1(new_n646_), .B2(KEYINPUT106), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n638_), .A2(new_n643_), .A3(new_n639_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n643_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n634_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  AOI22_X1  g555(.A1(new_n756_), .A2(new_n636_), .B1(new_n640_), .B2(new_n637_), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n538_), .A2(new_n753_), .A3(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT106), .ZN(new_n759_));
  OAI21_X1  g558(.A(KEYINPUT43), .B1(new_n757_), .B2(new_n759_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n529_), .A2(new_n532_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n326_), .A2(new_n327_), .ZN(new_n762_));
  AOI22_X1  g561(.A1(new_n428_), .A2(new_n429_), .B1(new_n343_), .B2(new_n517_), .ZN(new_n763_));
  AOI22_X1  g562(.A1(new_n761_), .A2(new_n762_), .B1(new_n519_), .B2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n430_), .ZN(new_n765_));
  AND4_X1   g564(.A1(new_n460_), .A2(new_n510_), .A3(new_n468_), .A4(new_n512_), .ZN(new_n766_));
  AOI22_X1  g565(.A1(new_n460_), .A2(new_n468_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n765_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  OAI22_X1  g567(.A1(new_n764_), .A2(new_n536_), .B1(new_n768_), .B2(new_n733_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n760_), .B1(new_n769_), .B2(new_n646_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n751_), .B1(new_n758_), .B2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT44), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  OAI211_X1 g572(.A(KEYINPUT44), .B(new_n751_), .C1(new_n758_), .C2(new_n770_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(G29gat), .B1(new_n775_), .B2(new_n765_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n714_), .A2(new_n756_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n726_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(G29gat), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n778_), .A2(new_n779_), .A3(new_n430_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n776_), .A2(new_n780_), .ZN(G1328gat));
  INV_X1    g580(.A(G36gat), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n778_), .A2(new_n782_), .A3(new_n733_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT45), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n773_), .A2(new_n733_), .A3(new_n774_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT107), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT107), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n773_), .A2(new_n787_), .A3(new_n733_), .A4(new_n774_), .ZN(new_n788_));
  AND4_X1   g587(.A1(KEYINPUT108), .A2(new_n786_), .A3(G36gat), .A4(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n782_), .B1(new_n785_), .B2(KEYINPUT107), .ZN(new_n790_));
  AOI21_X1  g589(.A(KEYINPUT108), .B1(new_n790_), .B2(new_n788_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n784_), .B1(new_n789_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT46), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  OAI211_X1 g593(.A(KEYINPUT46), .B(new_n784_), .C1(new_n789_), .C2(new_n791_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(G1329gat));
  NAND3_X1  g595(.A1(new_n773_), .A2(new_n513_), .A3(new_n774_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n535_), .A2(G43gat), .ZN(new_n798_));
  AOI22_X1  g597(.A1(new_n797_), .A2(G43gat), .B1(new_n778_), .B2(new_n798_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n799_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g599(.A(G50gat), .B1(new_n775_), .B2(new_n469_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n746_), .A2(new_n441_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(KEYINPUT109), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n778_), .A2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n801_), .A2(new_n804_), .ZN(G1331gat));
  NOR3_X1   g604(.A1(new_n538_), .A2(new_n724_), .A3(new_n582_), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n806_), .A2(new_n757_), .A3(new_n714_), .ZN(new_n807_));
  AOI21_X1  g606(.A(G57gat), .B1(new_n807_), .B2(new_n430_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n728_), .ZN(new_n809_));
  XOR2_X1   g608(.A(new_n809_), .B(KEYINPUT110), .Z(new_n810_));
  AND2_X1   g609(.A1(new_n430_), .A2(G57gat), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n808_), .B1(new_n810_), .B2(new_n811_), .ZN(G1332gat));
  INV_X1    g611(.A(G64gat), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n813_), .B1(new_n810_), .B2(new_n733_), .ZN(new_n814_));
  XOR2_X1   g613(.A(new_n814_), .B(KEYINPUT48), .Z(new_n815_));
  NAND3_X1  g614(.A1(new_n807_), .A2(new_n813_), .A3(new_n733_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(G1333gat));
  INV_X1    g616(.A(G71gat), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n818_), .B1(new_n810_), .B2(new_n513_), .ZN(new_n819_));
  XOR2_X1   g618(.A(new_n819_), .B(KEYINPUT49), .Z(new_n820_));
  NAND3_X1  g619(.A1(new_n807_), .A2(new_n818_), .A3(new_n513_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(G1334gat));
  INV_X1    g621(.A(G78gat), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n823_), .B1(new_n810_), .B2(new_n746_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n824_), .B(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n807_), .A2(new_n823_), .A3(new_n746_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(G1335gat));
  NAND2_X1  g627(.A1(new_n806_), .A2(new_n777_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n829_), .B(KEYINPUT112), .ZN(new_n830_));
  AOI21_X1  g629(.A(G85gat), .B1(new_n830_), .B2(new_n430_), .ZN(new_n831_));
  XNOR2_X1  g630(.A(new_n831_), .B(KEYINPUT113), .ZN(new_n832_));
  OR2_X1    g631(.A1(new_n758_), .A2(new_n770_), .ZN(new_n833_));
  NOR3_X1   g632(.A1(new_n714_), .A2(new_n724_), .A3(new_n582_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n430_), .A2(G85gat), .ZN(new_n836_));
  XOR2_X1   g635(.A(new_n836_), .B(KEYINPUT114), .Z(new_n837_));
  AOI21_X1  g636(.A(new_n832_), .B1(new_n835_), .B2(new_n837_), .ZN(G1336gat));
  AOI21_X1  g637(.A(G92gat), .B1(new_n830_), .B2(new_n733_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n346_), .A2(new_n316_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n839_), .B1(new_n835_), .B2(new_n840_), .ZN(G1337gat));
  NAND2_X1  g640(.A1(new_n593_), .A2(new_n595_), .ZN(new_n842_));
  AND3_X1   g641(.A1(new_n830_), .A2(new_n842_), .A3(new_n513_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n592_), .B1(new_n835_), .B2(new_n513_), .ZN(new_n844_));
  OAI22_X1  g643(.A1(new_n843_), .A2(new_n844_), .B1(KEYINPUT115), .B2(KEYINPUT51), .ZN(new_n845_));
  NAND2_X1  g644(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n845_), .B(new_n846_), .ZN(G1338gat));
  NAND3_X1  g646(.A1(new_n833_), .A2(new_n746_), .A3(new_n834_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(KEYINPUT116), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT116), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n833_), .A2(new_n850_), .A3(new_n746_), .A4(new_n834_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n849_), .A2(G106gat), .A3(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(KEYINPUT52), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n849_), .A2(new_n854_), .A3(G106gat), .A4(new_n851_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n469_), .A2(G106gat), .ZN(new_n856_));
  AOI22_X1  g655(.A1(new_n853_), .A2(new_n855_), .B1(new_n830_), .B2(new_n856_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n857_), .B(new_n859_), .ZN(G1339gat));
  INV_X1    g659(.A(KEYINPUT55), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n667_), .A2(KEYINPUT65), .ZN(new_n862_));
  AOI211_X1 g661(.A(new_n613_), .B(new_n661_), .C1(new_n665_), .C2(new_n666_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n655_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n668_), .A2(KEYINPUT66), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n672_), .A2(new_n658_), .A3(new_n654_), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n864_), .A2(new_n865_), .A3(new_n671_), .A4(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n861_), .B1(new_n867_), .B2(new_n674_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n867_), .A2(new_n674_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n659_), .A2(KEYINPUT55), .A3(new_n660_), .A4(new_n669_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n683_), .B1(new_n870_), .B2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(KEYINPUT56), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n574_), .A2(new_n578_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n571_), .A2(new_n569_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n578_), .ZN(new_n877_));
  OR2_X1    g676(.A1(new_n877_), .A2(KEYINPUT119), .ZN(new_n878_));
  AOI22_X1  g677(.A1(new_n877_), .A2(KEYINPUT119), .B1(new_n572_), .B2(new_n568_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n875_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n660_), .B1(new_n659_), .B2(new_n669_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n670_), .B1(new_n881_), .B2(new_n861_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n682_), .B1(new_n882_), .B2(new_n871_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT56), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  NAND4_X1  g684(.A1(new_n874_), .A2(new_n880_), .A3(new_n685_), .A4(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT58), .ZN(new_n887_));
  OAI21_X1  g686(.A(KEYINPUT120), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n757_), .B1(new_n886_), .B2(new_n887_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n685_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n890_));
  AOI211_X1 g689(.A(KEYINPUT56), .B(new_n682_), .C1(new_n882_), .C2(new_n871_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT120), .ZN(new_n893_));
  NAND4_X1  g692(.A1(new_n892_), .A2(new_n893_), .A3(KEYINPUT58), .A4(new_n880_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n888_), .A2(new_n889_), .A3(new_n894_), .ZN(new_n895_));
  NOR3_X1   g694(.A1(new_n890_), .A2(new_n581_), .A3(new_n891_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n880_), .A2(new_n686_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n756_), .B1(new_n896_), .B2(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT57), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  NAND4_X1  g700(.A1(new_n874_), .A2(new_n582_), .A3(new_n685_), .A4(new_n885_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(new_n897_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n903_), .A2(KEYINPUT57), .A3(new_n756_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n895_), .A2(new_n901_), .A3(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(new_n713_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n710_), .A2(new_n712_), .A3(new_n581_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(KEYINPUT118), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT118), .ZN(new_n909_));
  NAND4_X1  g708(.A1(new_n710_), .A2(new_n712_), .A3(new_n581_), .A4(new_n909_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n908_), .A2(new_n691_), .A3(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT54), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(new_n913_));
  NAND4_X1  g712(.A1(new_n908_), .A2(new_n691_), .A3(KEYINPUT54), .A4(new_n910_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n906_), .A2(new_n916_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n733_), .A2(new_n765_), .ZN(new_n918_));
  AND2_X1   g717(.A1(new_n917_), .A2(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(new_n767_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n920_), .ZN(new_n921_));
  AOI21_X1  g720(.A(G113gat), .B1(new_n921_), .B2(new_n582_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n920_), .A2(KEYINPUT59), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n917_), .A2(new_n918_), .ZN(new_n924_));
  OR3_X1    g723(.A1(new_n924_), .A2(KEYINPUT59), .A3(new_n514_), .ZN(new_n925_));
  AND2_X1   g724(.A1(new_n923_), .A2(new_n925_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n581_), .A2(new_n359_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n922_), .B1(new_n926_), .B2(new_n927_), .ZN(G1340gat));
  NAND3_X1  g727(.A1(new_n923_), .A2(new_n690_), .A3(new_n925_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(G120gat), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n360_), .B1(new_n724_), .B2(KEYINPUT60), .ZN(new_n931_));
  OAI211_X1 g730(.A(new_n921_), .B(new_n931_), .C1(KEYINPUT60), .C2(new_n360_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n930_), .A2(new_n932_), .ZN(G1341gat));
  NAND2_X1  g732(.A1(new_n714_), .A2(G127gat), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n934_), .B(KEYINPUT122), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n350_), .B1(new_n920_), .B2(new_n713_), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT121), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n936_), .A2(new_n937_), .ZN(new_n938_));
  OAI211_X1 g737(.A(KEYINPUT121), .B(new_n350_), .C1(new_n920_), .C2(new_n713_), .ZN(new_n939_));
  AOI22_X1  g738(.A1(new_n926_), .A2(new_n935_), .B1(new_n938_), .B2(new_n939_), .ZN(G1342gat));
  AOI21_X1  g739(.A(G134gat), .B1(new_n921_), .B2(new_n727_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n757_), .A2(new_n351_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n941_), .B1(new_n926_), .B2(new_n942_), .ZN(G1343gat));
  NOR2_X1   g742(.A1(new_n924_), .A2(new_n515_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n944_), .A2(new_n582_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(new_n945_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g745(.A1(new_n944_), .A2(new_n690_), .ZN(new_n947_));
  XNOR2_X1  g746(.A(new_n947_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g747(.A1(new_n944_), .A2(new_n714_), .ZN(new_n949_));
  XNOR2_X1  g748(.A(KEYINPUT61), .B(G155gat), .ZN(new_n950_));
  XNOR2_X1  g749(.A(new_n949_), .B(new_n950_), .ZN(G1346gat));
  AOI21_X1  g750(.A(G162gat), .B1(new_n944_), .B2(new_n727_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n646_), .A2(G162gat), .ZN(new_n953_));
  XNOR2_X1  g752(.A(new_n953_), .B(KEYINPUT123), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n952_), .B1(new_n944_), .B2(new_n954_), .ZN(G1347gat));
  NOR2_X1   g754(.A1(new_n346_), .A2(new_n430_), .ZN(new_n956_));
  AOI21_X1  g755(.A(KEYINPUT57), .B1(new_n903_), .B2(new_n756_), .ZN(new_n957_));
  AOI211_X1 g756(.A(new_n900_), .B(new_n645_), .C1(new_n902_), .C2(new_n897_), .ZN(new_n958_));
  NOR2_X1   g757(.A1(new_n957_), .A2(new_n958_), .ZN(new_n959_));
  AOI21_X1  g758(.A(new_n714_), .B1(new_n959_), .B2(new_n895_), .ZN(new_n960_));
  OAI211_X1 g759(.A(new_n767_), .B(new_n956_), .C1(new_n960_), .C2(new_n915_), .ZN(new_n961_));
  OAI21_X1  g760(.A(G169gat), .B1(new_n961_), .B2(new_n581_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n962_), .A2(KEYINPUT124), .ZN(new_n963_));
  INV_X1    g762(.A(KEYINPUT124), .ZN(new_n964_));
  OAI211_X1 g763(.A(new_n964_), .B(G169gat), .C1(new_n961_), .C2(new_n581_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n963_), .A2(new_n965_), .ZN(new_n966_));
  INV_X1    g765(.A(KEYINPUT62), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n966_), .A2(new_n967_), .ZN(new_n968_));
  INV_X1    g767(.A(KEYINPUT125), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n961_), .A2(new_n969_), .ZN(new_n970_));
  NAND4_X1  g769(.A1(new_n917_), .A2(KEYINPUT125), .A3(new_n767_), .A4(new_n956_), .ZN(new_n971_));
  AOI21_X1  g770(.A(new_n581_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n972_));
  NAND3_X1  g771(.A1(new_n970_), .A2(new_n971_), .A3(new_n972_), .ZN(new_n973_));
  NAND3_X1  g772(.A1(new_n963_), .A2(KEYINPUT62), .A3(new_n965_), .ZN(new_n974_));
  NAND3_X1  g773(.A1(new_n968_), .A2(new_n973_), .A3(new_n974_), .ZN(G1348gat));
  NOR3_X1   g774(.A1(new_n961_), .A2(new_n207_), .A3(new_n724_), .ZN(new_n976_));
  NAND3_X1  g775(.A1(new_n970_), .A2(new_n690_), .A3(new_n971_), .ZN(new_n977_));
  AOI21_X1  g776(.A(new_n976_), .B1(new_n977_), .B2(new_n207_), .ZN(G1349gat));
  NAND4_X1  g777(.A1(new_n970_), .A2(new_n714_), .A3(new_n971_), .A4(new_n218_), .ZN(new_n979_));
  OAI21_X1  g778(.A(new_n301_), .B1(new_n961_), .B2(new_n713_), .ZN(new_n980_));
  AND2_X1   g779(.A1(new_n979_), .A2(new_n980_), .ZN(G1350gat));
  NAND3_X1  g780(.A1(new_n970_), .A2(new_n646_), .A3(new_n971_), .ZN(new_n982_));
  NAND2_X1  g781(.A1(new_n982_), .A2(G190gat), .ZN(new_n983_));
  INV_X1    g782(.A(new_n727_), .ZN(new_n984_));
  NOR2_X1   g783(.A1(new_n984_), .A2(new_n273_), .ZN(new_n985_));
  XNOR2_X1  g784(.A(new_n985_), .B(KEYINPUT126), .ZN(new_n986_));
  NAND3_X1  g785(.A1(new_n970_), .A2(new_n971_), .A3(new_n986_), .ZN(new_n987_));
  NAND2_X1  g786(.A1(new_n983_), .A2(new_n987_), .ZN(new_n988_));
  NAND2_X1  g787(.A1(new_n988_), .A2(KEYINPUT127), .ZN(new_n989_));
  INV_X1    g788(.A(KEYINPUT127), .ZN(new_n990_));
  NAND3_X1  g789(.A1(new_n983_), .A2(new_n990_), .A3(new_n987_), .ZN(new_n991_));
  NAND2_X1  g790(.A1(new_n989_), .A2(new_n991_), .ZN(G1351gat));
  AND2_X1   g791(.A1(new_n917_), .A2(new_n956_), .ZN(new_n993_));
  NAND2_X1  g792(.A1(new_n993_), .A2(new_n766_), .ZN(new_n994_));
  NOR2_X1   g793(.A1(new_n994_), .A2(new_n581_), .ZN(new_n995_));
  XNOR2_X1  g794(.A(new_n995_), .B(new_n252_), .ZN(G1352gat));
  INV_X1    g795(.A(new_n994_), .ZN(new_n997_));
  NAND2_X1  g796(.A1(new_n997_), .A2(new_n690_), .ZN(new_n998_));
  NAND2_X1  g797(.A1(new_n998_), .A2(G204gat), .ZN(new_n999_));
  OAI21_X1  g798(.A(new_n999_), .B1(new_n998_), .B2(new_n254_), .ZN(G1353gat));
  NOR2_X1   g799(.A1(new_n994_), .A2(new_n713_), .ZN(new_n1001_));
  NOR2_X1   g800(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1002_));
  AND2_X1   g801(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1003_));
  OAI21_X1  g802(.A(new_n1001_), .B1(new_n1002_), .B2(new_n1003_), .ZN(new_n1004_));
  OAI21_X1  g803(.A(new_n1004_), .B1(new_n1001_), .B2(new_n1002_), .ZN(G1354gat));
  AND3_X1   g804(.A1(new_n997_), .A2(G218gat), .A3(new_n646_), .ZN(new_n1006_));
  AOI21_X1  g805(.A(G218gat), .B1(new_n997_), .B2(new_n727_), .ZN(new_n1007_));
  NOR2_X1   g806(.A1(new_n1006_), .A2(new_n1007_), .ZN(G1355gat));
endmodule


