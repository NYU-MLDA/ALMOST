//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 0 0 0 0 1 1 0 0 1 1 1 1 0 1 0 0 1 1 1 1 1 1 0 0 0 0 1 1 1 1 0 1 1 0 0 1 1 1 1 0 1 0 0 0 0 1 0 0 0 0 0 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n741_, new_n742_, new_n743_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n754_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n832_, new_n833_, new_n835_, new_n836_, new_n837_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n845_, new_n846_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n871_, new_n872_, new_n873_, new_n875_, new_n876_,
    new_n877_, new_n879_, new_n880_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_;
  INV_X1    g000(.A(KEYINPUT12), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G99gat), .A2(G106gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT6), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(KEYINPUT10), .B(G99gat), .Z(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT65), .ZN(new_n207_));
  INV_X1    g006(.A(G106gat), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n205_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT9), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT66), .B(G92gat), .ZN(new_n211_));
  INV_X1    g010(.A(G85gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n210_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT67), .ZN(new_n216_));
  OR2_X1    g015(.A1(G85gat), .A2(G92gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT67), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(new_n214_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n216_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n209_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G85gat), .A2(G92gat), .ZN(new_n222_));
  NOR2_X1   g021(.A1(G99gat), .A2(G106gat), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT7), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n223_), .B(new_n224_), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n217_), .B(new_n222_), .C1(new_n225_), .C2(new_n205_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT8), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n221_), .A2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G57gat), .B(G64gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT11), .ZN(new_n230_));
  XOR2_X1   g029(.A(G71gat), .B(G78gat), .Z(new_n231_));
  OR2_X1    g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n230_), .A2(new_n231_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n229_), .A2(KEYINPUT11), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n232_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n202_), .B1(new_n228_), .B2(new_n235_), .ZN(new_n236_));
  OR2_X1    g035(.A1(new_n235_), .A2(new_n202_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT68), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n227_), .B1(new_n221_), .B2(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(KEYINPUT68), .B1(new_n209_), .B2(new_n220_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n238_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G230gat), .A2(G233gat), .ZN(new_n243_));
  XOR2_X1   g042(.A(new_n243_), .B(KEYINPUT64), .Z(new_n244_));
  NAND2_X1  g043(.A1(new_n228_), .A2(new_n235_), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n236_), .A2(new_n242_), .A3(new_n244_), .A4(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n244_), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n228_), .A2(new_n235_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n228_), .A2(new_n235_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n247_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  XOR2_X1   g049(.A(G120gat), .B(G148gat), .Z(new_n251_));
  XNOR2_X1  g050(.A(G176gat), .B(G204gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n253_), .B(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n246_), .A2(new_n250_), .A3(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT71), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n246_), .A2(new_n250_), .A3(KEYINPUT71), .A4(new_n255_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n246_), .A2(new_n250_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n255_), .B(KEYINPUT70), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n260_), .A2(new_n263_), .ZN(new_n264_));
  XOR2_X1   g063(.A(KEYINPUT72), .B(KEYINPUT13), .Z(new_n265_));
  NOR2_X1   g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n267_), .B1(new_n260_), .B2(new_n263_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n266_), .A2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G29gat), .B(G36gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT73), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G43gat), .B(G50gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT15), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n274_), .B1(new_n241_), .B2(new_n240_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G232gat), .A2(G233gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT34), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT35), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  AOI22_X1  g080(.A1(new_n228_), .A2(new_n273_), .B1(new_n279_), .B2(new_n278_), .ZN(new_n282_));
  AND3_X1   g081(.A1(new_n275_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n281_), .B1(new_n275_), .B2(new_n282_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G190gat), .B(G218gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G134gat), .B(G162gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  OR2_X1    g086(.A1(new_n287_), .A2(KEYINPUT36), .ZN(new_n288_));
  OR3_X1    g087(.A1(new_n283_), .A2(new_n284_), .A3(new_n288_), .ZN(new_n289_));
  XOR2_X1   g088(.A(new_n287_), .B(KEYINPUT36), .Z(new_n290_));
  OAI21_X1  g089(.A(new_n290_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n289_), .A2(KEYINPUT37), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT74), .ZN(new_n294_));
  OR2_X1    g093(.A1(new_n291_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n291_), .A2(new_n294_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n295_), .A2(new_n296_), .A3(new_n289_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT37), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n293_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT76), .B(G1gat), .ZN(new_n301_));
  INV_X1    g100(.A(G8gat), .ZN(new_n302_));
  OAI21_X1  g101(.A(KEYINPUT14), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT77), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT75), .B(G15gat), .ZN(new_n305_));
  INV_X1    g104(.A(G22gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n304_), .A2(new_n307_), .ZN(new_n308_));
  XOR2_X1   g107(.A(G1gat), .B(G8gat), .Z(new_n309_));
  OR2_X1    g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n309_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G231gat), .A2(G233gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT78), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n312_), .B(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(new_n235_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G127gat), .B(G155gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT16), .ZN(new_n318_));
  XOR2_X1   g117(.A(G183gat), .B(G211gat), .Z(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT17), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n316_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT17), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n320_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n322_), .B1(new_n325_), .B2(new_n316_), .ZN(new_n326_));
  NOR3_X1   g125(.A1(new_n269_), .A2(new_n300_), .A3(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n274_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT79), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G229gat), .A2(G233gat), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n308_), .A2(new_n309_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n308_), .A2(new_n309_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n273_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n328_), .A2(new_n329_), .A3(new_n330_), .A4(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT15), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n273_), .B(new_n335_), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n333_), .B(new_n330_), .C1(new_n312_), .C2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT79), .ZN(new_n338_));
  INV_X1    g137(.A(new_n273_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n310_), .A2(new_n339_), .A3(new_n311_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n330_), .B1(new_n333_), .B2(new_n340_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n334_), .B1(new_n338_), .B2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G113gat), .B(G141gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G169gat), .B(G197gat), .ZN(new_n344_));
  XOR2_X1   g143(.A(new_n343_), .B(new_n344_), .Z(new_n345_));
  NAND2_X1  g144(.A1(new_n342_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n333_), .A2(new_n340_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n330_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n349_), .A2(KEYINPUT79), .A3(new_n337_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n345_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n350_), .A2(new_n334_), .A3(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n346_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT80), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT25), .B(G183gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT26), .B(G190gat), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G169gat), .A2(G176gat), .ZN(new_n360_));
  AOI22_X1  g159(.A1(new_n356_), .A2(new_n357_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G183gat), .A2(G190gat), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT23), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NOR3_X1   g165(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n361_), .A2(new_n368_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(G169gat), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n364_), .B(new_n365_), .C1(G183gat), .C2(G190gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n369_), .A2(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G71gat), .B(G99gat), .ZN(new_n375_));
  INV_X1    g174(.A(G43gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n374_), .A2(new_n377_), .ZN(new_n378_));
  AOI22_X1  g177(.A1(new_n361_), .A2(new_n368_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n377_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G227gat), .A2(G233gat), .ZN(new_n382_));
  XOR2_X1   g181(.A(new_n382_), .B(G15gat), .Z(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(KEYINPUT30), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  OR3_X1    g184(.A1(new_n378_), .A2(new_n381_), .A3(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n385_), .B1(new_n378_), .B2(new_n381_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n355_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  XOR2_X1   g187(.A(G127gat), .B(G134gat), .Z(new_n389_));
  XOR2_X1   g188(.A(G113gat), .B(G120gat), .Z(new_n390_));
  XOR2_X1   g189(.A(new_n389_), .B(new_n390_), .Z(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT31), .ZN(new_n392_));
  NOR3_X1   g191(.A1(new_n388_), .A2(KEYINPUT81), .A3(new_n392_), .ZN(new_n393_));
  OR2_X1    g192(.A1(new_n388_), .A2(KEYINPUT81), .ZN(new_n394_));
  INV_X1    g193(.A(new_n392_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n386_), .A2(new_n387_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n395_), .B1(new_n396_), .B2(KEYINPUT81), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n393_), .B1(new_n394_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(G204gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(G197gat), .ZN(new_n401_));
  INV_X1    g200(.A(G197gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(G204gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(KEYINPUT21), .ZN(new_n405_));
  INV_X1    g204(.A(G218gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(G211gat), .ZN(new_n407_));
  INV_X1    g206(.A(G211gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(G218gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT86), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n412_), .B1(new_n402_), .B2(G204gat), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n400_), .A2(KEYINPUT86), .A3(G197gat), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n413_), .A2(new_n403_), .A3(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(KEYINPUT87), .B(KEYINPUT21), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n405_), .B(new_n411_), .C1(new_n415_), .C2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT21), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n418_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT88), .ZN(new_n420_));
  AND3_X1   g219(.A1(new_n415_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n420_), .B1(new_n415_), .B2(new_n419_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n417_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(G155gat), .ZN(new_n424_));
  INV_X1    g223(.A(G162gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G155gat), .A2(G162gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(KEYINPUT82), .A2(G141gat), .A3(G148gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT85), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT2), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G141gat), .A2(G148gat), .ZN(new_n433_));
  AND2_X1   g232(.A1(KEYINPUT85), .A2(KEYINPUT2), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT82), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n433_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n432_), .A2(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(G141gat), .A2(G148gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(KEYINPUT3), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n428_), .B1(new_n437_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT84), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT1), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n442_), .A2(G155gat), .A3(G162gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(new_n426_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n427_), .A2(KEYINPUT1), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT83), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n427_), .A2(KEYINPUT83), .A3(KEYINPUT1), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n444_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(KEYINPUT82), .B1(G141gat), .B2(G148gat), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n450_), .A2(new_n438_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(new_n429_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n441_), .B1(new_n449_), .B2(new_n452_), .ZN(new_n453_));
  AND3_X1   g252(.A1(new_n427_), .A2(KEYINPUT83), .A3(KEYINPUT1), .ZN(new_n454_));
  AOI21_X1  g253(.A(KEYINPUT83), .B1(new_n427_), .B2(KEYINPUT1), .ZN(new_n455_));
  OAI211_X1 g254(.A(new_n426_), .B(new_n443_), .C1(new_n454_), .C2(new_n455_), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n451_), .A2(new_n429_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n456_), .A2(new_n457_), .A3(KEYINPUT84), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n440_), .B1(new_n453_), .B2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT29), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n423_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n461_), .A2(G228gat), .A3(G233gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G228gat), .A2(G233gat), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n463_), .B(new_n423_), .C1(new_n459_), .C2(new_n460_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G78gat), .B(G106gat), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n462_), .A2(new_n464_), .A3(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT89), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n459_), .A2(new_n460_), .ZN(new_n470_));
  XOR2_X1   g269(.A(G22gat), .B(G50gat), .Z(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT28), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n470_), .B(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n469_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n462_), .A2(new_n464_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(new_n465_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(new_n467_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n474_), .A2(new_n477_), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n476_), .A2(KEYINPUT89), .A3(new_n467_), .A4(new_n473_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n437_), .A2(new_n439_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n428_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NOR3_X1   g283(.A1(new_n449_), .A2(new_n441_), .A3(new_n452_), .ZN(new_n485_));
  AOI21_X1  g284(.A(KEYINPUT84), .B1(new_n456_), .B2(new_n457_), .ZN(new_n486_));
  OAI211_X1 g285(.A(KEYINPUT90), .B(new_n484_), .C1(new_n485_), .C2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n391_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n391_), .B1(new_n459_), .B2(KEYINPUT90), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT4), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G225gat), .A2(G233gat), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT4), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n391_), .A2(new_n494_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n493_), .B1(new_n459_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n491_), .A2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G1gat), .B(G29gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(KEYINPUT91), .B(G85gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(KEYINPUT0), .B(G57gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n487_), .A2(new_n488_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n459_), .A2(KEYINPUT90), .A3(new_n391_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n504_), .B1(new_n507_), .B2(new_n492_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n498_), .A2(KEYINPUT33), .A3(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G8gat), .B(G36gat), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT18), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G64gat), .B(G92gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT20), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n515_), .B1(new_n423_), .B2(new_n374_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G226gat), .A2(G233gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT19), .ZN(new_n518_));
  OAI211_X1 g317(.A(new_n379_), .B(new_n417_), .C1(new_n422_), .C2(new_n421_), .ZN(new_n519_));
  AND3_X1   g318(.A1(new_n516_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n518_), .B1(new_n516_), .B2(new_n519_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n514_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n518_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n415_), .A2(new_n419_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT88), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n415_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n526_));
  OR2_X1    g325(.A1(new_n415_), .A2(new_n416_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n410_), .B1(KEYINPUT21), .B2(new_n404_), .ZN(new_n528_));
  AOI22_X1  g327(.A1(new_n525_), .A2(new_n526_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT20), .B1(new_n529_), .B2(new_n379_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n423_), .A2(new_n374_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n523_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n514_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n516_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n532_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n522_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n507_), .A2(KEYINPUT93), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT93), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n505_), .A2(new_n506_), .A3(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n537_), .A2(new_n493_), .A3(new_n539_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n459_), .A2(new_n495_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n541_), .A2(new_n493_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n503_), .B1(new_n491_), .B2(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n536_), .B1(new_n540_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT92), .ZN(new_n545_));
  AOI211_X1 g344(.A(new_n545_), .B(KEYINPUT33), .C1(new_n498_), .C2(new_n508_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n492_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n494_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n548_));
  OAI211_X1 g347(.A(new_n547_), .B(new_n503_), .C1(new_n548_), .C2(new_n496_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT33), .ZN(new_n550_));
  AOI21_X1  g349(.A(KEYINPUT92), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n509_), .B(new_n544_), .C1(new_n546_), .C2(new_n551_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n548_), .A2(new_n496_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n547_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n504_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(KEYINPUT99), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT99), .ZN(new_n557_));
  OAI211_X1 g356(.A(new_n557_), .B(new_n504_), .C1(new_n553_), .C2(new_n554_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n556_), .A2(new_n558_), .A3(new_n549_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n514_), .A2(KEYINPUT32), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT95), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n532_), .A2(new_n534_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(KEYINPUT96), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT96), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n561_), .A2(new_n565_), .A3(new_n562_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n529_), .A2(KEYINPUT98), .A3(new_n379_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT98), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n374_), .B1(new_n423_), .B2(new_n568_), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n515_), .A2(KEYINPUT97), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n515_), .A2(KEYINPUT97), .ZN(new_n571_));
  NOR3_X1   g370(.A1(new_n523_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n567_), .A2(new_n569_), .A3(new_n572_), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n532_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n560_), .ZN(new_n575_));
  AOI22_X1  g374(.A1(new_n564_), .A2(new_n566_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  AOI22_X1  g375(.A1(new_n552_), .A2(KEYINPUT94), .B1(new_n559_), .B2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n549_), .A2(new_n550_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(new_n545_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n549_), .A2(KEYINPUT92), .A3(new_n550_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n543_), .A2(new_n540_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n536_), .ZN(new_n583_));
  AND3_X1   g382(.A1(new_n582_), .A2(new_n583_), .A3(new_n509_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT94), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n581_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n481_), .B1(new_n577_), .B2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n532_), .A2(new_n533_), .A3(new_n573_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT100), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n532_), .A2(KEYINPUT100), .A3(new_n533_), .A4(new_n573_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n592_), .A2(new_n522_), .A3(KEYINPUT27), .ZN(new_n593_));
  OAI21_X1  g392(.A(KEYINPUT101), .B1(new_n591_), .B2(new_n593_), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n522_), .A2(KEYINPUT27), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT101), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n595_), .A2(new_n596_), .A3(new_n590_), .A4(new_n592_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n594_), .A2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(KEYINPUT102), .B(KEYINPUT27), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n536_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT103), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n536_), .A2(KEYINPUT103), .A3(new_n599_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n598_), .A2(new_n604_), .ZN(new_n605_));
  AOI22_X1  g404(.A1(new_n555_), .A2(KEYINPUT99), .B1(new_n498_), .B2(new_n508_), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n606_), .A2(new_n478_), .A3(new_n558_), .A4(new_n479_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n399_), .B1(new_n587_), .B2(new_n608_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n598_), .A2(new_n604_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n399_), .A2(new_n559_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT104), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n610_), .A2(new_n611_), .A3(new_n612_), .A4(new_n480_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n598_), .A2(new_n480_), .A3(new_n604_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n398_), .A2(new_n606_), .A3(new_n558_), .ZN(new_n615_));
  OAI21_X1  g414(.A(KEYINPUT104), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n613_), .A2(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n354_), .B1(new_n609_), .B2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n327_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n620_), .A2(new_n301_), .A3(new_n559_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT38), .ZN(new_n622_));
  OR2_X1    g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(KEYINPUT105), .B1(new_n269_), .B2(new_n354_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n326_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT105), .ZN(new_n626_));
  OAI211_X1 g425(.A(new_n626_), .B(new_n353_), .C1(new_n266_), .C2(new_n268_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n624_), .A2(new_n625_), .A3(new_n627_), .ZN(new_n628_));
  OR2_X1    g427(.A1(new_n628_), .A2(KEYINPUT106), .ZN(new_n629_));
  INV_X1    g428(.A(new_n297_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n630_), .B1(new_n609_), .B2(new_n617_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n628_), .A2(KEYINPUT106), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n629_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n559_), .ZN(new_n634_));
  OAI21_X1  g433(.A(G1gat), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n621_), .A2(new_n622_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n623_), .A2(new_n635_), .A3(new_n636_), .ZN(G1324gat));
  NAND3_X1  g436(.A1(new_n620_), .A2(new_n302_), .A3(new_n605_), .ZN(new_n638_));
  OAI21_X1  g437(.A(G8gat), .B1(new_n633_), .B2(new_n610_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n639_), .A2(KEYINPUT39), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT39), .ZN(new_n641_));
  OAI211_X1 g440(.A(new_n641_), .B(G8gat), .C1(new_n633_), .C2(new_n610_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n638_), .B1(new_n640_), .B2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT40), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  OAI211_X1 g445(.A(KEYINPUT40), .B(new_n638_), .C1(new_n640_), .C2(new_n643_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(G1325gat));
  OAI21_X1  g447(.A(G15gat), .B1(new_n633_), .B2(new_n399_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(KEYINPUT107), .B(KEYINPUT41), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n649_), .A2(new_n650_), .ZN(new_n652_));
  OR3_X1    g451(.A1(new_n619_), .A2(G15gat), .A3(new_n399_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n651_), .A2(new_n652_), .A3(new_n653_), .ZN(G1326gat));
  NAND3_X1  g453(.A1(new_n620_), .A2(new_n306_), .A3(new_n481_), .ZN(new_n655_));
  OAI21_X1  g454(.A(G22gat), .B1(new_n633_), .B2(new_n480_), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n656_), .A2(KEYINPUT42), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n656_), .A2(KEYINPUT42), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n655_), .B1(new_n658_), .B2(new_n659_), .ZN(G1327gat));
  NAND2_X1  g459(.A1(new_n630_), .A2(new_n326_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n661_), .A2(new_n269_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n618_), .A2(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(G29gat), .B1(new_n663_), .B2(new_n559_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT110), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n624_), .A2(new_n326_), .A3(new_n627_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n546_), .A2(new_n551_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n582_), .A2(new_n583_), .A3(new_n509_), .ZN(new_n668_));
  OAI21_X1  g467(.A(KEYINPUT94), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n559_), .A2(new_n576_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n669_), .A2(new_n586_), .A3(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n608_), .B1(new_n671_), .B2(new_n480_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n617_), .B1(new_n672_), .B2(new_n398_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(new_n300_), .ZN(new_n674_));
  XOR2_X1   g473(.A(KEYINPUT108), .B(KEYINPUT43), .Z(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT43), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n673_), .A2(new_n677_), .A3(new_n300_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n666_), .B1(new_n676_), .B2(new_n678_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(KEYINPUT109), .B(KEYINPUT44), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n665_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n624_), .A2(new_n326_), .A3(new_n627_), .ZN(new_n682_));
  AOI211_X1 g481(.A(KEYINPUT43), .B(new_n299_), .C1(new_n609_), .C2(new_n617_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n675_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n684_), .B1(new_n673_), .B2(new_n300_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n682_), .B1(new_n683_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n680_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n686_), .A2(KEYINPUT110), .A3(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n681_), .A2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n679_), .A2(KEYINPUT44), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n559_), .A2(G29gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n664_), .B1(new_n691_), .B2(new_n692_), .ZN(G1328gat));
  INV_X1    g492(.A(G36gat), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n663_), .A2(new_n694_), .A3(new_n605_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT45), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT111), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n610_), .B1(new_n679_), .B2(KEYINPUT44), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n299_), .B1(new_n609_), .B2(new_n617_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n678_), .B1(new_n699_), .B2(new_n684_), .ZN(new_n700_));
  AOI211_X1 g499(.A(new_n665_), .B(new_n680_), .C1(new_n700_), .C2(new_n682_), .ZN(new_n701_));
  AOI21_X1  g500(.A(KEYINPUT110), .B1(new_n686_), .B2(new_n687_), .ZN(new_n702_));
  OAI211_X1 g501(.A(new_n697_), .B(new_n698_), .C1(new_n701_), .C2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(G36gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n697_), .B1(new_n689_), .B2(new_n698_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n696_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT46), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  OAI211_X1 g507(.A(KEYINPUT46), .B(new_n696_), .C1(new_n704_), .C2(new_n705_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1329gat));
  NAND4_X1  g509(.A1(new_n689_), .A2(G43gat), .A3(new_n398_), .A4(new_n690_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n663_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n376_), .B1(new_n712_), .B2(new_n399_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g514(.A(G50gat), .B1(new_n663_), .B2(new_n481_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n481_), .A2(G50gat), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n716_), .B1(new_n691_), .B2(new_n717_), .ZN(G1331gat));
  AOI21_X1  g517(.A(new_n353_), .B1(new_n609_), .B2(new_n617_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n300_), .A2(new_n326_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n719_), .A2(new_n269_), .A3(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT112), .ZN(new_n722_));
  AOI21_X1  g521(.A(G57gat), .B1(new_n722_), .B2(new_n559_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n269_), .A2(new_n354_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n724_), .A2(new_n326_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n631_), .A2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n634_), .A2(KEYINPUT113), .ZN(new_n728_));
  MUX2_X1   g527(.A(KEYINPUT113), .B(new_n728_), .S(G57gat), .Z(new_n729_));
  AOI21_X1  g528(.A(new_n723_), .B1(new_n727_), .B2(new_n729_), .ZN(G1332gat));
  OAI21_X1  g529(.A(G64gat), .B1(new_n726_), .B2(new_n610_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT48), .ZN(new_n732_));
  INV_X1    g531(.A(new_n722_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n610_), .A2(G64gat), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT114), .Z(new_n735_));
  OAI21_X1  g534(.A(new_n732_), .B1(new_n733_), .B2(new_n735_), .ZN(G1333gat));
  OAI21_X1  g535(.A(G71gat), .B1(new_n726_), .B2(new_n399_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT49), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n399_), .A2(G71gat), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n738_), .B1(new_n733_), .B2(new_n739_), .ZN(G1334gat));
  OAI21_X1  g539(.A(G78gat), .B1(new_n726_), .B2(new_n480_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT50), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n480_), .A2(G78gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n742_), .B1(new_n733_), .B2(new_n743_), .ZN(G1335gat));
  NAND4_X1  g543(.A1(new_n719_), .A2(new_n269_), .A3(new_n326_), .A4(new_n630_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n746_), .A2(new_n212_), .A3(new_n559_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n724_), .A2(new_n625_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n700_), .A2(new_n748_), .ZN(new_n749_));
  OR2_X1    g548(.A1(new_n749_), .A2(KEYINPUT115), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(KEYINPUT115), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n634_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n747_), .B1(new_n752_), .B2(new_n212_), .ZN(G1336gat));
  AOI21_X1  g552(.A(G92gat), .B1(new_n746_), .B2(new_n605_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n750_), .A2(new_n751_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n610_), .A2(new_n211_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n754_), .B1(new_n755_), .B2(new_n756_), .ZN(G1337gat));
  NAND3_X1  g556(.A1(new_n746_), .A2(new_n398_), .A3(new_n207_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n399_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n759_));
  INV_X1    g558(.A(G99gat), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n758_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g561(.A1(new_n746_), .A2(new_n208_), .A3(new_n481_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT52), .ZN(new_n764_));
  INV_X1    g563(.A(new_n749_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(new_n481_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n764_), .B1(new_n766_), .B2(G106gat), .ZN(new_n767_));
  AOI211_X1 g566(.A(KEYINPUT52), .B(new_n208_), .C1(new_n765_), .C2(new_n481_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n763_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g569(.A1(new_n244_), .A2(KEYINPUT119), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT55), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n771_), .B1(new_n772_), .B2(new_n244_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n236_), .A2(new_n242_), .A3(new_n245_), .A4(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n236_), .A2(new_n242_), .A3(new_n245_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n771_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n246_), .A2(new_n777_), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n774_), .B(new_n776_), .C1(new_n778_), .C2(KEYINPUT118), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n778_), .A2(KEYINPUT118), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n262_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  OR2_X1    g580(.A1(new_n781_), .A2(KEYINPUT56), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n328_), .A2(new_n333_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n330_), .B1(new_n783_), .B2(KEYINPUT121), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n784_), .B1(KEYINPUT121), .B2(new_n783_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n345_), .B1(new_n347_), .B2(new_n330_), .ZN(new_n786_));
  AOI22_X1  g585(.A1(new_n785_), .A2(new_n786_), .B1(new_n342_), .B2(new_n345_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n787_), .A2(new_n260_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n781_), .A2(KEYINPUT56), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n782_), .A2(new_n788_), .A3(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT58), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n299_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n792_), .B1(new_n791_), .B2(new_n790_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT57), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n353_), .A2(new_n260_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT116), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n353_), .A2(KEYINPUT116), .A3(new_n260_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n781_), .B1(KEYINPUT120), .B2(KEYINPUT56), .ZN(new_n799_));
  NOR2_X1   g598(.A1(KEYINPUT120), .A2(KEYINPUT56), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n262_), .B(new_n800_), .C1(new_n779_), .C2(new_n780_), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n797_), .A2(new_n798_), .A3(new_n799_), .A4(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n264_), .A2(new_n787_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n794_), .B1(new_n804_), .B2(new_n297_), .ZN(new_n805_));
  AOI211_X1 g604(.A(KEYINPUT57), .B(new_n630_), .C1(new_n802_), .C2(new_n803_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n793_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(new_n326_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n269_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n720_), .A2(new_n354_), .A3(new_n809_), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n810_), .B(KEYINPUT54), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n808_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT59), .ZN(new_n813_));
  NOR3_X1   g612(.A1(new_n614_), .A2(new_n634_), .A3(new_n399_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n812_), .A2(new_n813_), .A3(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n814_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT122), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n807_), .A2(new_n817_), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n793_), .B(KEYINPUT122), .C1(new_n805_), .C2(new_n806_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n818_), .A2(new_n326_), .A3(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n816_), .B1(new_n820_), .B2(new_n811_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n815_), .B1(new_n821_), .B2(new_n813_), .ZN(new_n822_));
  OAI21_X1  g621(.A(G113gat), .B1(new_n822_), .B2(new_n354_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n821_), .ZN(new_n824_));
  OR3_X1    g623(.A1(new_n824_), .A2(G113gat), .A3(new_n354_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n823_), .A2(new_n825_), .ZN(G1340gat));
  OAI21_X1  g625(.A(G120gat), .B1(new_n822_), .B2(new_n809_), .ZN(new_n827_));
  INV_X1    g626(.A(G120gat), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n828_), .B1(new_n809_), .B2(KEYINPUT60), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n821_), .B(new_n829_), .C1(KEYINPUT60), .C2(new_n828_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n827_), .A2(new_n830_), .ZN(G1341gat));
  OAI21_X1  g630(.A(G127gat), .B1(new_n822_), .B2(new_n326_), .ZN(new_n832_));
  OR3_X1    g631(.A1(new_n824_), .A2(G127gat), .A3(new_n326_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(G1342gat));
  OAI211_X1 g633(.A(new_n300_), .B(new_n815_), .C1(new_n821_), .C2(new_n813_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(G134gat), .ZN(new_n836_));
  OR2_X1    g635(.A1(new_n297_), .A2(G134gat), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n836_), .B1(new_n824_), .B2(new_n837_), .ZN(G1343gat));
  NAND2_X1  g637(.A1(new_n820_), .A2(new_n811_), .ZN(new_n839_));
  NOR3_X1   g638(.A1(new_n634_), .A2(new_n480_), .A3(new_n398_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n839_), .A2(new_n610_), .A3(new_n840_), .ZN(new_n841_));
  OR3_X1    g640(.A1(new_n841_), .A2(G141gat), .A3(new_n354_), .ZN(new_n842_));
  OAI21_X1  g641(.A(G141gat), .B1(new_n841_), .B2(new_n354_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(G1344gat));
  OR3_X1    g643(.A1(new_n841_), .A2(G148gat), .A3(new_n809_), .ZN(new_n845_));
  OAI21_X1  g644(.A(G148gat), .B1(new_n841_), .B2(new_n809_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(G1345gat));
  XNOR2_X1  g646(.A(KEYINPUT61), .B(G155gat), .ZN(new_n848_));
  OR3_X1    g647(.A1(new_n841_), .A2(new_n326_), .A3(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n848_), .B1(new_n841_), .B2(new_n326_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(G1346gat));
  OAI21_X1  g650(.A(G162gat), .B1(new_n841_), .B2(new_n299_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n630_), .A2(new_n425_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n841_), .B2(new_n853_), .ZN(G1347gat));
  AOI21_X1  g653(.A(new_n481_), .B1(new_n808_), .B2(new_n811_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n610_), .A2(new_n615_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n855_), .A2(new_n353_), .A3(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT62), .ZN(new_n858_));
  AND4_X1   g657(.A1(KEYINPUT123), .A2(new_n857_), .A3(new_n858_), .A4(G169gat), .ZN(new_n859_));
  INV_X1    g658(.A(G169gat), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT123), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n860_), .B1(new_n861_), .B2(KEYINPUT62), .ZN(new_n862_));
  AOI22_X1  g661(.A1(new_n857_), .A2(new_n862_), .B1(KEYINPUT123), .B2(new_n858_), .ZN(new_n863_));
  XOR2_X1   g662(.A(KEYINPUT22), .B(G169gat), .Z(new_n864_));
  OAI22_X1  g663(.A1(new_n859_), .A2(new_n863_), .B1(new_n857_), .B2(new_n864_), .ZN(G1348gat));
  AND2_X1   g664(.A1(new_n855_), .A2(new_n856_), .ZN(new_n866_));
  AOI21_X1  g665(.A(G176gat), .B1(new_n866_), .B2(new_n269_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n481_), .B1(new_n820_), .B2(new_n811_), .ZN(new_n868_));
  AND3_X1   g667(.A1(new_n269_), .A2(G176gat), .A3(new_n856_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n867_), .B1(new_n868_), .B2(new_n869_), .ZN(G1349gat));
  NOR3_X1   g669(.A1(new_n326_), .A2(new_n610_), .A3(new_n615_), .ZN(new_n871_));
  AOI21_X1  g670(.A(G183gat), .B1(new_n868_), .B2(new_n871_), .ZN(new_n872_));
  NOR4_X1   g671(.A1(new_n326_), .A2(new_n356_), .A3(new_n610_), .A4(new_n615_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n872_), .B1(new_n855_), .B2(new_n873_), .ZN(G1350gat));
  NAND2_X1  g673(.A1(new_n866_), .A2(new_n300_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(G190gat), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n866_), .A2(new_n357_), .A3(new_n630_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(G1351gat));
  NOR3_X1   g677(.A1(new_n610_), .A2(new_n607_), .A3(new_n398_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n880_), .B1(new_n820_), .B2(new_n811_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n353_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g682(.A1(new_n881_), .A2(new_n269_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(KEYINPUT125), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n884_), .B(new_n886_), .ZN(G1353gat));
  INV_X1    g686(.A(KEYINPUT126), .ZN(new_n888_));
  AOI211_X1 g687(.A(new_n326_), .B(new_n880_), .C1(new_n820_), .C2(new_n811_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n888_), .B1(new_n889_), .B2(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n881_), .A2(new_n625_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n893_), .A2(KEYINPUT126), .A3(new_n890_), .ZN(new_n894_));
  XOR2_X1   g693(.A(KEYINPUT63), .B(G211gat), .Z(new_n895_));
  AOI22_X1  g694(.A1(new_n892_), .A2(new_n894_), .B1(new_n889_), .B2(new_n895_), .ZN(G1354gat));
  INV_X1    g695(.A(KEYINPUT127), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n406_), .B1(new_n881_), .B2(new_n300_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n297_), .A2(G218gat), .ZN(new_n899_));
  AND3_X1   g698(.A1(new_n839_), .A2(new_n879_), .A3(new_n899_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n897_), .B1(new_n898_), .B2(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n881_), .A2(new_n899_), .ZN(new_n902_));
  AOI211_X1 g701(.A(new_n299_), .B(new_n880_), .C1(new_n820_), .C2(new_n811_), .ZN(new_n903_));
  OAI211_X1 g702(.A(new_n902_), .B(KEYINPUT127), .C1(new_n903_), .C2(new_n406_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n901_), .A2(new_n904_), .ZN(G1355gat));
endmodule


