//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 1 0 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 1 0 0 0 0 0 0 0 1 0 1 0 0 1 0 0 1 0 0 0 0 1 1 0 0 0 1 0 1 1 1 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n768_, new_n769_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n885_, new_n886_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n919_, new_n920_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_, new_n943_;
  AND2_X1   g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202_));
  NOR2_X1   g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  OR2_X1    g003(.A1(G141gat), .A2(G148gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT93), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT3), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT2), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210_));
  AOI22_X1  g009(.A1(new_n205_), .A2(new_n208_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n211_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(KEYINPUT93), .A2(KEYINPUT3), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n213_), .B1(new_n205_), .B2(new_n208_), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n204_), .B1(new_n212_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT94), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n215_), .B(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n202_), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n203_), .B1(new_n218_), .B2(KEYINPUT1), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n219_), .B1(KEYINPUT1), .B2(new_n218_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n220_), .A2(new_n205_), .A3(new_n210_), .ZN(new_n221_));
  AND2_X1   g020(.A1(new_n217_), .A2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G127gat), .B(G134gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G113gat), .B(G120gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n223_), .B(new_n224_), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n223_), .A2(new_n224_), .ZN(new_n226_));
  MUX2_X1   g025(.A(new_n225_), .B(new_n226_), .S(KEYINPUT91), .Z(new_n227_));
  NOR2_X1   g026(.A1(new_n222_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT4), .ZN(new_n229_));
  AOI21_X1  g028(.A(KEYINPUT104), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  XOR2_X1   g029(.A(new_n225_), .B(KEYINPUT103), .Z(new_n231_));
  NAND2_X1  g030(.A1(new_n222_), .A2(new_n231_), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n232_), .B(KEYINPUT4), .C1(new_n222_), .C2(new_n227_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n230_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n228_), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n235_), .A2(KEYINPUT104), .A3(KEYINPUT4), .A4(new_n232_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G225gat), .A2(G233gat), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n235_), .A2(new_n232_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n241_), .A2(new_n239_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G1gat), .B(G29gat), .ZN(new_n244_));
  INV_X1    g043(.A(G85gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT0), .B(G57gat), .ZN(new_n247_));
  XOR2_X1   g046(.A(new_n246_), .B(new_n247_), .Z(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n240_), .A2(new_n243_), .A3(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n238_), .B1(new_n234_), .B2(new_n236_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n248_), .B1(new_n251_), .B2(new_n242_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  XOR2_X1   g053(.A(KEYINPUT97), .B(G197gat), .Z(new_n255_));
  NOR2_X1   g054(.A1(new_n255_), .A2(G204gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT98), .B(G204gat), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n257_), .A2(G197gat), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT21), .B1(new_n256_), .B2(new_n258_), .ZN(new_n259_));
  AOI22_X1  g058(.A1(new_n255_), .A2(G204gat), .B1(new_n257_), .B2(G197gat), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT21), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G211gat), .B(G218gat), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n259_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  OR3_X1    g063(.A1(new_n260_), .A2(new_n261_), .A3(new_n263_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(G169gat), .ZN(new_n268_));
  INV_X1    g067(.A(G176gat), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT22), .B(G169gat), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n270_), .B1(new_n271_), .B2(new_n269_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT23), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n273_), .A2(G183gat), .A3(G190gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT88), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n273_), .B1(G183gat), .B2(G190gat), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(G183gat), .A2(G190gat), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n272_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT86), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n280_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n281_));
  OAI21_X1  g080(.A(KEYINPUT86), .B1(G169gat), .B2(G176gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT24), .ZN(new_n284_));
  OR3_X1    g083(.A1(new_n283_), .A2(new_n284_), .A3(new_n270_), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n285_), .A2(KEYINPUT87), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(KEYINPUT87), .ZN(new_n287_));
  INV_X1    g086(.A(new_n276_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(new_n274_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n283_), .A2(new_n284_), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n286_), .A2(new_n287_), .A3(new_n289_), .A4(new_n290_), .ZN(new_n291_));
  AND2_X1   g090(.A1(KEYINPUT83), .A2(KEYINPUT25), .ZN(new_n292_));
  NOR2_X1   g091(.A1(KEYINPUT83), .A2(KEYINPUT25), .ZN(new_n293_));
  OAI21_X1  g092(.A(G183gat), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT84), .ZN(new_n295_));
  OR2_X1    g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(G190gat), .ZN(new_n297_));
  OR2_X1    g096(.A1(new_n297_), .A2(KEYINPUT26), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT25), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n298_), .B1(new_n299_), .B2(G183gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n297_), .A2(KEYINPUT26), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n300_), .B1(KEYINPUT85), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n294_), .A2(new_n295_), .ZN(new_n303_));
  OR2_X1    g102(.A1(new_n301_), .A2(KEYINPUT85), .ZN(new_n304_));
  AND4_X1   g103(.A1(new_n296_), .A2(new_n302_), .A3(new_n303_), .A4(new_n304_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n279_), .B1(new_n291_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT89), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT89), .ZN(new_n308_));
  OAI211_X1 g107(.A(new_n308_), .B(new_n279_), .C1(new_n291_), .C2(new_n305_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n267_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G226gat), .A2(G233gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT19), .ZN(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT25), .B(G183gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n313_), .A2(new_n301_), .A3(new_n298_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n285_), .A2(new_n290_), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n272_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n278_), .B1(new_n288_), .B2(new_n274_), .ZN(new_n317_));
  OAI22_X1  g116(.A1(new_n315_), .A2(new_n277_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT20), .B1(new_n266_), .B2(new_n318_), .ZN(new_n319_));
  NOR3_X1   g118(.A1(new_n310_), .A2(new_n312_), .A3(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n312_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n307_), .A2(new_n267_), .A3(new_n309_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT20), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n323_), .B1(new_n266_), .B2(new_n318_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n321_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G8gat), .B(G36gat), .ZN(new_n326_));
  INV_X1    g125(.A(G92gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT18), .B(G64gat), .ZN(new_n329_));
  XOR2_X1   g128(.A(new_n328_), .B(new_n329_), .Z(new_n330_));
  NOR3_X1   g129(.A1(new_n320_), .A2(new_n325_), .A3(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n330_), .B1(new_n320_), .B2(new_n325_), .ZN(new_n333_));
  AOI21_X1  g132(.A(KEYINPUT27), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n310_), .A2(new_n319_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n335_), .A2(new_n321_), .ZN(new_n336_));
  AND3_X1   g135(.A1(new_n322_), .A2(new_n321_), .A3(new_n324_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n330_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT27), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n331_), .A2(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n334_), .B1(new_n338_), .B2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G22gat), .B(G50gat), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT95), .B(KEYINPUT28), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n217_), .A2(new_n221_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n344_), .B1(new_n345_), .B2(KEYINPUT29), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NOR3_X1   g146(.A1(new_n345_), .A2(KEYINPUT29), .A3(new_n344_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n343_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n348_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n350_), .A2(new_n342_), .A3(new_n346_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n349_), .A2(new_n351_), .ZN(new_n352_));
  XOR2_X1   g151(.A(G78gat), .B(G106gat), .Z(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT100), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT99), .B(KEYINPUT29), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n267_), .B1(new_n345_), .B2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(G228gat), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n357_), .A2(KEYINPUT96), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n357_), .A2(KEYINPUT96), .ZN(new_n359_));
  OAI21_X1  g158(.A(G233gat), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  OR2_X1    g159(.A1(new_n356_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n345_), .A2(KEYINPUT29), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n362_), .A2(new_n360_), .A3(new_n266_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n361_), .A2(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n352_), .A2(new_n354_), .A3(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n349_), .A2(new_n351_), .A3(KEYINPUT102), .ZN(new_n366_));
  XOR2_X1   g165(.A(new_n354_), .B(KEYINPUT101), .Z(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n368_), .B1(new_n361_), .B2(new_n363_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n361_), .A2(new_n368_), .A3(new_n363_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n366_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n366_), .A2(new_n371_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n365_), .B1(new_n372_), .B2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n307_), .A2(new_n309_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G71gat), .B(G99gat), .ZN(new_n377_));
  INV_X1    g176(.A(G43gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  AND2_X1   g178(.A1(G227gat), .A2(G233gat), .ZN(new_n380_));
  XOR2_X1   g179(.A(new_n379_), .B(new_n380_), .Z(new_n381_));
  NAND2_X1  g180(.A1(new_n376_), .A2(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT30), .B(G15gat), .ZN(new_n383_));
  XOR2_X1   g182(.A(new_n383_), .B(KEYINPUT90), .Z(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n381_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n307_), .A2(new_n309_), .A3(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n382_), .A2(new_n385_), .A3(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  XOR2_X1   g188(.A(new_n227_), .B(KEYINPUT31), .Z(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT92), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n385_), .B1(new_n382_), .B2(new_n387_), .ZN(new_n392_));
  OR3_X1    g191(.A1(new_n389_), .A2(new_n391_), .A3(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT92), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n390_), .A2(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n395_), .B1(new_n389_), .B2(new_n392_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n393_), .A2(new_n396_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n375_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n371_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n399_), .A2(new_n369_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n373_), .B1(new_n400_), .B2(new_n366_), .ZN(new_n401_));
  AOI22_X1  g200(.A1(new_n401_), .A2(new_n365_), .B1(new_n393_), .B2(new_n396_), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n254_), .B(new_n341_), .C1(new_n398_), .C2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n237_), .A2(new_n238_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n248_), .B1(new_n241_), .B2(new_n238_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n404_), .A2(KEYINPUT105), .A3(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT105), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n239_), .B1(new_n234_), .B2(new_n236_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n408_), .B1(new_n409_), .B2(new_n405_), .ZN(new_n410_));
  AND4_X1   g209(.A1(new_n332_), .A2(new_n407_), .A3(new_n333_), .A4(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n242_), .B1(new_n237_), .B2(new_n239_), .ZN(new_n412_));
  AOI21_X1  g211(.A(KEYINPUT33), .B1(new_n412_), .B2(new_n249_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT33), .ZN(new_n414_));
  NOR4_X1   g213(.A1(new_n251_), .A2(new_n414_), .A3(new_n242_), .A4(new_n248_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n330_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT32), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NOR3_X1   g218(.A1(new_n320_), .A2(new_n325_), .A3(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT106), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n419_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n420_), .A2(new_n421_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  AOI22_X1  g225(.A1(new_n411_), .A2(new_n416_), .B1(new_n253_), .B2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n397_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(new_n375_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n403_), .B1(new_n427_), .B2(new_n429_), .ZN(new_n430_));
  AND3_X1   g229(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n431_));
  AOI21_X1  g230(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n432_));
  NOR3_X1   g231(.A1(new_n431_), .A2(new_n432_), .A3(KEYINPUT64), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT64), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G99gat), .A2(G106gat), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT6), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n434_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n433_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n245_), .A2(new_n327_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G85gat), .A2(G92gat), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n441_), .A2(KEYINPUT9), .A3(new_n442_), .ZN(new_n443_));
  OR2_X1    g242(.A1(new_n442_), .A2(KEYINPUT9), .ZN(new_n444_));
  XNOR2_X1  g243(.A(KEYINPUT10), .B(G99gat), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n443_), .B(new_n444_), .C1(G106gat), .C2(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(KEYINPUT65), .B1(new_n440_), .B2(new_n446_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n442_), .A2(KEYINPUT9), .ZN(new_n448_));
  XOR2_X1   g247(.A(KEYINPUT10), .B(G99gat), .Z(new_n449_));
  INV_X1    g248(.A(G106gat), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n448_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(KEYINPUT64), .B1(new_n431_), .B2(new_n432_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n437_), .A2(new_n434_), .A3(new_n438_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT65), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n451_), .A2(new_n454_), .A3(new_n455_), .A4(new_n443_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT8), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT66), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT7), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n458_), .B(new_n459_), .C1(G99gat), .C2(G106gat), .ZN(new_n460_));
  INV_X1    g259(.A(G99gat), .ZN(new_n461_));
  OAI211_X1 g260(.A(new_n461_), .B(new_n450_), .C1(KEYINPUT66), .C2(KEYINPUT7), .ZN(new_n462_));
  NAND2_X1  g261(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n460_), .B1(new_n462_), .B2(new_n464_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n431_), .A2(new_n432_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  XOR2_X1   g266(.A(G85gat), .B(G92gat), .Z(new_n468_));
  AOI21_X1  g267(.A(new_n457_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n457_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n470_), .B1(new_n454_), .B2(new_n465_), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n447_), .B(new_n456_), .C1(new_n469_), .C2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT11), .ZN(new_n473_));
  INV_X1    g272(.A(G57gat), .ZN(new_n474_));
  INV_X1    g273(.A(G64gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G57gat), .A2(G64gat), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n473_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n476_), .A2(new_n473_), .A3(new_n477_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT67), .ZN(new_n481_));
  AND2_X1   g280(.A1(G71gat), .A2(G78gat), .ZN(new_n482_));
  NOR2_X1   g281(.A1(G71gat), .A2(G78gat), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n480_), .A2(new_n481_), .A3(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n481_), .B1(new_n480_), .B2(new_n484_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n479_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n480_), .A2(new_n484_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(KEYINPUT67), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n490_), .A2(new_n485_), .A3(new_n478_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n488_), .A2(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n472_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G230gat), .A2(G233gat), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n493_), .A2(new_n495_), .ZN(new_n496_));
  AND3_X1   g295(.A1(new_n488_), .A2(new_n491_), .A3(KEYINPUT69), .ZN(new_n497_));
  AOI21_X1  g296(.A(KEYINPUT69), .B1(new_n488_), .B2(new_n491_), .ZN(new_n498_));
  OAI211_X1 g297(.A(KEYINPUT12), .B(new_n472_), .C1(new_n497_), .C2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n472_), .A2(new_n492_), .ZN(new_n500_));
  XOR2_X1   g299(.A(KEYINPUT70), .B(KEYINPUT12), .Z(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n496_), .A2(new_n499_), .A3(new_n502_), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n488_), .A2(new_n491_), .ZN(new_n504_));
  AND2_X1   g303(.A1(new_n447_), .A2(new_n456_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT68), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n441_), .A2(new_n442_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n507_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n458_), .A2(new_n459_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(G99gat), .A2(G106gat), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n509_), .A2(new_n510_), .A3(new_n463_), .ZN(new_n511_));
  AOI22_X1  g310(.A1(new_n452_), .A2(new_n453_), .B1(new_n511_), .B2(new_n460_), .ZN(new_n512_));
  OAI22_X1  g311(.A1(new_n508_), .A2(new_n457_), .B1(new_n512_), .B2(new_n470_), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n504_), .A2(new_n505_), .A3(new_n506_), .A4(new_n513_), .ZN(new_n514_));
  OAI21_X1  g313(.A(KEYINPUT68), .B1(new_n472_), .B2(new_n492_), .ZN(new_n515_));
  AOI22_X1  g314(.A1(new_n514_), .A2(new_n515_), .B1(new_n472_), .B2(new_n492_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n503_), .B1(new_n516_), .B2(new_n494_), .ZN(new_n517_));
  XOR2_X1   g316(.A(G176gat), .B(G204gat), .Z(new_n518_));
  XNOR2_X1  g317(.A(G120gat), .B(G148gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n521_));
  XOR2_X1   g320(.A(new_n520_), .B(new_n521_), .Z(new_n522_));
  NAND2_X1  g321(.A1(new_n517_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n522_), .ZN(new_n524_));
  OAI211_X1 g323(.A(new_n503_), .B(new_n524_), .C1(new_n516_), .C2(new_n494_), .ZN(new_n525_));
  AND3_X1   g324(.A1(new_n523_), .A2(KEYINPUT13), .A3(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(KEYINPUT13), .B1(new_n523_), .B2(new_n525_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G229gat), .A2(G233gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G29gat), .B(G36gat), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G43gat), .B(G50gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n533_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(new_n531_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G1gat), .B(G8gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT77), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G15gat), .B(G22gat), .ZN(new_n541_));
  INV_X1    g340(.A(G1gat), .ZN(new_n542_));
  INV_X1    g341(.A(G8gat), .ZN(new_n543_));
  OAI21_X1  g342(.A(KEYINPUT14), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n541_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n540_), .A2(new_n545_), .ZN(new_n546_));
  OR2_X1    g345(.A1(new_n539_), .A2(KEYINPUT77), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n539_), .A2(KEYINPUT77), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n547_), .A2(new_n544_), .A3(new_n541_), .A4(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n538_), .A2(new_n546_), .A3(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(KEYINPUT73), .B(KEYINPUT15), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n537_), .A2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n534_), .A2(new_n536_), .A3(new_n552_), .ZN(new_n555_));
  AOI22_X1  g354(.A1(new_n554_), .A2(new_n555_), .B1(new_n546_), .B2(new_n549_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n530_), .B1(new_n551_), .B2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n546_), .A2(new_n549_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(new_n537_), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n559_), .A2(G229gat), .A3(G233gat), .A4(new_n550_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n557_), .A2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G113gat), .B(G141gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G169gat), .B(G197gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n561_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT81), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT82), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n566_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n564_), .B1(new_n557_), .B2(new_n560_), .ZN(new_n570_));
  OAI21_X1  g369(.A(KEYINPUT82), .B1(new_n570_), .B2(KEYINPUT81), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n561_), .A2(new_n565_), .ZN(new_n572_));
  AND3_X1   g371(.A1(new_n569_), .A2(new_n571_), .A3(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n572_), .B1(new_n569_), .B2(new_n571_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n529_), .A2(new_n576_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n430_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G231gat), .A2(G233gat), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n579_), .B(KEYINPUT78), .Z(new_n580_));
  XNOR2_X1  g379(.A(new_n558_), .B(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT69), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n492_), .A2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n488_), .A2(new_n491_), .A3(KEYINPUT69), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n581_), .B(new_n585_), .ZN(new_n586_));
  XOR2_X1   g385(.A(KEYINPUT80), .B(KEYINPUT17), .Z(new_n587_));
  XOR2_X1   g386(.A(G183gat), .B(G211gat), .Z(new_n588_));
  XNOR2_X1  g387(.A(G127gat), .B(G155gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  NOR3_X1   g391(.A1(new_n586_), .A2(new_n587_), .A3(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(KEYINPUT17), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n594_), .B1(new_n504_), .B2(new_n581_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n595_), .B1(new_n504_), .B2(new_n581_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n593_), .A2(new_n596_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n513_), .A2(new_n538_), .A3(new_n447_), .A4(new_n456_), .ZN(new_n598_));
  XOR2_X1   g397(.A(KEYINPUT72), .B(KEYINPUT34), .Z(new_n599_));
  NAND2_X1  g398(.A1(G232gat), .A2(G233gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT35), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n598_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT74), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n554_), .A2(new_n555_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n472_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n605_), .B1(new_n472_), .B2(new_n606_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n604_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n601_), .A2(new_n602_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G190gat), .B(G218gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G134gat), .B(G162gat), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n612_), .B(new_n613_), .Z(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n615_), .A2(KEYINPUT36), .ZN(new_n616_));
  INV_X1    g415(.A(new_n610_), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n604_), .B(new_n617_), .C1(new_n607_), .C2(new_n608_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n611_), .A2(new_n616_), .A3(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT75), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n611_), .A2(KEYINPUT75), .A3(new_n616_), .A4(new_n618_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n611_), .A2(new_n618_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n614_), .B(KEYINPUT36), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n623_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT37), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n627_), .A2(KEYINPUT76), .A3(new_n628_), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n628_), .A2(KEYINPUT76), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(KEYINPUT76), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n623_), .A2(new_n626_), .A3(new_n630_), .A4(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n629_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n578_), .A2(new_n597_), .A3(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n253_), .B(KEYINPUT107), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n635_), .A2(new_n542_), .A3(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT38), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT108), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n627_), .A2(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n623_), .A2(KEYINPUT108), .A3(new_n626_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n597_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n578_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  OAI21_X1  g448(.A(G1gat), .B1(new_n649_), .B2(new_n254_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n638_), .A2(new_n639_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n640_), .A2(new_n650_), .A3(new_n651_), .ZN(G1324gat));
  INV_X1    g451(.A(new_n341_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n635_), .A2(new_n543_), .A3(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT39), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n648_), .A2(new_n653_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n655_), .B1(new_n656_), .B2(G8gat), .ZN(new_n657_));
  AOI211_X1 g456(.A(KEYINPUT39), .B(new_n543_), .C1(new_n648_), .C2(new_n653_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n654_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT40), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  OAI211_X1 g460(.A(KEYINPUT40), .B(new_n654_), .C1(new_n657_), .C2(new_n658_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1325gat));
  OAI21_X1  g462(.A(G15gat), .B1(new_n649_), .B2(new_n428_), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n664_), .A2(KEYINPUT41), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(KEYINPUT41), .ZN(new_n666_));
  INV_X1    g465(.A(G15gat), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n635_), .A2(new_n667_), .A3(new_n397_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n665_), .A2(new_n666_), .A3(new_n668_), .ZN(G1326gat));
  INV_X1    g468(.A(G22gat), .ZN(new_n670_));
  INV_X1    g469(.A(new_n375_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n670_), .B1(new_n648_), .B2(new_n671_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(KEYINPUT109), .B(KEYINPUT42), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n672_), .B(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n635_), .A2(new_n670_), .A3(new_n671_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(G1327gat));
  NOR2_X1   g475(.A1(new_n644_), .A2(new_n597_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n578_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(G29gat), .B1(new_n679_), .B2(new_n253_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n577_), .A2(new_n646_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n424_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n425_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n682_), .A2(new_n253_), .A3(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n415_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n250_), .A2(new_n414_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n407_), .A2(new_n410_), .A3(new_n332_), .A4(new_n333_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n684_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n429_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n340_), .A2(new_n338_), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n691_), .A2(new_n253_), .A3(new_n334_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n375_), .A2(new_n397_), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n401_), .A2(new_n365_), .A3(new_n393_), .A4(new_n396_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  AOI22_X1  g494(.A1(new_n689_), .A2(new_n690_), .B1(new_n692_), .B2(new_n695_), .ZN(new_n696_));
  OAI21_X1  g495(.A(KEYINPUT43), .B1(new_n696_), .B2(new_n634_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT43), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n430_), .A2(new_n698_), .A3(new_n633_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n681_), .B1(new_n697_), .B2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  AND3_X1   g502(.A1(new_n703_), .A2(G29gat), .A3(new_n637_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n681_), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n696_), .A2(KEYINPUT43), .A3(new_n634_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n698_), .B1(new_n430_), .B2(new_n633_), .ZN(new_n707_));
  OAI211_X1 g506(.A(KEYINPUT44), .B(new_n705_), .C1(new_n706_), .C2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(KEYINPUT110), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT110), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n700_), .A2(new_n710_), .A3(KEYINPUT44), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n709_), .A2(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n680_), .B1(new_n704_), .B2(new_n712_), .ZN(G1328gat));
  INV_X1    g512(.A(KEYINPUT46), .ZN(new_n714_));
  INV_X1    g513(.A(G36gat), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n653_), .B1(new_n700_), .B2(KEYINPUT44), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n715_), .B1(new_n712_), .B2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n653_), .A2(new_n715_), .ZN(new_n719_));
  OR3_X1    g518(.A1(new_n678_), .A2(KEYINPUT45), .A3(new_n719_), .ZN(new_n720_));
  OAI21_X1  g519(.A(KEYINPUT45), .B1(new_n678_), .B2(new_n719_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n714_), .B1(new_n718_), .B2(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n716_), .B1(new_n709_), .B2(new_n711_), .ZN(new_n725_));
  OAI211_X1 g524(.A(KEYINPUT46), .B(new_n722_), .C1(new_n725_), .C2(new_n715_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(G1329gat));
  OAI211_X1 g526(.A(G43gat), .B(new_n397_), .C1(new_n700_), .C2(KEYINPUT44), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n728_), .B1(new_n709_), .B2(new_n711_), .ZN(new_n729_));
  AOI21_X1  g528(.A(G43gat), .B1(new_n679_), .B2(new_n397_), .ZN(new_n730_));
  OAI21_X1  g529(.A(KEYINPUT47), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT47), .ZN(new_n732_));
  INV_X1    g531(.A(new_n730_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n712_), .ZN(new_n734_));
  OAI211_X1 g533(.A(new_n732_), .B(new_n733_), .C1(new_n734_), .C2(new_n728_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n731_), .A2(new_n735_), .ZN(G1330gat));
  AOI21_X1  g535(.A(G50gat), .B1(new_n679_), .B2(new_n671_), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n703_), .A2(G50gat), .A3(new_n671_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n737_), .B1(new_n738_), .B2(new_n712_), .ZN(G1331gat));
  NOR2_X1   g538(.A1(new_n528_), .A2(new_n575_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n430_), .A2(new_n740_), .ZN(new_n741_));
  NOR3_X1   g540(.A1(new_n741_), .A2(new_n646_), .A3(new_n633_), .ZN(new_n742_));
  AOI21_X1  g541(.A(G57gat), .B1(new_n742_), .B2(new_n637_), .ZN(new_n743_));
  NOR3_X1   g542(.A1(new_n741_), .A2(new_n646_), .A3(new_n645_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n254_), .A2(new_n474_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n743_), .B1(new_n744_), .B2(new_n745_), .ZN(G1332gat));
  AOI21_X1  g545(.A(new_n475_), .B1(new_n744_), .B2(new_n653_), .ZN(new_n747_));
  XOR2_X1   g546(.A(new_n747_), .B(KEYINPUT48), .Z(new_n748_));
  NAND3_X1  g547(.A1(new_n742_), .A2(new_n475_), .A3(new_n653_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(G1333gat));
  INV_X1    g549(.A(G71gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(new_n744_), .B2(new_n397_), .ZN(new_n752_));
  XOR2_X1   g551(.A(new_n752_), .B(KEYINPUT49), .Z(new_n753_));
  NAND3_X1  g552(.A1(new_n742_), .A2(new_n751_), .A3(new_n397_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(G1334gat));
  INV_X1    g554(.A(G78gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n756_), .B1(new_n744_), .B2(new_n671_), .ZN(new_n757_));
  XOR2_X1   g556(.A(new_n757_), .B(KEYINPUT50), .Z(new_n758_));
  NAND3_X1  g557(.A1(new_n742_), .A2(new_n756_), .A3(new_n671_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(G1335gat));
  NOR3_X1   g559(.A1(new_n741_), .A2(new_n597_), .A3(new_n644_), .ZN(new_n761_));
  AOI21_X1  g560(.A(G85gat), .B1(new_n761_), .B2(new_n637_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n740_), .A2(new_n646_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n763_), .B1(new_n697_), .B2(new_n699_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT111), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n254_), .A2(new_n245_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n762_), .B1(new_n765_), .B2(new_n766_), .ZN(G1336gat));
  AOI21_X1  g566(.A(G92gat), .B1(new_n761_), .B2(new_n653_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n341_), .A2(new_n327_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n768_), .B1(new_n765_), .B2(new_n769_), .ZN(G1337gat));
  AOI21_X1  g569(.A(new_n461_), .B1(new_n764_), .B2(new_n397_), .ZN(new_n771_));
  AND3_X1   g570(.A1(new_n761_), .A2(new_n449_), .A3(new_n397_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT112), .ZN(new_n773_));
  OAI22_X1  g572(.A1(new_n771_), .A2(new_n772_), .B1(new_n773_), .B2(KEYINPUT51), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(KEYINPUT51), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n774_), .B(new_n775_), .ZN(G1338gat));
  NAND3_X1  g575(.A1(new_n761_), .A2(new_n450_), .A3(new_n671_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n764_), .A2(new_n671_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n778_), .B1(new_n779_), .B2(G106gat), .ZN(new_n780_));
  AOI211_X1 g579(.A(KEYINPUT52), .B(new_n450_), .C1(new_n764_), .C2(new_n671_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n777_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT53), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT53), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n784_), .B(new_n777_), .C1(new_n780_), .C2(new_n781_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n785_), .ZN(G1339gat));
  NOR2_X1   g585(.A1(new_n636_), .A2(new_n653_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n402_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n574_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n569_), .A2(new_n571_), .A3(new_n572_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n789_), .A2(new_n790_), .A3(new_n525_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT113), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n503_), .A2(new_n792_), .A3(new_n793_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n496_), .A2(KEYINPUT55), .A3(new_n499_), .A4(new_n502_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT114), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n472_), .A2(KEYINPUT12), .ZN(new_n797_));
  AOI22_X1  g596(.A1(new_n797_), .A2(new_n585_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n798_), .A2(new_n799_), .A3(KEYINPUT55), .A4(new_n496_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n794_), .A2(new_n796_), .A3(new_n800_), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n514_), .A2(new_n515_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n499_), .A2(new_n502_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n495_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(KEYINPUT55), .B1(new_n798_), .B2(new_n496_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n804_), .B1(new_n805_), .B2(new_n792_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n522_), .B1(new_n801_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT56), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  OAI211_X1 g608(.A(KEYINPUT56), .B(new_n522_), .C1(new_n801_), .C2(new_n806_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n791_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n523_), .A2(new_n525_), .ZN(new_n812_));
  OR3_X1    g611(.A1(new_n551_), .A2(new_n556_), .A3(new_n530_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n559_), .A2(new_n550_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n565_), .B1(new_n814_), .B2(new_n530_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n570_), .B1(new_n813_), .B2(new_n815_), .ZN(new_n816_));
  AND2_X1   g615(.A1(new_n812_), .A2(new_n816_), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n644_), .B(KEYINPUT57), .C1(new_n811_), .C2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT115), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT57), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n809_), .A2(new_n810_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n791_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n817_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n820_), .B1(new_n823_), .B2(new_n645_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n819_), .A2(new_n824_), .ZN(new_n825_));
  OAI211_X1 g624(.A(KEYINPUT115), .B(new_n820_), .C1(new_n823_), .C2(new_n645_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n525_), .A2(new_n816_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(KEYINPUT116), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n821_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT58), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n821_), .A2(KEYINPUT58), .A3(new_n828_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n831_), .A2(new_n633_), .A3(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n825_), .A2(new_n826_), .A3(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n646_), .ZN(new_n835_));
  NOR3_X1   g634(.A1(new_n575_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n836_), .A2(new_n629_), .A3(new_n597_), .A4(new_n632_), .ZN(new_n837_));
  XOR2_X1   g636(.A(new_n837_), .B(KEYINPUT54), .Z(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n788_), .B1(new_n835_), .B2(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(G113gat), .B1(new_n840_), .B2(new_n575_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT59), .ZN(new_n842_));
  OAI21_X1  g641(.A(KEYINPUT117), .B1(new_n840_), .B2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT117), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n838_), .B1(new_n834_), .B2(new_n646_), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n844_), .B(KEYINPUT59), .C1(new_n845_), .C2(new_n788_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n833_), .A2(new_n824_), .A3(new_n818_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n646_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT118), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n847_), .A2(KEYINPUT118), .A3(new_n646_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n850_), .A2(new_n839_), .A3(new_n851_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n788_), .A2(KEYINPUT59), .ZN(new_n853_));
  AOI22_X1  g652(.A1(new_n843_), .A2(new_n846_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  AND2_X1   g653(.A1(new_n575_), .A2(G113gat), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n841_), .B1(new_n854_), .B2(new_n855_), .ZN(G1340gat));
  INV_X1    g655(.A(G120gat), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n857_), .B1(new_n528_), .B2(KEYINPUT60), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n840_), .B(new_n858_), .C1(KEYINPUT60), .C2(new_n857_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n852_), .A2(new_n853_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n846_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n788_), .ZN(new_n862_));
  AOI22_X1  g661(.A1(new_n829_), .A2(new_n830_), .B1(new_n632_), .B2(new_n629_), .ZN(new_n863_));
  AOI22_X1  g662(.A1(new_n819_), .A2(new_n824_), .B1(new_n832_), .B2(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n597_), .B1(new_n864_), .B2(new_n826_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n862_), .B1(new_n865_), .B2(new_n838_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n844_), .B1(new_n866_), .B2(KEYINPUT59), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n529_), .B(new_n860_), .C1(new_n861_), .C2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT119), .ZN(new_n869_));
  OAI21_X1  g668(.A(G120gat), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(KEYINPUT119), .B1(new_n854_), .B2(new_n529_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n859_), .B1(new_n870_), .B2(new_n871_), .ZN(G1341gat));
  AOI21_X1  g671(.A(G127gat), .B1(new_n840_), .B2(new_n597_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(KEYINPUT120), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n597_), .A2(G127gat), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n874_), .B1(new_n854_), .B2(new_n875_), .ZN(G1342gat));
  AOI21_X1  g675(.A(G134gat), .B1(new_n840_), .B2(new_n645_), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n633_), .A2(G134gat), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n877_), .B1(new_n854_), .B2(new_n878_), .ZN(G1343gat));
  INV_X1    g678(.A(new_n845_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n880_), .A2(new_n398_), .A3(new_n787_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n881_), .A2(new_n576_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(KEYINPUT121), .B(G141gat), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n882_), .B(new_n883_), .ZN(G1344gat));
  INV_X1    g683(.A(new_n881_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n529_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(G148gat), .ZN(G1345gat));
  OR3_X1    g686(.A1(new_n881_), .A2(KEYINPUT122), .A3(new_n646_), .ZN(new_n888_));
  OAI21_X1  g687(.A(KEYINPUT122), .B1(new_n881_), .B2(new_n646_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(KEYINPUT61), .B(G155gat), .ZN(new_n890_));
  AND3_X1   g689(.A1(new_n888_), .A2(new_n889_), .A3(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n890_), .B1(new_n888_), .B2(new_n889_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n891_), .A2(new_n892_), .ZN(G1346gat));
  INV_X1    g692(.A(G162gat), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n881_), .A2(new_n894_), .A3(new_n634_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n885_), .A2(new_n645_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n895_), .B1(new_n896_), .B2(new_n894_), .ZN(G1347gat));
  NAND3_X1  g696(.A1(new_n636_), .A2(new_n397_), .A3(new_n653_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(new_n671_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n852_), .A2(new_n899_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n901_), .A2(new_n575_), .A3(new_n271_), .ZN(new_n902_));
  OAI21_X1  g701(.A(G169gat), .B1(new_n900_), .B2(new_n576_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT124), .ZN(new_n904_));
  XOR2_X1   g703(.A(KEYINPUT123), .B(KEYINPUT62), .Z(new_n905_));
  NAND3_X1  g704(.A1(new_n903_), .A2(new_n904_), .A3(new_n905_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n906_), .B1(new_n903_), .B2(new_n905_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n904_), .B1(new_n903_), .B2(new_n905_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n902_), .B1(new_n907_), .B2(new_n908_), .ZN(G1348gat));
  AOI21_X1  g708(.A(G176gat), .B1(new_n901_), .B2(new_n529_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n845_), .A2(new_n671_), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n898_), .A2(new_n269_), .A3(new_n528_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n910_), .B1(new_n911_), .B2(new_n912_), .ZN(G1349gat));
  NOR3_X1   g712(.A1(new_n900_), .A2(new_n313_), .A3(new_n646_), .ZN(new_n914_));
  INV_X1    g713(.A(G183gat), .ZN(new_n915_));
  INV_X1    g714(.A(new_n898_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n911_), .A2(new_n597_), .A3(new_n916_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n914_), .B1(new_n915_), .B2(new_n917_), .ZN(G1350gat));
  OAI21_X1  g717(.A(G190gat), .B1(new_n900_), .B2(new_n634_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n645_), .A2(new_n301_), .A3(new_n298_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n919_), .B1(new_n900_), .B2(new_n920_), .ZN(G1351gat));
  NOR2_X1   g720(.A1(new_n341_), .A2(new_n253_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n880_), .A2(new_n398_), .A3(new_n922_), .ZN(new_n923_));
  INV_X1    g722(.A(new_n923_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(new_n575_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g725(.A1(new_n923_), .A2(new_n528_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT125), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n927_), .B1(new_n928_), .B2(G204gat), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n257_), .B1(KEYINPUT125), .B2(G204gat), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n929_), .B1(new_n927_), .B2(new_n930_), .ZN(G1353gat));
  NAND2_X1  g730(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n597_), .A2(new_n932_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(KEYINPUT126), .ZN(new_n934_));
  OR3_X1    g733(.A1(new_n923_), .A2(KEYINPUT127), .A3(new_n934_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n936_));
  OAI21_X1  g735(.A(KEYINPUT127), .B1(new_n923_), .B2(new_n934_), .ZN(new_n937_));
  AND3_X1   g736(.A1(new_n935_), .A2(new_n936_), .A3(new_n937_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n936_), .B1(new_n935_), .B2(new_n937_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n938_), .A2(new_n939_), .ZN(G1354gat));
  INV_X1    g739(.A(G218gat), .ZN(new_n941_));
  NOR3_X1   g740(.A1(new_n923_), .A2(new_n941_), .A3(new_n634_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n924_), .A2(new_n645_), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n942_), .B1(new_n943_), .B2(new_n941_), .ZN(G1355gat));
endmodule


