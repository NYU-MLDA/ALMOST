//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 1 1 1 1 1 0 1 0 1 0 0 0 0 0 0 0 1 0 0 0 1 1 1 1 0 0 1 1 0 0 1 1 1 1 1 0 0 1 1 0 1 0 0 0 0 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n764_, new_n765_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n778_, new_n779_, new_n780_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n805_, new_n806_, new_n807_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n898_, new_n900_,
    new_n902_, new_n903_, new_n905_, new_n906_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n937_, new_n939_,
    new_n940_, new_n941_, new_n943_, new_n944_;
  NAND2_X1  g000(.A1(G141gat), .A2(G148gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT88), .ZN(new_n203_));
  NOR3_X1   g002(.A1(new_n203_), .A2(G141gat), .A3(G148gat), .ZN(new_n204_));
  INV_X1    g003(.A(G141gat), .ZN(new_n205_));
  INV_X1    g004(.A(G148gat), .ZN(new_n206_));
  AOI21_X1  g005(.A(KEYINPUT88), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n202_), .B1(new_n204_), .B2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209_));
  AOI21_X1  g008(.A(KEYINPUT89), .B1(new_n209_), .B2(KEYINPUT1), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n209_), .A2(KEYINPUT89), .A3(KEYINPUT1), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n209_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT1), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n214_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n208_), .B1(new_n213_), .B2(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n215_), .A2(new_n214_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT3), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT90), .ZN(new_n223_));
  NOR2_X1   g022(.A1(G141gat), .A2(G148gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT90), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(new_n225_), .A3(new_n221_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n223_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT2), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n202_), .A2(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n231_));
  AND3_X1   g030(.A1(new_n229_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n220_), .B1(new_n227_), .B2(new_n232_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n218_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT29), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT28), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G22gat), .B(G50gat), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n238_), .A2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n236_), .B(KEYINPUT28), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(new_n239_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  XOR2_X1   g043(.A(G78gat), .B(G106gat), .Z(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT92), .ZN(new_n247_));
  AND2_X1   g046(.A1(G197gat), .A2(G204gat), .ZN(new_n248_));
  NOR2_X1   g047(.A1(G197gat), .A2(G204gat), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n247_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT21), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G211gat), .B(G218gat), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n250_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n253_));
  OR2_X1    g052(.A1(G197gat), .A2(G204gat), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT93), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G197gat), .A2(G204gat), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n254_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT93), .B1(new_n248_), .B2(new_n249_), .ZN(new_n258_));
  INV_X1    g057(.A(G218gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(G211gat), .ZN(new_n260_));
  INV_X1    g059(.A(G211gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(G218gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  AND3_X1   g062(.A1(new_n257_), .A2(new_n258_), .A3(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(KEYINPUT92), .B1(new_n254_), .B2(new_n256_), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT21), .B1(new_n265_), .B2(new_n263_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n253_), .B1(new_n264_), .B2(new_n266_), .ZN(new_n267_));
  XOR2_X1   g066(.A(KEYINPUT94), .B(KEYINPUT29), .Z(new_n268_));
  OAI21_X1  g067(.A(new_n267_), .B1(new_n234_), .B2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(G233gat), .ZN(new_n270_));
  AND2_X1   g069(.A1(new_n270_), .A2(KEYINPUT91), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n270_), .A2(KEYINPUT91), .ZN(new_n272_));
  OAI21_X1  g071(.A(G228gat), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n269_), .A2(new_n274_), .ZN(new_n275_));
  OAI211_X1 g074(.A(new_n273_), .B(new_n267_), .C1(new_n234_), .C2(new_n235_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n246_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  AND3_X1   g076(.A1(new_n275_), .A2(new_n246_), .A3(new_n276_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n244_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n278_), .A2(new_n277_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n280_), .A2(new_n241_), .A3(new_n243_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n279_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT20), .ZN(new_n283_));
  NOR3_X1   g082(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT24), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n285_), .B1(G169gat), .B2(G176gat), .ZN(new_n286_));
  INV_X1    g085(.A(G169gat), .ZN(new_n287_));
  INV_X1    g086(.A(G176gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n284_), .B1(new_n286_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G183gat), .A2(G190gat), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT81), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n293_), .A2(KEYINPUT23), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT23), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n295_), .A2(KEYINPUT81), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n292_), .B1(new_n294_), .B2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n291_), .A2(new_n295_), .ZN(new_n298_));
  INV_X1    g097(.A(G183gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT25), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT25), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(G183gat), .ZN(new_n302_));
  INV_X1    g101(.A(G190gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT26), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT26), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(G190gat), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n300_), .A2(new_n302_), .A3(new_n304_), .A4(new_n306_), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n290_), .A2(new_n297_), .A3(new_n298_), .A4(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(G183gat), .A2(G190gat), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n291_), .B1(new_n294_), .B2(new_n296_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n291_), .A2(KEYINPUT23), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n309_), .B1(new_n310_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G169gat), .A2(G176gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT95), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT95), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n316_), .A2(G169gat), .A3(G176gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(KEYINPUT22), .B(G169gat), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n318_), .B1(new_n320_), .B2(G176gat), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n308_), .B1(new_n313_), .B2(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n283_), .B1(new_n322_), .B2(new_n267_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n309_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT81), .B(KEYINPUT23), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n324_), .B(new_n298_), .C1(new_n325_), .C2(new_n291_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(KEYINPUT83), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT83), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n297_), .A2(new_n328_), .A3(new_n324_), .A4(new_n298_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n314_), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n287_), .A2(KEYINPUT22), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n287_), .A2(KEYINPUT22), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT82), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n287_), .A2(KEYINPUT22), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT82), .ZN(new_n335_));
  AOI21_X1  g134(.A(G176gat), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n330_), .B1(new_n333_), .B2(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n327_), .A2(new_n329_), .A3(new_n337_), .ZN(new_n338_));
  AND3_X1   g137(.A1(new_n250_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n257_), .A2(new_n258_), .A3(new_n263_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n251_), .B1(new_n250_), .B2(new_n252_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n339_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  AND2_X1   g141(.A1(new_n304_), .A2(new_n306_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT80), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n300_), .A2(new_n344_), .ZN(new_n345_));
  AND2_X1   g144(.A1(new_n300_), .A2(new_n302_), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n343_), .B(new_n345_), .C1(new_n346_), .C2(new_n344_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n310_), .A2(new_n312_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n347_), .A2(new_n348_), .A3(new_n290_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n338_), .A2(new_n342_), .A3(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n323_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G226gat), .A2(G233gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT19), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  XOR2_X1   g153(.A(G8gat), .B(G36gat), .Z(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT18), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G64gat), .B(G92gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n338_), .A2(new_n349_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(new_n267_), .ZN(new_n360_));
  AND3_X1   g159(.A1(new_n297_), .A2(new_n307_), .A3(new_n298_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n295_), .A2(KEYINPUT81), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n293_), .A2(KEYINPUT23), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n292_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n324_), .B1(new_n364_), .B2(new_n311_), .ZN(new_n365_));
  AOI22_X1  g164(.A1(new_n319_), .A2(new_n288_), .B1(new_n315_), .B2(new_n317_), .ZN(new_n366_));
  AOI22_X1  g165(.A1(new_n361_), .A2(new_n290_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n283_), .B1(new_n367_), .B2(new_n342_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n353_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n360_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n354_), .A2(new_n358_), .A3(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n351_), .A2(new_n353_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n369_), .B1(new_n360_), .B2(new_n368_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  OAI211_X1 g173(.A(KEYINPUT27), .B(new_n371_), .C1(new_n374_), .C2(new_n358_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT96), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n371_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n358_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n342_), .B1(new_n338_), .B2(new_n349_), .ZN(new_n379_));
  OAI21_X1  g178(.A(KEYINPUT20), .B1(new_n322_), .B2(new_n267_), .ZN(new_n380_));
  NOR3_X1   g179(.A1(new_n379_), .A2(new_n380_), .A3(new_n353_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n369_), .B1(new_n323_), .B2(new_n350_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n378_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n354_), .A2(new_n370_), .A3(KEYINPUT96), .A4(new_n358_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n377_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT105), .ZN(new_n386_));
  XOR2_X1   g185(.A(KEYINPUT104), .B(KEYINPUT27), .Z(new_n387_));
  AND3_X1   g186(.A1(new_n385_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n386_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n375_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT106), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n371_), .A2(new_n376_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n383_), .A2(new_n384_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n387_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(KEYINPUT105), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n385_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n398_), .A2(KEYINPUT106), .A3(new_n375_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n282_), .B1(new_n392_), .B2(new_n399_), .ZN(new_n400_));
  XOR2_X1   g199(.A(KEYINPUT84), .B(G43gat), .Z(new_n401_));
  INV_X1    g200(.A(KEYINPUT85), .ZN(new_n402_));
  INV_X1    g201(.A(G99gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(G71gat), .ZN(new_n404_));
  INV_X1    g203(.A(G71gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(G99gat), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n402_), .B1(new_n404_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(G15gat), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n404_), .A2(new_n406_), .A3(new_n402_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n408_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n410_), .ZN(new_n412_));
  OAI21_X1  g211(.A(G15gat), .B1(new_n412_), .B2(new_n407_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n411_), .A2(new_n413_), .A3(G227gat), .A4(G233gat), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  AOI22_X1  g214(.A1(new_n411_), .A2(new_n413_), .B1(G227gat), .B2(G233gat), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n401_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n416_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n401_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(new_n419_), .A3(new_n414_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n417_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT30), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n359_), .A2(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n338_), .A2(KEYINPUT30), .A3(new_n349_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n423_), .A2(KEYINPUT86), .A3(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(KEYINPUT86), .B1(new_n423_), .B2(new_n424_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n421_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT31), .ZN(new_n429_));
  INV_X1    g228(.A(new_n427_), .ZN(new_n430_));
  NOR3_X1   g229(.A1(new_n415_), .A2(new_n401_), .A3(new_n416_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n419_), .B1(new_n418_), .B2(new_n414_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n430_), .A2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n428_), .A2(new_n429_), .A3(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n429_), .B1(new_n428_), .B2(new_n434_), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT87), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G127gat), .B(G134gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G113gat), .B(G120gat), .ZN(new_n440_));
  XOR2_X1   g239(.A(new_n439_), .B(new_n440_), .Z(new_n441_));
  AOI21_X1  g240(.A(new_n433_), .B1(new_n430_), .B2(new_n425_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n421_), .A2(new_n427_), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT31), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT87), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n444_), .A2(new_n435_), .A3(new_n445_), .ZN(new_n446_));
  AND3_X1   g245(.A1(new_n438_), .A2(new_n441_), .A3(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n441_), .B1(new_n438_), .B2(new_n446_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G225gat), .A2(G233gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(KEYINPUT97), .ZN(new_n450_));
  XOR2_X1   g249(.A(new_n450_), .B(KEYINPUT98), .Z(new_n451_));
  XNOR2_X1  g250(.A(new_n439_), .B(new_n440_), .ZN(new_n452_));
  NOR4_X1   g251(.A1(KEYINPUT90), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n225_), .B1(new_n224_), .B2(new_n221_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n229_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n219_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n212_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n217_), .B1(new_n458_), .B2(new_n210_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n224_), .A2(KEYINPUT88), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n203_), .B1(G141gat), .B2(G148gat), .ZN(new_n461_));
  AOI22_X1  g260(.A1(new_n460_), .A2(new_n461_), .B1(G141gat), .B2(G148gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n459_), .A2(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n452_), .B1(new_n457_), .B2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT4), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n451_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n441_), .B1(new_n218_), .B2(new_n233_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n457_), .A2(new_n463_), .A3(new_n452_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n467_), .A2(KEYINPUT4), .A3(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT99), .ZN(new_n470_));
  AND3_X1   g269(.A1(new_n466_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n470_), .B1(new_n466_), .B2(new_n469_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT102), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G1gat), .B(G29gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(G85gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(KEYINPUT0), .B(G57gat), .ZN(new_n477_));
  XOR2_X1   g276(.A(new_n476_), .B(new_n477_), .Z(new_n478_));
  NAND3_X1  g277(.A1(new_n467_), .A2(new_n468_), .A3(new_n450_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT100), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT100), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n467_), .A2(new_n481_), .A3(new_n468_), .A4(new_n450_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n473_), .A2(new_n474_), .A3(new_n478_), .A4(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n466_), .A2(new_n469_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT99), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n466_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n486_), .A2(new_n483_), .A3(new_n478_), .A4(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT102), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n486_), .A2(new_n483_), .A3(new_n487_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n478_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n484_), .A2(new_n489_), .A3(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT103), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n484_), .A2(new_n489_), .A3(KEYINPUT103), .A4(new_n492_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NOR3_X1   g296(.A1(new_n447_), .A2(new_n448_), .A3(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n495_), .A2(new_n496_), .A3(new_n282_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n473_), .A2(KEYINPUT33), .A3(new_n478_), .A4(new_n483_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT33), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n488_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n467_), .A2(new_n468_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n469_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n450_), .B1(new_n467_), .B2(KEYINPUT4), .ZN(new_n505_));
  OAI221_X1 g304(.A(new_n491_), .B1(new_n503_), .B2(new_n451_), .C1(new_n504_), .C2(new_n505_), .ZN(new_n506_));
  AND3_X1   g305(.A1(new_n500_), .A2(new_n502_), .A3(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n385_), .ZN(new_n508_));
  AND2_X1   g307(.A1(new_n358_), .A2(KEYINPUT32), .ZN(new_n509_));
  NOR3_X1   g308(.A1(new_n381_), .A2(new_n509_), .A3(new_n382_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n509_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(KEYINPUT101), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT101), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n513_), .B(new_n509_), .C1(new_n372_), .C2(new_n373_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n510_), .B1(new_n512_), .B2(new_n514_), .ZN(new_n515_));
  AOI22_X1  g314(.A1(new_n507_), .A2(new_n508_), .B1(new_n493_), .B2(new_n515_), .ZN(new_n516_));
  OAI22_X1  g315(.A1(new_n390_), .A2(new_n499_), .B1(new_n516_), .B2(new_n282_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n438_), .A2(new_n446_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(new_n452_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n438_), .A2(new_n441_), .A3(new_n446_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  AOI22_X1  g320(.A1(new_n400_), .A2(new_n498_), .B1(new_n517_), .B2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT77), .B(G15gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(G22gat), .ZN(new_n524_));
  INV_X1    g323(.A(G1gat), .ZN(new_n525_));
  INV_X1    g324(.A(G8gat), .ZN(new_n526_));
  OAI21_X1  g325(.A(KEYINPUT14), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n524_), .A2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G1gat), .B(G8gat), .ZN(new_n529_));
  OR2_X1    g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n528_), .A2(new_n529_), .ZN(new_n531_));
  AND2_X1   g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G29gat), .B(G36gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G43gat), .B(G50gat), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n533_), .B(new_n534_), .Z(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n532_), .B(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT78), .ZN(new_n538_));
  OR2_X1    g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n537_), .A2(new_n538_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n539_), .A2(G229gat), .A3(G233gat), .A4(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n532_), .ZN(new_n542_));
  XOR2_X1   g341(.A(new_n535_), .B(KEYINPUT15), .Z(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G229gat), .A2(G233gat), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n544_), .B(new_n545_), .C1(new_n542_), .C2(new_n535_), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n541_), .A2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G113gat), .B(G141gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G169gat), .B(G197gat), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n548_), .B(new_n549_), .Z(new_n550_));
  OR2_X1    g349(.A1(new_n547_), .A2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n541_), .A2(new_n546_), .A3(new_n550_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT79), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n541_), .A2(KEYINPUT79), .A3(new_n546_), .A4(new_n550_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n551_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n522_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT107), .ZN(new_n560_));
  XOR2_X1   g359(.A(G120gat), .B(G148gat), .Z(new_n561_));
  XNOR2_X1  g360(.A(G176gat), .B(G204gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n564_));
  XOR2_X1   g363(.A(new_n563_), .B(new_n564_), .Z(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n566_), .A2(KEYINPUT71), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G99gat), .A2(G106gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT6), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT65), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(G85gat), .ZN(new_n573_));
  INV_X1    g372(.A(G92gat), .ZN(new_n574_));
  NOR3_X1   g373(.A1(new_n573_), .A2(new_n574_), .A3(KEYINPUT9), .ZN(new_n575_));
  XOR2_X1   g374(.A(G85gat), .B(G92gat), .Z(new_n576_));
  AOI21_X1  g375(.A(new_n575_), .B1(new_n576_), .B2(KEYINPUT9), .ZN(new_n577_));
  XOR2_X1   g376(.A(KEYINPUT10), .B(G99gat), .Z(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n572_), .B(new_n577_), .C1(G106gat), .C2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT8), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n576_), .A2(new_n581_), .ZN(new_n582_));
  NOR3_X1   g381(.A1(KEYINPUT66), .A2(G99gat), .A3(G106gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT7), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n582_), .B1(new_n572_), .B2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n570_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n581_), .B1(new_n586_), .B2(new_n576_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n580_), .B1(new_n585_), .B2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT67), .ZN(new_n589_));
  XOR2_X1   g388(.A(G57gat), .B(G64gat), .Z(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT68), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT11), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  XOR2_X1   g392(.A(G71gat), .B(G78gat), .Z(new_n594_));
  OR2_X1    g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n591_), .A2(new_n592_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n593_), .A2(new_n596_), .A3(new_n594_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n589_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT12), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n599_), .A2(KEYINPUT12), .A3(new_n588_), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n588_), .B(KEYINPUT67), .Z(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(new_n598_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n602_), .A2(new_n603_), .A3(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(G230gat), .A2(G233gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT64), .ZN(new_n608_));
  OAI21_X1  g407(.A(KEYINPUT70), .B1(new_n606_), .B2(new_n608_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n605_), .A2(new_n603_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT70), .ZN(new_n611_));
  INV_X1    g410(.A(new_n608_), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n610_), .A2(new_n611_), .A3(new_n612_), .A4(new_n602_), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n609_), .A2(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n612_), .B1(new_n605_), .B2(new_n600_), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n615_), .B(KEYINPUT69), .Z(new_n616_));
  AOI21_X1  g415(.A(new_n568_), .B1(new_n614_), .B2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n614_), .A2(new_n616_), .A3(new_n568_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n618_), .A2(KEYINPUT13), .A3(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT13), .ZN(new_n621_));
  INV_X1    g420(.A(new_n619_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n621_), .B1(new_n622_), .B2(new_n617_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n620_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(G231gat), .A2(G233gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n532_), .B(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(new_n598_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G127gat), .B(G155gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT16), .ZN(new_n629_));
  XOR2_X1   g428(.A(G183gat), .B(G211gat), .Z(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT17), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n631_), .A2(new_n632_), .ZN(new_n634_));
  NOR3_X1   g433(.A1(new_n627_), .A2(new_n633_), .A3(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n635_), .B1(new_n633_), .B2(new_n627_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(G232gat), .A2(G233gat), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT34), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(KEYINPUT35), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n640_), .A2(KEYINPUT74), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n639_), .A2(KEYINPUT35), .ZN(new_n642_));
  AOI211_X1 g441(.A(new_n641_), .B(new_n642_), .C1(new_n588_), .C2(new_n543_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n643_), .B1(new_n589_), .B2(new_n535_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n640_), .A2(KEYINPUT74), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n644_), .A2(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n644_), .A2(new_n646_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(G190gat), .B(G218gat), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT73), .ZN(new_n651_));
  XNOR2_X1  g450(.A(G134gat), .B(G162gat), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n651_), .B(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT36), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT75), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n649_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT36), .ZN(new_n657_));
  OAI211_X1 g456(.A(new_n657_), .B(new_n653_), .C1(new_n647_), .C2(new_n648_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(KEYINPUT37), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n649_), .A2(new_n654_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(new_n658_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(KEYINPUT76), .B(KEYINPUT37), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n660_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NOR3_X1   g464(.A1(new_n624_), .A2(new_n637_), .A3(new_n665_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n560_), .A2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n667_), .A2(new_n525_), .A3(new_n497_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT38), .ZN(new_n669_));
  OR2_X1    g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n624_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n662_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n522_), .A2(new_n672_), .ZN(new_n673_));
  NAND4_X1  g472(.A1(new_n671_), .A2(new_n557_), .A3(new_n636_), .A4(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n497_), .ZN(new_n675_));
  OAI21_X1  g474(.A(G1gat), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n668_), .A2(new_n669_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n670_), .A2(new_n676_), .A3(new_n677_), .ZN(G1324gat));
  NAND2_X1  g477(.A1(new_n392_), .A2(new_n399_), .ZN(new_n679_));
  OR3_X1    g478(.A1(new_n674_), .A2(KEYINPUT109), .A3(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(KEYINPUT109), .B1(new_n674_), .B2(new_n679_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n680_), .A2(G8gat), .A3(new_n681_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT39), .ZN(new_n683_));
  INV_X1    g482(.A(new_n679_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n667_), .A2(new_n526_), .A3(new_n684_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT108), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n683_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT40), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n687_), .B(new_n688_), .ZN(G1325gat));
  OAI21_X1  g488(.A(G15gat), .B1(new_n674_), .B2(new_n521_), .ZN(new_n690_));
  XOR2_X1   g489(.A(new_n690_), .B(KEYINPUT41), .Z(new_n691_));
  INV_X1    g490(.A(new_n521_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n667_), .A2(new_n409_), .A3(new_n692_), .ZN(new_n693_));
  OR2_X1    g492(.A1(new_n693_), .A2(KEYINPUT110), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(KEYINPUT110), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n691_), .A2(new_n694_), .A3(new_n695_), .ZN(G1326gat));
  INV_X1    g495(.A(new_n282_), .ZN(new_n697_));
  OAI21_X1  g496(.A(G22gat), .B1(new_n674_), .B2(new_n697_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT42), .ZN(new_n699_));
  INV_X1    g498(.A(new_n667_), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n697_), .A2(G22gat), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n699_), .B1(new_n700_), .B2(new_n701_), .ZN(G1327gat));
  NOR2_X1   g501(.A1(new_n636_), .A2(new_n662_), .ZN(new_n703_));
  AND3_X1   g502(.A1(new_n560_), .A2(new_n671_), .A3(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(G29gat), .B1(new_n704_), .B2(new_n497_), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n522_), .A2(KEYINPUT43), .A3(new_n664_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT113), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT43), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n517_), .A2(new_n521_), .ZN(new_n710_));
  AOI21_X1  g509(.A(KEYINPUT106), .B1(new_n398_), .B2(new_n375_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n375_), .ZN(new_n712_));
  AOI211_X1 g511(.A(new_n391_), .B(new_n712_), .C1(new_n396_), .C2(new_n397_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n697_), .B1(new_n711_), .B2(new_n713_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n519_), .A2(new_n675_), .A3(new_n520_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n710_), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT112), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n664_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  OAI211_X1 g517(.A(new_n710_), .B(KEYINPUT112), .C1(new_n714_), .C2(new_n715_), .ZN(new_n719_));
  AOI211_X1 g518(.A(new_n708_), .B(new_n709_), .C1(new_n718_), .C2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n716_), .A2(new_n717_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n721_), .A2(new_n665_), .A3(new_n719_), .ZN(new_n722_));
  AOI21_X1  g521(.A(KEYINPUT113), .B1(new_n722_), .B2(KEYINPUT43), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n707_), .B1(new_n720_), .B2(new_n723_), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n620_), .A2(new_n623_), .A3(new_n557_), .A4(new_n637_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT111), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n725_), .B(new_n726_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n724_), .A2(KEYINPUT44), .A3(new_n727_), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n728_), .A2(G29gat), .A3(new_n497_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n665_), .B1(new_n522_), .B2(KEYINPUT112), .ZN(new_n731_));
  INV_X1    g530(.A(new_n719_), .ZN(new_n732_));
  OAI21_X1  g531(.A(KEYINPUT43), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(new_n708_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n722_), .A2(KEYINPUT113), .A3(KEYINPUT43), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n706_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n725_), .B(KEYINPUT111), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n730_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n705_), .B1(new_n729_), .B2(new_n738_), .ZN(G1328gat));
  INV_X1    g538(.A(G36gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n704_), .A2(new_n740_), .A3(new_n684_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT45), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n738_), .A2(new_n684_), .A3(new_n728_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT114), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n743_), .A2(new_n744_), .A3(G36gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n743_), .B2(G36gat), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n742_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT46), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  OAI211_X1 g548(.A(KEYINPUT46), .B(new_n742_), .C1(new_n745_), .C2(new_n746_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1329gat));
  NAND2_X1  g550(.A1(new_n704_), .A2(new_n692_), .ZN(new_n752_));
  INV_X1    g551(.A(G43gat), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n521_), .A2(new_n753_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n728_), .A2(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(KEYINPUT115), .B1(new_n756_), .B2(new_n738_), .ZN(new_n757_));
  AND4_X1   g556(.A1(KEYINPUT115), .A2(new_n738_), .A3(new_n728_), .A4(new_n755_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n754_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(KEYINPUT47), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT47), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n761_), .B(new_n754_), .C1(new_n757_), .C2(new_n758_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(G1330gat));
  AOI21_X1  g562(.A(G50gat), .B1(new_n704_), .B2(new_n282_), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n728_), .A2(G50gat), .A3(new_n282_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n765_), .B2(new_n738_), .ZN(G1331gat));
  INV_X1    g565(.A(G57gat), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n665_), .A2(new_n637_), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n624_), .A2(new_n768_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n522_), .A2(new_n557_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n767_), .B1(new_n771_), .B2(new_n675_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT116), .ZN(new_n773_));
  NOR3_X1   g572(.A1(new_n671_), .A2(new_n557_), .A3(new_n637_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n673_), .ZN(new_n775_));
  NOR3_X1   g574(.A1(new_n775_), .A2(new_n767_), .A3(new_n675_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n773_), .A2(new_n776_), .ZN(G1332gat));
  OAI21_X1  g576(.A(G64gat), .B1(new_n775_), .B2(new_n679_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT48), .ZN(new_n779_));
  OR2_X1    g578(.A1(new_n679_), .A2(G64gat), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n779_), .B1(new_n771_), .B2(new_n780_), .ZN(G1333gat));
  INV_X1    g580(.A(KEYINPUT49), .ZN(new_n782_));
  INV_X1    g581(.A(new_n775_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n692_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n782_), .B1(new_n784_), .B2(G71gat), .ZN(new_n785_));
  AOI211_X1 g584(.A(KEYINPUT49), .B(new_n405_), .C1(new_n783_), .C2(new_n692_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n692_), .A2(new_n405_), .ZN(new_n787_));
  OAI22_X1  g586(.A1(new_n785_), .A2(new_n786_), .B1(new_n771_), .B2(new_n787_), .ZN(new_n788_));
  XOR2_X1   g587(.A(new_n788_), .B(KEYINPUT117), .Z(G1334gat));
  OR3_X1    g588(.A1(new_n771_), .A2(G78gat), .A3(new_n697_), .ZN(new_n790_));
  OAI21_X1  g589(.A(G78gat), .B1(new_n775_), .B2(new_n697_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(KEYINPUT118), .B(KEYINPUT50), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n792_), .A2(new_n793_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n790_), .B1(new_n794_), .B2(new_n795_), .ZN(G1335gat));
  AND2_X1   g595(.A1(new_n624_), .A2(new_n703_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n770_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n573_), .B1(new_n798_), .B2(new_n675_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n799_), .B(KEYINPUT119), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n624_), .A2(new_n558_), .A3(new_n637_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n736_), .A2(new_n801_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n675_), .A2(new_n573_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n800_), .B1(new_n802_), .B2(new_n803_), .ZN(G1336gat));
  NOR3_X1   g603(.A1(new_n798_), .A2(G92gat), .A3(new_n679_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n802_), .A2(new_n684_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n805_), .B1(new_n806_), .B2(G92gat), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n807_), .B(KEYINPUT120), .ZN(G1337gat));
  NAND4_X1  g607(.A1(new_n797_), .A2(new_n692_), .A3(new_n578_), .A4(new_n770_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT51), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n736_), .A2(new_n521_), .A3(new_n801_), .ZN(new_n811_));
  OAI221_X1 g610(.A(new_n809_), .B1(KEYINPUT121), .B2(new_n810_), .C1(new_n811_), .C2(new_n403_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(KEYINPUT121), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n812_), .B(new_n813_), .ZN(G1338gat));
  XNOR2_X1  g613(.A(KEYINPUT122), .B(KEYINPUT53), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n802_), .A2(new_n282_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(G106gat), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(KEYINPUT52), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT52), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n816_), .A2(new_n819_), .A3(G106gat), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n820_), .ZN(new_n821_));
  NOR3_X1   g620(.A1(new_n798_), .A2(G106gat), .A3(new_n697_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n815_), .B1(new_n821_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n815_), .ZN(new_n825_));
  AOI211_X1 g624(.A(new_n822_), .B(new_n825_), .C1(new_n818_), .C2(new_n820_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n824_), .A2(new_n826_), .ZN(G1339gat));
  NAND3_X1  g626(.A1(new_n671_), .A2(new_n558_), .A3(new_n768_), .ZN(new_n828_));
  XOR2_X1   g627(.A(new_n828_), .B(KEYINPUT54), .Z(new_n829_));
  NAND3_X1  g628(.A1(new_n614_), .A2(new_n616_), .A3(new_n566_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n539_), .A2(new_n545_), .A3(new_n540_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n545_), .B1(new_n532_), .B2(new_n536_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n550_), .B1(new_n544_), .B2(new_n832_), .ZN(new_n833_));
  AOI22_X1  g632(.A1(new_n554_), .A2(new_n555_), .B1(new_n831_), .B2(new_n833_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n830_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT55), .ZN(new_n836_));
  NOR3_X1   g635(.A1(new_n606_), .A2(new_n836_), .A3(new_n608_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n612_), .B1(new_n610_), .B2(new_n602_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n609_), .A2(new_n613_), .A3(new_n836_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(KEYINPUT56), .B1(new_n841_), .B2(new_n565_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT56), .ZN(new_n843_));
  AOI211_X1 g642(.A(new_n843_), .B(new_n566_), .C1(new_n839_), .C2(new_n840_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n835_), .B1(new_n842_), .B2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT58), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n835_), .B(KEYINPUT58), .C1(new_n842_), .C2(new_n844_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n847_), .A2(new_n665_), .A3(new_n848_), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n557_), .B(new_n830_), .C1(new_n842_), .C2(new_n844_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n834_), .B1(new_n622_), .B2(new_n617_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n672_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n849_), .B1(KEYINPUT57), .B2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(KEYINPUT123), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT123), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n849_), .B(new_n855_), .C1(KEYINPUT57), .C2(new_n852_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n852_), .A2(KEYINPUT57), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n854_), .A2(new_n856_), .A3(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n829_), .B1(new_n858_), .B2(new_n637_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n521_), .A2(new_n675_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n400_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n861_), .A2(KEYINPUT59), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  OAI21_X1  g662(.A(KEYINPUT124), .B1(new_n859_), .B2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT124), .ZN(new_n865_));
  INV_X1    g664(.A(new_n857_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n866_), .B1(new_n853_), .B2(KEYINPUT123), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n636_), .B1(new_n867_), .B2(new_n856_), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n865_), .B(new_n862_), .C1(new_n868_), .C2(new_n829_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n637_), .B1(new_n853_), .B2(new_n866_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n828_), .B(KEYINPUT54), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n861_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(KEYINPUT59), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n864_), .A2(new_n869_), .A3(new_n557_), .A4(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(G113gat), .ZN(new_n877_));
  OR3_X1    g676(.A1(new_n874_), .A2(G113gat), .A3(new_n558_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(G1340gat));
  NAND4_X1  g678(.A1(new_n864_), .A2(new_n869_), .A3(new_n624_), .A4(new_n875_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(G120gat), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT60), .ZN(new_n882_));
  AOI21_X1  g681(.A(G120gat), .B1(new_n624_), .B2(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n883_), .B1(new_n882_), .B2(G120gat), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n872_), .A2(new_n873_), .A3(new_n884_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(KEYINPUT125), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n881_), .A2(new_n886_), .ZN(G1341gat));
  NAND4_X1  g686(.A1(new_n864_), .A2(new_n869_), .A3(new_n636_), .A4(new_n875_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(G127gat), .ZN(new_n889_));
  OR3_X1    g688(.A1(new_n874_), .A2(G127gat), .A3(new_n637_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(G1342gat));
  NAND4_X1  g690(.A1(new_n864_), .A2(new_n869_), .A3(new_n665_), .A4(new_n875_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(G134gat), .ZN(new_n893_));
  OR3_X1    g692(.A1(new_n874_), .A2(G134gat), .A3(new_n662_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(G1343gat));
  NOR3_X1   g694(.A1(new_n692_), .A2(new_n675_), .A3(new_n697_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n872_), .A2(new_n679_), .A3(new_n896_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n897_), .A2(new_n558_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(new_n205_), .ZN(G1344gat));
  NOR2_X1   g698(.A1(new_n897_), .A2(new_n671_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(new_n206_), .ZN(G1345gat));
  NOR2_X1   g700(.A1(new_n897_), .A2(new_n637_), .ZN(new_n902_));
  XOR2_X1   g701(.A(KEYINPUT61), .B(G155gat), .Z(new_n903_));
  XNOR2_X1  g702(.A(new_n902_), .B(new_n903_), .ZN(G1346gat));
  OAI21_X1  g703(.A(G162gat), .B1(new_n897_), .B2(new_n664_), .ZN(new_n905_));
  OR2_X1    g704(.A1(new_n662_), .A2(G162gat), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n905_), .B1(new_n897_), .B2(new_n906_), .ZN(G1347gat));
  NOR3_X1   g706(.A1(new_n679_), .A2(new_n715_), .A3(new_n282_), .ZN(new_n908_));
  OAI211_X1 g707(.A(new_n557_), .B(new_n908_), .C1(new_n868_), .C2(new_n829_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(G169gat), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT62), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n909_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n913_));
  OAI211_X1 g712(.A(new_n912_), .B(new_n913_), .C1(new_n320_), .C2(new_n909_), .ZN(G1348gat));
  NOR2_X1   g713(.A1(new_n679_), .A2(new_n715_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n624_), .A2(G176gat), .A3(new_n915_), .ZN(new_n916_));
  AOI211_X1 g715(.A(new_n282_), .B(new_n916_), .C1(new_n870_), .C2(new_n871_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n859_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n918_), .A2(new_n624_), .A3(new_n908_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n917_), .B1(new_n919_), .B2(new_n288_), .ZN(G1349gat));
  NAND2_X1  g719(.A1(new_n918_), .A2(new_n908_), .ZN(new_n921_));
  NOR3_X1   g720(.A1(new_n921_), .A2(new_n346_), .A3(new_n637_), .ZN(new_n922_));
  NAND4_X1  g721(.A1(new_n872_), .A2(new_n697_), .A3(new_n636_), .A4(new_n915_), .ZN(new_n923_));
  AND2_X1   g722(.A1(new_n923_), .A2(new_n299_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n922_), .A2(new_n924_), .ZN(G1350gat));
  OAI211_X1 g724(.A(new_n665_), .B(new_n908_), .C1(new_n868_), .C2(new_n829_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT126), .ZN(new_n927_));
  AND3_X1   g726(.A1(new_n926_), .A2(new_n927_), .A3(G190gat), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n927_), .B1(new_n926_), .B2(G190gat), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n672_), .A2(new_n343_), .ZN(new_n930_));
  OAI22_X1  g729(.A1(new_n928_), .A2(new_n929_), .B1(new_n921_), .B2(new_n930_), .ZN(G1351gat));
  NOR3_X1   g730(.A1(new_n692_), .A2(new_n679_), .A3(new_n499_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n872_), .A2(new_n932_), .ZN(new_n933_));
  INV_X1    g732(.A(new_n933_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(new_n557_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g735(.A1(new_n934_), .A2(new_n624_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g737(.A(KEYINPUT63), .B(G211gat), .C1(new_n934_), .C2(new_n636_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(KEYINPUT63), .B(G211gat), .ZN(new_n940_));
  NOR3_X1   g739(.A1(new_n933_), .A2(new_n637_), .A3(new_n940_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n939_), .A2(new_n941_), .ZN(G1354gat));
  OAI21_X1  g741(.A(G218gat), .B1(new_n933_), .B2(new_n664_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n672_), .A2(new_n259_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n943_), .B1(new_n933_), .B2(new_n944_), .ZN(G1355gat));
endmodule


