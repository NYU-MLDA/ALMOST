//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 0 0 0 0 1 0 0 0 1 0 1 0 1 0 1 1 1 1 1 1 0 1 0 0 0 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n584_, new_n586_, new_n587_, new_n588_,
    new_n589_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n656_, new_n657_, new_n658_, new_n659_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n815_, new_n816_, new_n817_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n827_, new_n829_,
    new_n830_, new_n832_, new_n833_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n845_, new_n846_, new_n847_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n855_, new_n856_, new_n857_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT85), .ZN(new_n205_));
  XOR2_X1   g004(.A(KEYINPUT84), .B(KEYINPUT30), .Z(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT23), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n209_), .B1(G183gat), .B2(G190gat), .ZN(new_n210_));
  INV_X1    g009(.A(G169gat), .ZN(new_n211_));
  INV_X1    g010(.A(G176gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT83), .ZN(new_n215_));
  NOR3_X1   g014(.A1(new_n215_), .A2(new_n211_), .A3(KEYINPUT22), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT22), .B1(new_n215_), .B2(new_n211_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(new_n212_), .ZN(new_n218_));
  OAI211_X1 g017(.A(new_n210_), .B(new_n214_), .C1(new_n216_), .C2(new_n218_), .ZN(new_n219_));
  NOR3_X1   g018(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT25), .B(G183gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT26), .B(G190gat), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n220_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n224_));
  OAI211_X1 g023(.A(new_n223_), .B(new_n209_), .C1(new_n213_), .C2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n219_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n207_), .B(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n228_), .B(G43gat), .ZN(new_n229_));
  XOR2_X1   g028(.A(KEYINPUT86), .B(KEYINPUT31), .Z(new_n230_));
  XNOR2_X1  g029(.A(G71gat), .B(G99gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n230_), .B(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G227gat), .A2(G233gat), .ZN(new_n233_));
  INV_X1    g032(.A(G15gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n232_), .B(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n229_), .B(new_n236_), .ZN(new_n237_));
  XOR2_X1   g036(.A(G78gat), .B(G106gat), .Z(new_n238_));
  INV_X1    g037(.A(KEYINPUT87), .ZN(new_n239_));
  OAI22_X1  g038(.A1(new_n239_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n240_), .B1(KEYINPUT87), .B2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G141gat), .A2(G148gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT2), .ZN(new_n244_));
  OR2_X1    g043(.A1(G141gat), .A2(G148gat), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n245_), .A2(new_n239_), .A3(KEYINPUT3), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n242_), .A2(new_n244_), .A3(new_n246_), .ZN(new_n247_));
  OR2_X1    g046(.A1(G155gat), .A2(G162gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G155gat), .A2(G162gat), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n247_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(KEYINPUT1), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(new_n248_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n249_), .A2(KEYINPUT1), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n245_), .B(new_n243_), .C1(new_n252_), .C2(new_n253_), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n250_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT29), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT28), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(G22gat), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT28), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n257_), .B(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(G22gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  AND3_X1   g062(.A1(new_n259_), .A2(new_n263_), .A3(G50gat), .ZN(new_n264_));
  AOI21_X1  g063(.A(G50gat), .B1(new_n259_), .B2(new_n263_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n238_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G228gat), .A2(G233gat), .ZN(new_n267_));
  XOR2_X1   g066(.A(new_n267_), .B(KEYINPUT90), .Z(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(G50gat), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n261_), .A2(new_n262_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n258_), .A2(G22gat), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n270_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n259_), .A2(new_n263_), .A3(G50gat), .ZN(new_n274_));
  INV_X1    g073(.A(new_n238_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(KEYINPUT89), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n273_), .A2(new_n274_), .A3(new_n277_), .ZN(new_n278_));
  AND3_X1   g077(.A1(new_n266_), .A2(new_n269_), .A3(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n269_), .B1(new_n266_), .B2(new_n278_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G197gat), .A2(G204gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT88), .B(G197gat), .ZN(new_n282_));
  OAI211_X1 g081(.A(KEYINPUT21), .B(new_n281_), .C1(new_n282_), .C2(G204gat), .ZN(new_n283_));
  XOR2_X1   g082(.A(G211gat), .B(G218gat), .Z(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(G204gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(G197gat), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n287_), .B1(new_n282_), .B2(new_n286_), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n283_), .B(new_n285_), .C1(new_n288_), .C2(KEYINPUT21), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n288_), .A2(KEYINPUT21), .A3(new_n284_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n250_), .A2(new_n254_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n292_), .B1(KEYINPUT29), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NOR3_X1   g094(.A1(new_n279_), .A2(new_n280_), .A3(new_n295_), .ZN(new_n296_));
  NOR3_X1   g095(.A1(new_n264_), .A2(new_n265_), .A3(new_n276_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n275_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n268_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n266_), .A2(new_n278_), .A3(new_n269_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n294_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n205_), .A2(new_n255_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n302_), .A2(KEYINPUT4), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT91), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n255_), .A2(new_n204_), .ZN(new_n306_));
  OAI21_X1  g105(.A(KEYINPUT91), .B1(new_n205_), .B2(new_n255_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n305_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n303_), .B1(new_n308_), .B2(KEYINPUT4), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G225gat), .A2(G233gat), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  OR2_X1    g110(.A1(new_n309_), .A2(new_n311_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n308_), .A2(new_n310_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G1gat), .B(G29gat), .ZN(new_n314_));
  INV_X1    g113(.A(G85gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT0), .B(G57gat), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n316_), .B(new_n317_), .Z(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n313_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n312_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n226_), .A2(new_n291_), .ZN(new_n322_));
  XOR2_X1   g121(.A(KEYINPUT22), .B(G169gat), .Z(new_n323_));
  OAI211_X1 g122(.A(new_n210_), .B(new_n214_), .C1(G176gat), .C2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(new_n225_), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n322_), .B(KEYINPUT20), .C1(new_n291_), .C2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n291_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT20), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n328_), .B1(new_n292_), .B2(new_n227_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G226gat), .A2(G233gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT19), .ZN(new_n331_));
  MUX2_X1   g130(.A(new_n326_), .B(new_n329_), .S(new_n331_), .Z(new_n332_));
  XNOR2_X1  g131(.A(G8gat), .B(G36gat), .ZN(new_n333_));
  INV_X1    g132(.A(G92gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT18), .B(G64gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n332_), .A2(new_n337_), .ZN(new_n338_));
  OR2_X1    g137(.A1(new_n332_), .A2(new_n337_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n321_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  OR3_X1    g139(.A1(new_n308_), .A2(KEYINPUT92), .A3(new_n311_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n309_), .A2(new_n310_), .ZN(new_n342_));
  OAI21_X1  g141(.A(KEYINPUT92), .B1(new_n308_), .B2(new_n311_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n341_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(new_n319_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT33), .ZN(new_n346_));
  INV_X1    g145(.A(new_n343_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n347_), .B1(new_n310_), .B2(new_n309_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n318_), .B1(new_n348_), .B2(new_n341_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT33), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n340_), .B1(new_n346_), .B2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n337_), .A2(KEYINPUT32), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n332_), .A2(new_n353_), .ZN(new_n354_));
  AOI211_X1 g153(.A(new_n331_), .B(new_n328_), .C1(new_n292_), .C2(new_n227_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n355_), .B1(new_n331_), .B2(new_n326_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n354_), .B1(new_n353_), .B2(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n348_), .A2(new_n318_), .A3(new_n341_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n357_), .B1(new_n345_), .B2(new_n358_), .ZN(new_n359_));
  OAI22_X1  g158(.A1(new_n296_), .A2(new_n301_), .B1(new_n352_), .B2(new_n359_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n344_), .A2(new_n319_), .ZN(new_n361_));
  OAI21_X1  g160(.A(KEYINPUT93), .B1(new_n361_), .B2(new_n349_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT93), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n345_), .A2(new_n358_), .A3(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n339_), .A2(new_n338_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT27), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  XOR2_X1   g167(.A(new_n337_), .B(KEYINPUT94), .Z(new_n369_));
  OAI211_X1 g168(.A(new_n338_), .B(KEYINPUT27), .C1(new_n356_), .C2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n295_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n299_), .A2(new_n294_), .A3(new_n300_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n365_), .A2(new_n372_), .A3(new_n373_), .A4(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n237_), .B1(new_n360_), .B2(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n296_), .A2(new_n301_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n365_), .A2(new_n237_), .ZN(new_n378_));
  NOR3_X1   g177(.A1(new_n377_), .A2(new_n378_), .A3(new_n371_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n376_), .A2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G15gat), .B(G22gat), .ZN(new_n381_));
  INV_X1    g180(.A(G1gat), .ZN(new_n382_));
  INV_X1    g181(.A(G8gat), .ZN(new_n383_));
  OAI21_X1  g182(.A(KEYINPUT14), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n381_), .A2(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G1gat), .B(G8gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G29gat), .B(G36gat), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G43gat), .B(G50gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n390_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(new_n388_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n391_), .A2(new_n393_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n387_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT15), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n394_), .B(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n395_), .B1(new_n397_), .B2(new_n387_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G229gat), .A2(G233gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT80), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n398_), .A2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n387_), .B(new_n394_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n403_), .A2(G229gat), .A3(G233gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G169gat), .B(G197gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(KEYINPUT81), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G113gat), .B(G141gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n402_), .A2(new_n404_), .A3(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT82), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n409_), .B1(new_n402_), .B2(new_n404_), .ZN(new_n413_));
  OR3_X1    g212(.A1(new_n411_), .A2(new_n412_), .A3(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n412_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT8), .ZN(new_n418_));
  AND2_X1   g217(.A1(G85gat), .A2(G92gat), .ZN(new_n419_));
  NOR2_X1   g218(.A1(G85gat), .A2(G92gat), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT69), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n315_), .A2(new_n334_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT69), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G85gat), .A2(G92gat), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n422_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n421_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT7), .ZN(new_n427_));
  INV_X1    g226(.A(G99gat), .ZN(new_n428_));
  INV_X1    g227(.A(G106gat), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n427_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(G99gat), .A2(G106gat), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT6), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n430_), .A2(new_n433_), .A3(new_n434_), .A4(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n418_), .B1(new_n426_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT68), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(KEYINPUT8), .B1(new_n421_), .B2(new_n425_), .ZN(new_n440_));
  AND3_X1   g239(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n441_));
  AOI21_X1  g240(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n443_), .A2(KEYINPUT68), .A3(new_n435_), .A4(new_n430_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n439_), .A2(new_n440_), .A3(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT70), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT70), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n439_), .A2(new_n440_), .A3(new_n444_), .A4(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n437_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n449_));
  XOR2_X1   g248(.A(KEYINPUT10), .B(G99gat), .Z(new_n450_));
  XNOR2_X1  g249(.A(KEYINPUT65), .B(G106gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  OR2_X1    g251(.A1(new_n452_), .A2(KEYINPUT66), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT9), .ZN(new_n454_));
  OR3_X1    g253(.A1(new_n424_), .A2(new_n454_), .A3(KEYINPUT67), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n420_), .B1(new_n454_), .B2(new_n424_), .ZN(new_n456_));
  OAI21_X1  g255(.A(KEYINPUT67), .B1(new_n424_), .B2(new_n454_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n455_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n452_), .A2(KEYINPUT66), .ZN(new_n459_));
  AND4_X1   g258(.A1(new_n443_), .A2(new_n453_), .A3(new_n458_), .A4(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(G57gat), .ZN(new_n461_));
  INV_X1    g260(.A(G64gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT11), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G57gat), .A2(G64gat), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n463_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n466_));
  AND2_X1   g265(.A1(G71gat), .A2(G78gat), .ZN(new_n467_));
  NOR2_X1   g266(.A1(G71gat), .A2(G78gat), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n466_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT71), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n464_), .B1(new_n463_), .B2(new_n465_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT71), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n466_), .A2(new_n473_), .A3(new_n469_), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n471_), .A2(new_n472_), .A3(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n472_), .B1(new_n471_), .B2(new_n474_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NOR3_X1   g276(.A1(new_n449_), .A2(new_n460_), .A3(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n477_), .B1(new_n449_), .B2(new_n460_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(KEYINPUT72), .B(KEYINPUT12), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n478_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G230gat), .A2(G233gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT64), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  OAI211_X1 g283(.A(KEYINPUT12), .B(new_n477_), .C1(new_n449_), .C2(new_n460_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n481_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  OR3_X1    g285(.A1(new_n449_), .A2(new_n460_), .A3(new_n477_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(new_n479_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(new_n483_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n486_), .A2(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(G120gat), .B(G148gat), .Z(new_n491_));
  XNOR2_X1  g290(.A(KEYINPUT75), .B(KEYINPUT76), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G176gat), .B(G204gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(KEYINPUT74), .B(KEYINPUT5), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n498_), .A2(KEYINPUT73), .ZN(new_n499_));
  XOR2_X1   g298(.A(new_n490_), .B(new_n499_), .Z(new_n500_));
  OR2_X1    g299(.A1(new_n500_), .A2(KEYINPUT13), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(KEYINPUT13), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NOR3_X1   g302(.A1(new_n380_), .A2(new_n417_), .A3(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G190gat), .B(G218gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G134gat), .B(G162gat), .ZN(new_n506_));
  XOR2_X1   g305(.A(new_n505_), .B(new_n506_), .Z(new_n507_));
  INV_X1    g306(.A(KEYINPUT36), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  OR2_X1    g308(.A1(new_n507_), .A2(new_n508_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n397_), .B1(new_n449_), .B2(new_n460_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NOR3_X1   g311(.A1(new_n449_), .A2(new_n460_), .A3(new_n394_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G232gat), .A2(G233gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT34), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT35), .ZN(new_n517_));
  AND2_X1   g316(.A1(new_n517_), .A2(KEYINPUT78), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n517_), .A2(KEYINPUT78), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n516_), .A2(KEYINPUT35), .ZN(new_n520_));
  NOR3_X1   g319(.A1(new_n518_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n514_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n513_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n517_), .B1(new_n523_), .B2(new_n511_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n522_), .B1(new_n524_), .B2(KEYINPUT77), .ZN(new_n525_));
  OAI211_X1 g324(.A(KEYINPUT35), .B(new_n516_), .C1(new_n512_), .C2(new_n513_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT77), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n509_), .B(new_n510_), .C1(new_n525_), .C2(new_n528_), .ZN(new_n529_));
  AOI22_X1  g328(.A1(new_n526_), .A2(new_n527_), .B1(new_n514_), .B2(new_n521_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n524_), .A2(KEYINPUT77), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n530_), .A2(new_n508_), .A3(new_n507_), .A4(new_n531_), .ZN(new_n532_));
  XOR2_X1   g331(.A(KEYINPUT79), .B(KEYINPUT37), .Z(new_n533_));
  AND3_X1   g332(.A1(new_n529_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n533_), .B1(new_n529_), .B2(new_n532_), .ZN(new_n535_));
  OR2_X1    g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G231gat), .A2(G233gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n387_), .B(new_n537_), .ZN(new_n538_));
  XOR2_X1   g337(.A(new_n538_), .B(new_n477_), .Z(new_n539_));
  XOR2_X1   g338(.A(G127gat), .B(G155gat), .Z(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(G211gat), .ZN(new_n541_));
  XOR2_X1   g340(.A(KEYINPUT16), .B(G183gat), .Z(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT17), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n543_), .A2(KEYINPUT17), .ZN(new_n545_));
  AND3_X1   g344(.A1(new_n539_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n539_), .A2(new_n544_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n536_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n504_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n365_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n552_), .A2(new_n382_), .A3(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT38), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n529_), .A2(new_n532_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n557_), .A2(new_n549_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n504_), .A2(new_n558_), .ZN(new_n559_));
  OAI21_X1  g358(.A(G1gat), .B1(new_n559_), .B2(new_n365_), .ZN(new_n560_));
  OR2_X1    g359(.A1(new_n560_), .A2(KEYINPUT95), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(KEYINPUT95), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n555_), .A2(new_n561_), .A3(new_n562_), .ZN(G1324gat));
  NAND3_X1  g362(.A1(new_n552_), .A2(new_n383_), .A3(new_n371_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n504_), .A2(new_n371_), .A3(new_n558_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(G8gat), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(KEYINPUT39), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(KEYINPUT96), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT96), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n566_), .A2(new_n569_), .A3(KEYINPUT39), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT39), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n565_), .A2(new_n572_), .A3(G8gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT97), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n564_), .B1(new_n571_), .B2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT40), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  OAI211_X1 g376(.A(KEYINPUT40), .B(new_n564_), .C1(new_n571_), .C2(new_n574_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(G1325gat));
  INV_X1    g378(.A(new_n237_), .ZN(new_n580_));
  OAI21_X1  g379(.A(G15gat), .B1(new_n559_), .B2(new_n580_), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n581_), .A2(KEYINPUT41), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(KEYINPUT41), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n552_), .A2(new_n234_), .A3(new_n237_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n582_), .A2(new_n583_), .A3(new_n584_), .ZN(G1326gat));
  INV_X1    g384(.A(new_n377_), .ZN(new_n586_));
  OAI21_X1  g385(.A(G22gat), .B1(new_n559_), .B2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT42), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n552_), .A2(new_n262_), .A3(new_n377_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(G1327gat));
  NOR2_X1   g389(.A1(new_n556_), .A2(new_n548_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n504_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(G29gat), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n593_), .A2(new_n594_), .A3(new_n553_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n534_), .A2(new_n535_), .ZN(new_n596_));
  AND4_X1   g395(.A1(new_n365_), .A2(new_n374_), .A3(new_n372_), .A4(new_n373_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n346_), .A2(new_n351_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n340_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n359_), .ZN(new_n601_));
  AOI22_X1  g400(.A1(new_n600_), .A2(new_n601_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n580_), .B1(new_n597_), .B2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n378_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n586_), .A2(new_n604_), .A3(new_n372_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n596_), .B1(new_n603_), .B2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT43), .ZN(new_n607_));
  OAI21_X1  g406(.A(KEYINPUT98), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n606_), .A2(KEYINPUT99), .A3(new_n607_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT98), .ZN(new_n610_));
  OAI211_X1 g409(.A(new_n610_), .B(KEYINPUT43), .C1(new_n380_), .C2(new_n596_), .ZN(new_n611_));
  OAI211_X1 g410(.A(new_n607_), .B(new_n536_), .C1(new_n376_), .C2(new_n379_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT99), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n608_), .A2(new_n609_), .A3(new_n611_), .A4(new_n614_), .ZN(new_n615_));
  NOR3_X1   g414(.A1(new_n503_), .A2(new_n417_), .A3(new_n548_), .ZN(new_n616_));
  AND3_X1   g415(.A1(new_n615_), .A2(KEYINPUT44), .A3(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(KEYINPUT44), .B1(new_n615_), .B2(new_n616_), .ZN(new_n618_));
  NOR3_X1   g417(.A1(new_n617_), .A2(new_n618_), .A3(new_n365_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n595_), .B1(new_n619_), .B2(new_n594_), .ZN(G1328gat));
  INV_X1    g419(.A(G36gat), .ZN(new_n621_));
  XOR2_X1   g420(.A(new_n371_), .B(KEYINPUT100), .Z(new_n622_));
  NAND3_X1  g421(.A1(new_n593_), .A2(new_n621_), .A3(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT45), .ZN(new_n624_));
  NOR3_X1   g423(.A1(new_n617_), .A2(new_n618_), .A3(new_n372_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n624_), .B1(new_n625_), .B2(new_n621_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT46), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  OAI211_X1 g427(.A(new_n624_), .B(KEYINPUT46), .C1(new_n625_), .C2(new_n621_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(G1329gat));
  AOI21_X1  g429(.A(G43gat), .B1(new_n593_), .B2(new_n237_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT101), .ZN(new_n632_));
  INV_X1    g431(.A(new_n618_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n615_), .A2(KEYINPUT44), .A3(new_n616_), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n633_), .A2(G43gat), .A3(new_n237_), .A4(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n632_), .A2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(KEYINPUT47), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT47), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n632_), .A2(new_n635_), .A3(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(G1330gat));
  NAND3_X1  g439(.A1(new_n633_), .A2(new_n377_), .A3(new_n634_), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n641_), .A2(KEYINPUT102), .A3(G50gat), .ZN(new_n642_));
  AOI21_X1  g441(.A(KEYINPUT102), .B1(new_n641_), .B2(G50gat), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n377_), .A2(new_n270_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT103), .ZN(new_n645_));
  OAI22_X1  g444(.A1(new_n642_), .A2(new_n643_), .B1(new_n592_), .B2(new_n645_), .ZN(G1331gat));
  INV_X1    g445(.A(new_n503_), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n380_), .A2(new_n416_), .A3(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(new_n550_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n461_), .B1(new_n649_), .B2(new_n365_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n648_), .A2(new_n558_), .ZN(new_n651_));
  OAI21_X1  g450(.A(G57gat), .B1(new_n365_), .B2(KEYINPUT104), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n652_), .B1(KEYINPUT104), .B2(G57gat), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n650_), .B1(new_n651_), .B2(new_n653_), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT105), .Z(G1332gat));
  INV_X1    g454(.A(new_n622_), .ZN(new_n656_));
  OAI21_X1  g455(.A(G64gat), .B1(new_n651_), .B2(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT48), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n622_), .A2(new_n462_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n658_), .B1(new_n649_), .B2(new_n659_), .ZN(G1333gat));
  OAI21_X1  g459(.A(G71gat), .B1(new_n651_), .B2(new_n580_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT49), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n580_), .A2(G71gat), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n662_), .B1(new_n649_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT106), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n664_), .B(new_n665_), .ZN(G1334gat));
  OAI21_X1  g465(.A(G78gat), .B1(new_n651_), .B2(new_n586_), .ZN(new_n667_));
  XOR2_X1   g466(.A(KEYINPUT107), .B(KEYINPUT50), .Z(new_n668_));
  OR2_X1    g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n668_), .ZN(new_n670_));
  OR3_X1    g469(.A1(new_n649_), .A2(G78gat), .A3(new_n586_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n669_), .A2(new_n670_), .A3(new_n671_), .ZN(G1335gat));
  NAND3_X1  g471(.A1(new_n648_), .A2(new_n553_), .A3(new_n591_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(new_n315_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT108), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n647_), .A2(new_n416_), .A3(new_n548_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n615_), .A2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT109), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n615_), .A2(KEYINPUT109), .A3(new_n676_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n365_), .A2(new_n315_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n675_), .B1(new_n681_), .B2(new_n682_), .ZN(G1336gat));
  NAND4_X1  g482(.A1(new_n648_), .A2(new_n334_), .A3(new_n371_), .A4(new_n591_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n656_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n684_), .B1(new_n685_), .B2(new_n334_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(KEYINPUT110), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT110), .ZN(new_n688_));
  OAI211_X1 g487(.A(new_n688_), .B(new_n684_), .C1(new_n685_), .C2(new_n334_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n689_), .ZN(G1337gat));
  NOR2_X1   g489(.A1(new_n677_), .A2(new_n580_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n691_), .A2(new_n428_), .ZN(new_n692_));
  AND4_X1   g491(.A1(new_n450_), .A2(new_n648_), .A3(new_n237_), .A4(new_n591_), .ZN(new_n693_));
  OAI22_X1  g492(.A1(new_n692_), .A2(new_n693_), .B1(KEYINPUT111), .B2(KEYINPUT51), .ZN(new_n694_));
  NAND2_X1  g493(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT112), .Z(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n694_), .A2(new_n697_), .ZN(new_n698_));
  OAI221_X1 g497(.A(new_n696_), .B1(KEYINPUT111), .B2(KEYINPUT51), .C1(new_n692_), .C2(new_n693_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1338gat));
  NAND4_X1  g499(.A1(new_n648_), .A2(new_n451_), .A3(new_n377_), .A4(new_n591_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n615_), .A2(new_n377_), .A3(new_n676_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT52), .ZN(new_n703_));
  AND3_X1   g502(.A1(new_n702_), .A2(new_n703_), .A3(G106gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n703_), .B1(new_n702_), .B2(G106gat), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n701_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g506(.A1(new_n486_), .A2(new_n489_), .A3(new_n498_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n416_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n484_), .B1(new_n481_), .B2(new_n485_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT55), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n486_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n479_), .A2(new_n480_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n714_), .A2(new_n487_), .A3(new_n485_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n715_), .A2(new_n712_), .A3(new_n483_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n713_), .A2(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(KEYINPUT56), .B1(new_n718_), .B2(new_n497_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT56), .ZN(new_n720_));
  AOI211_X1 g519(.A(new_n720_), .B(new_n498_), .C1(new_n713_), .C2(new_n717_), .ZN(new_n721_));
  OAI211_X1 g520(.A(KEYINPUT114), .B(new_n710_), .C1(new_n719_), .C2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n398_), .A2(new_n400_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n403_), .A2(new_n401_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n723_), .A2(new_n408_), .A3(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(KEYINPUT115), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT115), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n723_), .A2(new_n727_), .A3(new_n408_), .A4(new_n724_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n726_), .A2(new_n410_), .A3(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT116), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n726_), .A2(KEYINPUT116), .A3(new_n410_), .A4(new_n728_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n500_), .A2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n722_), .A2(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n712_), .B1(new_n715_), .B2(new_n483_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n715_), .A2(new_n483_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n497_), .B1(new_n739_), .B2(new_n716_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(new_n720_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n718_), .A2(KEYINPUT56), .A3(new_n497_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(KEYINPUT114), .B1(new_n743_), .B2(new_n710_), .ZN(new_n744_));
  OAI211_X1 g543(.A(KEYINPUT57), .B(new_n556_), .C1(new_n736_), .C2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT119), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n500_), .A2(new_n734_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n709_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n749_), .B2(KEYINPUT114), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT114), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n719_), .A2(new_n721_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n751_), .B1(new_n752_), .B2(new_n709_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n750_), .A2(new_n753_), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n754_), .A2(KEYINPUT119), .A3(KEYINPUT57), .A4(new_n556_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n747_), .A2(new_n755_), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n708_), .B(new_n733_), .C1(new_n719_), .C2(new_n721_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT58), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n596_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT118), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n743_), .A2(KEYINPUT58), .A3(new_n708_), .A4(new_n733_), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n759_), .A2(new_n760_), .A3(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n760_), .B1(new_n759_), .B2(new_n761_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n756_), .A2(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n556_), .B1(new_n736_), .B2(new_n744_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT57), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n766_), .A2(KEYINPUT117), .A3(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(KEYINPUT117), .B1(new_n766_), .B2(new_n767_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  OAI21_X1  g569(.A(KEYINPUT120), .B1(new_n765_), .B2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n766_), .A2(new_n767_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT117), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n766_), .A2(KEYINPUT117), .A3(new_n767_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT120), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n776_), .A2(new_n777_), .A3(new_n756_), .A4(new_n764_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n771_), .A2(new_n549_), .A3(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n550_), .A2(new_n647_), .A3(new_n417_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n780_), .A2(KEYINPUT54), .ZN(new_n781_));
  OR2_X1    g580(.A1(new_n781_), .A2(KEYINPUT113), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(KEYINPUT54), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(KEYINPUT113), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n782_), .A2(new_n783_), .A3(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n779_), .A2(new_n785_), .ZN(new_n786_));
  NOR4_X1   g585(.A1(new_n377_), .A2(new_n365_), .A3(new_n371_), .A4(new_n580_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT59), .ZN(new_n789_));
  AOI22_X1  g588(.A1(new_n766_), .A2(new_n767_), .B1(new_n761_), .B2(new_n759_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n548_), .B1(new_n756_), .B2(new_n790_), .ZN(new_n791_));
  OR2_X1    g590(.A1(new_n791_), .A2(KEYINPUT121), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(KEYINPUT121), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n792_), .A2(new_n785_), .A3(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT59), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n794_), .A2(new_n795_), .A3(new_n787_), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n789_), .A2(G113gat), .A3(new_n416_), .A4(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n788_), .ZN(new_n799_));
  AOI21_X1  g598(.A(G113gat), .B1(new_n799_), .B2(new_n416_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n798_), .A2(new_n800_), .ZN(G1340gat));
  INV_X1    g600(.A(G120gat), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n802_), .B1(new_n647_), .B2(KEYINPUT60), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n799_), .B(new_n803_), .C1(KEYINPUT60), .C2(new_n802_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n789_), .A2(new_n503_), .A3(new_n796_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n804_), .B1(new_n806_), .B2(new_n802_), .ZN(G1341gat));
  INV_X1    g606(.A(G127gat), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n808_), .B1(new_n788_), .B2(new_n549_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT122), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n789_), .A2(G127gat), .A3(new_n548_), .A4(new_n796_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT122), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n812_), .B(new_n808_), .C1(new_n788_), .C2(new_n549_), .ZN(new_n813_));
  AND3_X1   g612(.A1(new_n810_), .A2(new_n811_), .A3(new_n813_), .ZN(G1342gat));
  NAND4_X1  g613(.A1(new_n789_), .A2(G134gat), .A3(new_n536_), .A4(new_n796_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(G134gat), .B1(new_n799_), .B2(new_n557_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n816_), .A2(new_n817_), .ZN(G1343gat));
  AND3_X1   g617(.A1(new_n782_), .A2(new_n783_), .A3(new_n784_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n756_), .B(new_n764_), .C1(new_n769_), .C2(new_n768_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n548_), .B1(new_n820_), .B2(KEYINPUT120), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n819_), .B1(new_n821_), .B2(new_n778_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n656_), .A2(new_n377_), .A3(new_n580_), .ZN(new_n823_));
  NOR3_X1   g622(.A1(new_n822_), .A2(new_n365_), .A3(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n416_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n825_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n503_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g627(.A1(new_n824_), .A2(new_n548_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(KEYINPUT61), .B(G155gat), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n829_), .B(new_n830_), .ZN(G1346gat));
  AOI21_X1  g630(.A(G162gat), .B1(new_n824_), .B2(new_n557_), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n536_), .A2(G162gat), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n832_), .B1(new_n824_), .B2(new_n833_), .ZN(G1347gat));
  NAND2_X1  g633(.A1(new_n622_), .A2(new_n604_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n835_), .A2(new_n417_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n836_), .B(KEYINPUT123), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n837_), .A2(new_n377_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n211_), .B1(new_n794_), .B2(new_n838_), .ZN(new_n839_));
  XOR2_X1   g638(.A(new_n839_), .B(KEYINPUT62), .Z(new_n840_));
  AND4_X1   g639(.A1(new_n586_), .A2(new_n794_), .A3(new_n604_), .A4(new_n622_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n417_), .A2(new_n323_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n840_), .A2(new_n843_), .ZN(G1348gat));
  AOI21_X1  g643(.A(G176gat), .B1(new_n841_), .B2(new_n503_), .ZN(new_n845_));
  NOR3_X1   g644(.A1(new_n822_), .A2(new_n377_), .A3(new_n835_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n647_), .A2(new_n212_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n845_), .B1(new_n846_), .B2(new_n847_), .ZN(G1349gat));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n548_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT124), .ZN(new_n850_));
  AOI21_X1  g649(.A(G183gat), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n846_), .A2(KEYINPUT124), .A3(new_n548_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n549_), .A2(new_n221_), .ZN(new_n853_));
  AOI22_X1  g652(.A1(new_n851_), .A2(new_n852_), .B1(new_n841_), .B2(new_n853_), .ZN(G1350gat));
  NAND2_X1  g653(.A1(new_n841_), .A2(new_n536_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(G190gat), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n841_), .A2(new_n222_), .A3(new_n557_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(G1351gat));
  INV_X1    g657(.A(KEYINPUT126), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n377_), .A2(new_n365_), .A3(new_n580_), .ZN(new_n860_));
  XOR2_X1   g659(.A(new_n860_), .B(KEYINPUT125), .Z(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n622_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n859_), .B1(new_n822_), .B2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n862_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n786_), .A2(KEYINPUT126), .A3(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n863_), .A2(new_n865_), .ZN(new_n866_));
  AND3_X1   g665(.A1(new_n866_), .A2(G197gat), .A3(new_n416_), .ZN(new_n867_));
  AOI21_X1  g666(.A(G197gat), .B1(new_n866_), .B2(new_n416_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n867_), .A2(new_n868_), .ZN(G1352gat));
  AOI21_X1  g668(.A(new_n647_), .B1(new_n863_), .B2(new_n865_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(new_n286_), .ZN(G1353gat));
  INV_X1    g670(.A(KEYINPUT127), .ZN(new_n872_));
  XOR2_X1   g671(.A(KEYINPUT63), .B(G211gat), .Z(new_n873_));
  NAND4_X1  g672(.A1(new_n866_), .A2(new_n872_), .A3(new_n548_), .A4(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(KEYINPUT126), .B1(new_n786_), .B2(new_n864_), .ZN(new_n875_));
  AOI211_X1 g674(.A(new_n859_), .B(new_n862_), .C1(new_n779_), .C2(new_n785_), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n548_), .B(new_n873_), .C1(new_n875_), .C2(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(KEYINPUT127), .ZN(new_n878_));
  OR2_X1    g677(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n879_), .B1(new_n866_), .B2(new_n548_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n874_), .B1(new_n878_), .B2(new_n880_), .ZN(G1354gat));
  AOI21_X1  g680(.A(G218gat), .B1(new_n866_), .B2(new_n557_), .ZN(new_n882_));
  AND2_X1   g681(.A1(new_n536_), .A2(G218gat), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n882_), .B1(new_n866_), .B2(new_n883_), .ZN(G1355gat));
endmodule


