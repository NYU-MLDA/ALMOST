//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 1 1 1 1 0 1 0 0 1 0 1 0 1 0 1 0 0 1 0 1 0 1 0 0 0 1 0 1 1 0 0 0 1 1 1 1 1 0 1 1 0 0 1 0 1 1 1 1 0 1 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n701_, new_n702_, new_n703_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n750_, new_n751_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n854_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n860_, new_n862_, new_n863_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n899_,
    new_n900_, new_n902_, new_n903_, new_n904_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n921_, new_n922_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n930_;
  XOR2_X1   g000(.A(G169gat), .B(G176gat), .Z(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT24), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT25), .B(G183gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT26), .B(G190gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT24), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n203_), .A2(new_n206_), .A3(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n211_), .B1(G183gat), .B2(G190gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT77), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT77), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n215_), .A2(G183gat), .A3(G190gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n212_), .B1(new_n217_), .B2(new_n211_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n210_), .A2(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n220_));
  INV_X1    g019(.A(G169gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n220_), .B(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n214_), .A2(new_n216_), .A3(KEYINPUT23), .ZN(new_n223_));
  OR3_X1    g022(.A1(new_n213_), .A2(KEYINPUT78), .A3(KEYINPUT23), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT78), .B1(new_n213_), .B2(KEYINPUT23), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n223_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(G183gat), .A2(G190gat), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n222_), .B1(new_n226_), .B2(new_n228_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n219_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G71gat), .B(G99gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(KEYINPUT80), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G15gat), .B(G43gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n230_), .B(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G227gat), .A2(G233gat), .ZN(new_n236_));
  XOR2_X1   g035(.A(new_n236_), .B(KEYINPUT79), .Z(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT30), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n235_), .B(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT81), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G127gat), .B(G134gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G113gat), .B(G120gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n242_), .A2(new_n243_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n241_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  OR2_X1    g046(.A1(new_n242_), .A2(new_n243_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n248_), .A2(KEYINPUT81), .A3(new_n244_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT31), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n240_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT83), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n251_), .B(KEYINPUT82), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n253_), .B1(new_n239_), .B2(new_n254_), .ZN(new_n255_));
  AND2_X1   g054(.A1(new_n252_), .A2(new_n255_), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n239_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G1gat), .B(G29gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(G85gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT0), .B(G57gat), .ZN(new_n261_));
  XOR2_X1   g060(.A(new_n260_), .B(new_n261_), .Z(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G225gat), .A2(G233gat), .ZN(new_n264_));
  XOR2_X1   g063(.A(new_n264_), .B(KEYINPUT99), .Z(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  XOR2_X1   g065(.A(G155gat), .B(G162gat), .Z(new_n267_));
  INV_X1    g066(.A(KEYINPUT3), .ZN(new_n268_));
  INV_X1    g067(.A(G141gat), .ZN(new_n269_));
  INV_X1    g068(.A(G148gat), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n268_), .A2(new_n269_), .A3(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G141gat), .A2(G148gat), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT2), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  OAI21_X1  g073(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n271_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT84), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT84), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n279_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n267_), .B1(new_n276_), .B2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT85), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  OAI211_X1 g083(.A(KEYINPUT85), .B(new_n267_), .C1(new_n276_), .C2(new_n281_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n269_), .A2(new_n270_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n286_), .A2(new_n272_), .A3(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT1), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n288_), .B1(new_n267_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n284_), .A2(new_n285_), .A3(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(new_n250_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n293_), .A2(KEYINPUT4), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n290_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT98), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n248_), .A2(new_n244_), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n295_), .A2(new_n296_), .A3(new_n297_), .A4(new_n285_), .ZN(new_n298_));
  NAND4_X1  g097(.A1(new_n284_), .A2(new_n297_), .A3(new_n285_), .A4(new_n291_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT98), .ZN(new_n300_));
  AOI22_X1  g099(.A1(new_n295_), .A2(new_n285_), .B1(new_n247_), .B2(new_n249_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n298_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  AOI211_X1 g101(.A(new_n266_), .B(new_n294_), .C1(new_n302_), .C2(KEYINPUT4), .ZN(new_n303_));
  INV_X1    g102(.A(new_n264_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n293_), .A2(KEYINPUT98), .A3(new_n299_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n304_), .B1(new_n305_), .B2(new_n298_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n263_), .B1(new_n303_), .B2(new_n306_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n294_), .B1(new_n302_), .B2(KEYINPUT4), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(new_n265_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n306_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n309_), .A2(new_n310_), .A3(new_n262_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n307_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n258_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT94), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n292_), .A2(KEYINPUT29), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G228gat), .A2(G233gat), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n317_), .B(KEYINPUT87), .Z(new_n318_));
  XNOR2_X1  g117(.A(G197gat), .B(G204gat), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT21), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G211gat), .B(G218gat), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n321_), .A2(KEYINPUT88), .A3(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(KEYINPUT88), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n324_), .B1(new_n320_), .B2(new_n319_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n323_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n322_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n319_), .A2(new_n320_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT89), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT89), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n319_), .A2(new_n330_), .A3(new_n320_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n327_), .B1(new_n329_), .B2(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n326_), .A2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n316_), .A2(new_n318_), .A3(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n318_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT29), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n336_), .B1(new_n295_), .B2(new_n285_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n321_), .B(new_n324_), .ZN(new_n338_));
  AND2_X1   g137(.A1(new_n329_), .A2(new_n331_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n338_), .B1(new_n339_), .B2(new_n327_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n335_), .B1(new_n337_), .B2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G78gat), .B(G106gat), .ZN(new_n342_));
  XOR2_X1   g141(.A(new_n342_), .B(KEYINPUT90), .Z(new_n343_));
  NAND3_X1  g142(.A1(new_n334_), .A2(new_n341_), .A3(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT93), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n284_), .A2(new_n336_), .A3(new_n285_), .A4(new_n291_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT28), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT28), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n295_), .A2(new_n348_), .A3(new_n336_), .A4(new_n285_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G22gat), .B(G50gat), .ZN(new_n350_));
  XOR2_X1   g149(.A(new_n350_), .B(KEYINPUT86), .Z(new_n351_));
  NAND3_X1  g150(.A1(new_n347_), .A2(new_n349_), .A3(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n351_), .B1(new_n347_), .B2(new_n349_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n345_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT93), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n334_), .A2(new_n341_), .A3(new_n357_), .A4(new_n343_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n342_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n359_), .B1(new_n334_), .B2(new_n341_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n358_), .B1(new_n360_), .B2(KEYINPUT92), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n334_), .A2(new_n341_), .ZN(new_n362_));
  AND3_X1   g161(.A1(new_n362_), .A2(KEYINPUT92), .A3(new_n342_), .ZN(new_n363_));
  NOR3_X1   g162(.A1(new_n356_), .A2(new_n361_), .A3(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT91), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n344_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n343_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n362_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n366_), .A2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n362_), .A2(new_n365_), .A3(new_n367_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n355_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n315_), .B1(new_n364_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n361_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n347_), .A2(new_n349_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n351_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(new_n352_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n377_), .B1(KEYINPUT93), .B2(new_n344_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n363_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n373_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n343_), .B1(new_n334_), .B2(new_n341_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n381_), .B1(new_n365_), .B2(new_n344_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n370_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n377_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n380_), .A2(KEYINPUT94), .A3(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n372_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT27), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G226gat), .A2(G233gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  XOR2_X1   g190(.A(KEYINPUT96), .B(KEYINPUT24), .Z(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  AOI22_X1  g192(.A1(new_n393_), .A2(new_n202_), .B1(new_n204_), .B2(new_n205_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT97), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n392_), .A2(new_n207_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n226_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n395_), .B1(new_n226_), .B2(new_n396_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n394_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n218_), .A2(new_n227_), .ZN(new_n401_));
  OR2_X1    g200(.A1(new_n401_), .A2(new_n222_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n340_), .B1(new_n400_), .B2(new_n402_), .ZN(new_n403_));
  AND2_X1   g202(.A1(new_n226_), .A2(new_n228_), .ZN(new_n404_));
  OAI22_X1  g203(.A1(new_n404_), .A2(new_n222_), .B1(new_n218_), .B2(new_n210_), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT20), .B1(new_n405_), .B2(new_n333_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n391_), .B1(new_n403_), .B2(new_n406_), .ZN(new_n407_));
  XOR2_X1   g206(.A(G8gat), .B(G36gat), .Z(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT18), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G64gat), .B(G92gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n400_), .A2(new_n340_), .A3(new_n402_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT20), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n413_), .B1(new_n405_), .B2(new_n333_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n412_), .A2(new_n414_), .A3(new_n390_), .ZN(new_n415_));
  AND3_X1   g214(.A1(new_n407_), .A2(new_n411_), .A3(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n411_), .B1(new_n407_), .B2(new_n415_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n387_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n411_), .ZN(new_n419_));
  NOR3_X1   g218(.A1(new_n403_), .A2(new_n406_), .A3(new_n391_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n390_), .B1(new_n412_), .B2(new_n414_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n419_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n407_), .A2(new_n411_), .A3(new_n415_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n422_), .A2(KEYINPUT27), .A3(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n418_), .A2(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT102), .B1(new_n386_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n425_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT102), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n372_), .A2(new_n427_), .A3(new_n428_), .A4(new_n385_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n314_), .B1(new_n426_), .B2(new_n429_), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n418_), .A2(new_n424_), .A3(new_n307_), .A4(new_n311_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NOR3_X1   g231(.A1(new_n364_), .A2(new_n371_), .A3(new_n315_), .ZN(new_n433_));
  AOI21_X1  g232(.A(KEYINPUT94), .B1(new_n380_), .B2(new_n384_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n432_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n433_), .A2(new_n434_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n411_), .A2(KEYINPUT32), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n438_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n407_), .A2(new_n415_), .A3(new_n437_), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n312_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT100), .ZN(new_n443_));
  AOI211_X1 g242(.A(new_n304_), .B(new_n294_), .C1(new_n302_), .C2(KEYINPUT4), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n262_), .B1(new_n302_), .B2(new_n265_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n443_), .B1(new_n444_), .B2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n308_), .A2(new_n264_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n448_), .A2(KEYINPUT100), .A3(new_n445_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n407_), .A2(new_n415_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(new_n419_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(new_n423_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n450_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT33), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n311_), .A2(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n306_), .B1(new_n308_), .B2(new_n265_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n458_), .A2(KEYINPUT33), .A3(new_n262_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n442_), .B1(new_n455_), .B2(new_n460_), .ZN(new_n461_));
  AOI22_X1  g260(.A1(new_n435_), .A2(KEYINPUT101), .B1(new_n436_), .B2(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n431_), .B1(new_n372_), .B2(new_n385_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT101), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n462_), .A2(new_n465_), .ZN(new_n466_));
  OR2_X1    g265(.A1(new_n256_), .A2(new_n257_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n430_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G29gat), .B(G36gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G43gat), .B(G50gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT15), .ZN(new_n472_));
  XOR2_X1   g271(.A(G1gat), .B(G8gat), .Z(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G15gat), .B(G22gat), .ZN(new_n475_));
  INV_X1    g274(.A(G1gat), .ZN(new_n476_));
  INV_X1    g275(.A(G8gat), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT14), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n475_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT73), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n479_), .A2(KEYINPUT73), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n474_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n482_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n484_), .A2(new_n473_), .A3(new_n480_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n472_), .A2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n483_), .A2(new_n485_), .A3(new_n471_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G229gat), .A2(G233gat), .ZN(new_n489_));
  AND3_X1   g288(.A1(new_n487_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n471_), .B1(new_n483_), .B2(new_n485_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n489_), .B1(new_n492_), .B2(new_n488_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n490_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT76), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G113gat), .B(G141gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G169gat), .B(G197gat), .ZN(new_n497_));
  XOR2_X1   g296(.A(new_n496_), .B(new_n497_), .Z(new_n498_));
  OAI21_X1  g297(.A(new_n494_), .B1(new_n495_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n498_), .ZN(new_n500_));
  OAI211_X1 g299(.A(KEYINPUT76), .B(new_n500_), .C1(new_n490_), .C2(new_n493_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G99gat), .A2(G106gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(KEYINPUT6), .ZN(new_n505_));
  XOR2_X1   g304(.A(KEYINPUT10), .B(G99gat), .Z(new_n506_));
  INV_X1    g305(.A(G106gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G85gat), .A2(G92gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  AND2_X1   g310(.A1(new_n511_), .A2(KEYINPUT65), .ZN(new_n512_));
  NOR2_X1   g311(.A1(G85gat), .A2(G92gat), .ZN(new_n513_));
  INV_X1    g312(.A(new_n510_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n513_), .B1(new_n514_), .B2(KEYINPUT9), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n515_), .B1(new_n511_), .B2(KEYINPUT65), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n505_), .B(new_n508_), .C1(new_n512_), .C2(new_n516_), .ZN(new_n517_));
  OAI21_X1  g316(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n518_));
  OR2_X1    g317(.A1(new_n518_), .A2(KEYINPUT66), .ZN(new_n519_));
  OR3_X1    g318(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n518_), .A2(KEYINPUT66), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n505_), .A2(new_n519_), .A3(new_n520_), .A4(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT8), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n514_), .A2(new_n513_), .ZN(new_n524_));
  AND3_X1   g323(.A1(new_n522_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n523_), .B1(new_n522_), .B2(new_n524_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n517_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G57gat), .B(G64gat), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT11), .ZN(new_n529_));
  XOR2_X1   g328(.A(G71gat), .B(G78gat), .Z(new_n530_));
  NOR2_X1   g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  AND2_X1   g330(.A1(new_n529_), .A2(new_n530_), .ZN(new_n532_));
  OR2_X1    g331(.A1(new_n528_), .A2(KEYINPUT11), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n531_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  AND2_X1   g333(.A1(new_n527_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT12), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n527_), .A2(new_n534_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n534_), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n539_), .B(new_n517_), .C1(new_n526_), .C2(new_n525_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n538_), .A2(KEYINPUT12), .A3(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n537_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G230gat), .A2(G233gat), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n543_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n540_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n545_), .B1(new_n535_), .B2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n544_), .A2(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(G120gat), .B(G148gat), .Z(new_n549_));
  XNOR2_X1  g348(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G176gat), .B(G204gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  XOR2_X1   g352(.A(new_n553_), .B(KEYINPUT68), .Z(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n548_), .A2(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n544_), .A2(new_n547_), .A3(new_n553_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  XOR2_X1   g357(.A(KEYINPUT69), .B(KEYINPUT13), .Z(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT13), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n556_), .B(new_n557_), .C1(KEYINPUT69), .C2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n560_), .A2(new_n562_), .ZN(new_n563_));
  XOR2_X1   g362(.A(new_n563_), .B(KEYINPUT70), .Z(new_n564_));
  INV_X1    g363(.A(KEYINPUT71), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n527_), .A2(new_n472_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G232gat), .A2(G233gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT34), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT35), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  OAI211_X1 g370(.A(new_n517_), .B(new_n471_), .C1(new_n525_), .C2(new_n526_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n566_), .A2(new_n571_), .A3(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n569_), .A2(new_n570_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n574_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n566_), .A2(new_n576_), .A3(new_n571_), .A4(new_n572_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n565_), .B1(new_n575_), .B2(new_n577_), .ZN(new_n578_));
  XOR2_X1   g377(.A(G190gat), .B(G218gat), .Z(new_n579_));
  XNOR2_X1  g378(.A(G134gat), .B(G162gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(KEYINPUT36), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n583_), .B1(new_n575_), .B2(new_n577_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n582_), .A2(KEYINPUT36), .ZN(new_n585_));
  NOR3_X1   g384(.A1(new_n578_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n585_), .ZN(new_n587_));
  AOI221_X4 g386(.A(new_n565_), .B1(new_n587_), .B2(new_n583_), .C1(new_n575_), .C2(new_n577_), .ZN(new_n588_));
  OAI21_X1  g387(.A(KEYINPUT72), .B1(new_n586_), .B2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT37), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n584_), .A2(new_n585_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n578_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n588_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n596_), .A2(KEYINPUT72), .A3(KEYINPUT37), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n591_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(G231gat), .A2(G233gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT74), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n486_), .B(new_n601_), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n602_), .A2(new_n539_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n539_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  XOR2_X1   g404(.A(G127gat), .B(G155gat), .Z(new_n606_));
  XNOR2_X1  g405(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G183gat), .B(G211gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n610_), .B(KEYINPUT17), .Z(new_n611_));
  NAND2_X1  g410(.A1(new_n605_), .A2(new_n611_), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n603_), .A2(KEYINPUT17), .A3(new_n610_), .A4(new_n604_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n599_), .A2(new_n615_), .ZN(new_n616_));
  NOR4_X1   g415(.A1(new_n468_), .A2(new_n503_), .A3(new_n564_), .A4(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n617_), .A2(new_n476_), .A3(new_n312_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT38), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n468_), .A2(new_n596_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n563_), .A2(new_n502_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n622_), .A2(new_n614_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  OAI21_X1  g423(.A(G1gat), .B1(new_n624_), .B2(new_n313_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n618_), .A2(new_n619_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n620_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT103), .ZN(G1324gat));
  NAND3_X1  g427(.A1(new_n617_), .A2(new_n477_), .A3(new_n425_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT39), .ZN(new_n630_));
  INV_X1    g429(.A(new_n624_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(new_n425_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n630_), .B1(new_n632_), .B2(G8gat), .ZN(new_n633_));
  AOI211_X1 g432(.A(KEYINPUT39), .B(new_n477_), .C1(new_n631_), .C2(new_n425_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n629_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT40), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  OAI211_X1 g436(.A(KEYINPUT40), .B(new_n629_), .C1(new_n633_), .C2(new_n634_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(G1325gat));
  OAI21_X1  g438(.A(G15gat), .B1(new_n624_), .B2(new_n467_), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT41), .Z(new_n641_));
  INV_X1    g440(.A(G15gat), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n617_), .A2(new_n642_), .A3(new_n258_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n643_), .ZN(G1326gat));
  OAI21_X1  g443(.A(G22gat), .B1(new_n624_), .B2(new_n436_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT42), .ZN(new_n646_));
  INV_X1    g445(.A(G22gat), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n617_), .A2(new_n647_), .A3(new_n386_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(G1327gat));
  NOR2_X1   g448(.A1(new_n468_), .A2(new_n503_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n596_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n651_), .A2(new_n615_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n652_), .A2(new_n563_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n650_), .A2(new_n653_), .ZN(new_n654_));
  OR3_X1    g453(.A1(new_n654_), .A2(G29gat), .A3(new_n313_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT44), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT43), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n598_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n439_), .A2(new_n440_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n659_), .B1(new_n307_), .B2(new_n311_), .ZN(new_n660_));
  NOR4_X1   g459(.A1(new_n303_), .A2(new_n456_), .A3(new_n306_), .A4(new_n263_), .ZN(new_n661_));
  AOI21_X1  g460(.A(KEYINPUT33), .B1(new_n458_), .B2(new_n262_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n453_), .B1(new_n447_), .B2(new_n449_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n660_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  OAI22_X1  g464(.A1(new_n463_), .A2(new_n464_), .B1(new_n665_), .B2(new_n386_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n435_), .A2(KEYINPUT101), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n467_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n426_), .A2(new_n429_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n314_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n658_), .B1(new_n668_), .B2(new_n671_), .ZN(new_n672_));
  AND3_X1   g471(.A1(new_n591_), .A2(new_n597_), .A3(KEYINPUT104), .ZN(new_n673_));
  AOI21_X1  g472(.A(KEYINPUT104), .B1(new_n591_), .B2(new_n597_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n258_), .B1(new_n462_), .B2(new_n465_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n675_), .B1(new_n676_), .B2(new_n430_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n672_), .B1(new_n677_), .B2(KEYINPUT43), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n622_), .A2(new_n615_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n656_), .B1(new_n678_), .B2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n668_), .A2(new_n671_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n657_), .B1(new_n682_), .B2(new_n675_), .ZN(new_n683_));
  OAI211_X1 g482(.A(KEYINPUT44), .B(new_n679_), .C1(new_n683_), .C2(new_n672_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n681_), .A2(new_n312_), .A3(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT105), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n685_), .A2(new_n686_), .A3(G29gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n686_), .B1(new_n685_), .B2(G29gat), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n655_), .B1(new_n687_), .B2(new_n688_), .ZN(G1328gat));
  NOR2_X1   g488(.A1(new_n427_), .A2(G36gat), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n682_), .A2(new_n502_), .A3(new_n653_), .A4(new_n690_), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT45), .Z(new_n692_));
  NAND3_X1  g491(.A1(new_n681_), .A2(new_n425_), .A3(new_n684_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n692_), .B1(new_n693_), .B2(G36gat), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT46), .ZN(new_n695_));
  AND3_X1   g494(.A1(new_n694_), .A2(KEYINPUT106), .A3(new_n695_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n695_), .A2(KEYINPUT106), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n695_), .A2(KEYINPUT106), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n694_), .A2(new_n697_), .A3(new_n698_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n696_), .A2(new_n699_), .ZN(G1329gat));
  NAND4_X1  g499(.A1(new_n681_), .A2(G43gat), .A3(new_n258_), .A4(new_n684_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n654_), .A2(new_n467_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n701_), .B1(G43gat), .B2(new_n702_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g503(.A(new_n654_), .ZN(new_n705_));
  AOI21_X1  g504(.A(G50gat), .B1(new_n705_), .B2(new_n386_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n681_), .A2(new_n684_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n386_), .A2(G50gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n706_), .B1(new_n707_), .B2(new_n708_), .ZN(G1331gat));
  NAND2_X1  g508(.A1(new_n682_), .A2(new_n503_), .ZN(new_n710_));
  NOR3_X1   g509(.A1(new_n710_), .A2(new_n563_), .A3(new_n616_), .ZN(new_n711_));
  AOI21_X1  g510(.A(G57gat), .B1(new_n711_), .B2(new_n312_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT107), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n614_), .A2(new_n502_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n621_), .A2(new_n564_), .A3(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT108), .ZN(new_n716_));
  XOR2_X1   g515(.A(KEYINPUT109), .B(G57gat), .Z(new_n717_));
  NOR2_X1   g516(.A1(new_n313_), .A2(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n713_), .B1(new_n716_), .B2(new_n718_), .ZN(G1332gat));
  INV_X1    g518(.A(G64gat), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n711_), .A2(new_n720_), .A3(new_n425_), .ZN(new_n721_));
  XOR2_X1   g520(.A(KEYINPUT110), .B(KEYINPUT48), .Z(new_n722_));
  NAND2_X1  g521(.A1(new_n716_), .A2(new_n425_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n722_), .B1(new_n723_), .B2(G64gat), .ZN(new_n724_));
  INV_X1    g523(.A(new_n722_), .ZN(new_n725_));
  AOI211_X1 g524(.A(new_n720_), .B(new_n725_), .C1(new_n716_), .C2(new_n425_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n721_), .B1(new_n724_), .B2(new_n726_), .ZN(G1333gat));
  INV_X1    g526(.A(G71gat), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n711_), .A2(new_n728_), .A3(new_n258_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT49), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n716_), .A2(new_n258_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n731_), .B2(G71gat), .ZN(new_n732_));
  AOI211_X1 g531(.A(KEYINPUT49), .B(new_n728_), .C1(new_n716_), .C2(new_n258_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n729_), .B1(new_n732_), .B2(new_n733_), .ZN(G1334gat));
  INV_X1    g533(.A(G78gat), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n711_), .A2(new_n735_), .A3(new_n386_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT50), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n716_), .A2(new_n386_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n737_), .B1(new_n738_), .B2(G78gat), .ZN(new_n739_));
  AOI211_X1 g538(.A(KEYINPUT50), .B(new_n735_), .C1(new_n716_), .C2(new_n386_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n736_), .B1(new_n739_), .B2(new_n740_), .ZN(G1335gat));
  NOR3_X1   g540(.A1(new_n563_), .A2(new_n502_), .A3(new_n615_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n742_), .B1(new_n683_), .B2(new_n672_), .ZN(new_n743_));
  OAI21_X1  g542(.A(G85gat), .B1(new_n743_), .B2(new_n313_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n564_), .ZN(new_n745_));
  NOR4_X1   g544(.A1(new_n710_), .A2(new_n745_), .A3(new_n615_), .A4(new_n651_), .ZN(new_n746_));
  INV_X1    g545(.A(G85gat), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n746_), .A2(new_n747_), .A3(new_n312_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n744_), .A2(new_n748_), .ZN(G1336gat));
  INV_X1    g548(.A(G92gat), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n746_), .A2(new_n750_), .A3(new_n425_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n743_), .A2(new_n427_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n751_), .B1(new_n752_), .B2(new_n750_), .ZN(new_n753_));
  XOR2_X1   g552(.A(new_n753_), .B(KEYINPUT111), .Z(G1337gat));
  OAI21_X1  g553(.A(G99gat), .B1(new_n743_), .B2(new_n467_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n746_), .A2(new_n258_), .A3(new_n506_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI211_X1 g557(.A(new_n386_), .B(new_n742_), .C1(new_n683_), .C2(new_n672_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n759_), .A2(KEYINPUT112), .A3(G106gat), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(KEYINPUT112), .B1(new_n759_), .B2(G106gat), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT52), .ZN(new_n763_));
  NOR3_X1   g562(.A1(new_n761_), .A2(new_n762_), .A3(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n762_), .A2(new_n763_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n746_), .A2(new_n507_), .A3(new_n386_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(KEYINPUT53), .B1(new_n764_), .B2(new_n767_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n762_), .A2(new_n763_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(new_n760_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT53), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n770_), .A2(new_n771_), .A3(new_n765_), .A4(new_n766_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n768_), .A2(new_n772_), .ZN(G1339gat));
  NAND3_X1  g572(.A1(new_n537_), .A2(new_n545_), .A3(new_n541_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n544_), .A2(KEYINPUT55), .A3(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n545_), .B1(new_n537_), .B2(new_n541_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT55), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n554_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n775_), .A2(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n779_), .A2(KEYINPUT113), .A3(KEYINPUT56), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n502_), .A2(new_n557_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT113), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n784_), .B1(new_n775_), .B2(new_n778_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n785_), .A2(KEYINPUT56), .ZN(new_n786_));
  OAI21_X1  g585(.A(KEYINPUT114), .B1(new_n783_), .B2(new_n786_), .ZN(new_n787_));
  OR2_X1    g586(.A1(new_n785_), .A2(KEYINPUT56), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n781_), .B1(new_n785_), .B2(KEYINPUT56), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT114), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n788_), .A2(new_n789_), .A3(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n494_), .A2(new_n498_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT116), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT115), .ZN(new_n794_));
  INV_X1    g593(.A(new_n489_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n795_), .B1(new_n492_), .B2(new_n488_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n794_), .B1(new_n796_), .B2(new_n498_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n488_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n489_), .B1(new_n798_), .B2(new_n491_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n799_), .A2(KEYINPUT115), .A3(new_n500_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n797_), .A2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n487_), .A2(new_n488_), .A3(new_n795_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n793_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n801_), .A2(new_n802_), .A3(new_n793_), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n558_), .B(new_n792_), .C1(new_n803_), .C2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n787_), .A2(new_n791_), .A3(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT57), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(KEYINPUT117), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n806_), .A2(new_n651_), .A3(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(KEYINPUT56), .B1(new_n775_), .B2(new_n778_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n775_), .A2(KEYINPUT56), .A3(new_n778_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n811_), .A2(KEYINPUT118), .A3(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT118), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n810_), .A2(new_n814_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n557_), .B(new_n792_), .C1(new_n804_), .C2(new_n803_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n813_), .A2(new_n815_), .A3(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT58), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n813_), .A2(new_n817_), .A3(KEYINPUT58), .A4(new_n815_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n820_), .A2(new_n598_), .A3(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n809_), .A2(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n808_), .B1(new_n806_), .B2(new_n651_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n614_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n563_), .A2(new_n714_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n826_), .A2(new_n598_), .ZN(new_n827_));
  XOR2_X1   g626(.A(new_n827_), .B(KEYINPUT54), .Z(new_n828_));
  NAND2_X1  g627(.A1(new_n825_), .A2(new_n828_), .ZN(new_n829_));
  AOI211_X1 g628(.A(new_n313_), .B(new_n467_), .C1(new_n426_), .C2(new_n429_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  OR2_X1    g630(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  XOR2_X1   g632(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n829_), .A2(new_n830_), .A3(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n833_), .A2(new_n502_), .A3(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(G113gat), .ZN(new_n838_));
  OR2_X1    g637(.A1(new_n503_), .A2(G113gat), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n838_), .B1(new_n831_), .B2(new_n839_), .ZN(G1340gat));
  AND3_X1   g639(.A1(new_n833_), .A2(new_n564_), .A3(new_n836_), .ZN(new_n841_));
  INV_X1    g640(.A(G120gat), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n842_), .B1(new_n563_), .B2(KEYINPUT60), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n843_), .B1(KEYINPUT60), .B2(new_n842_), .ZN(new_n844_));
  OAI22_X1  g643(.A1(new_n841_), .A2(new_n842_), .B1(new_n831_), .B2(new_n844_), .ZN(G1341gat));
  NAND4_X1  g644(.A1(new_n833_), .A2(G127gat), .A3(new_n615_), .A4(new_n836_), .ZN(new_n846_));
  INV_X1    g645(.A(G127gat), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n847_), .B1(new_n831_), .B2(new_n614_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT120), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n846_), .A2(KEYINPUT120), .A3(new_n848_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(G1342gat));
  NAND3_X1  g652(.A1(new_n833_), .A2(new_n598_), .A3(new_n836_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(G134gat), .ZN(new_n855_));
  OR2_X1    g654(.A1(new_n651_), .A2(G134gat), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n855_), .B1(new_n831_), .B2(new_n856_), .ZN(G1343gat));
  NOR4_X1   g656(.A1(new_n258_), .A2(new_n436_), .A3(new_n313_), .A4(new_n425_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n829_), .A2(new_n858_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n859_), .A2(new_n503_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(new_n269_), .ZN(G1344gat));
  NOR2_X1   g660(.A1(new_n859_), .A2(new_n745_), .ZN(new_n862_));
  XOR2_X1   g661(.A(KEYINPUT121), .B(G148gat), .Z(new_n863_));
  XNOR2_X1  g662(.A(new_n862_), .B(new_n863_), .ZN(G1345gat));
  NOR2_X1   g663(.A1(new_n859_), .A2(new_n614_), .ZN(new_n865_));
  XOR2_X1   g664(.A(KEYINPUT61), .B(G155gat), .Z(new_n866_));
  XNOR2_X1  g665(.A(new_n865_), .B(new_n866_), .ZN(G1346gat));
  NOR2_X1   g666(.A1(new_n859_), .A2(new_n651_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n675_), .A2(G162gat), .ZN(new_n869_));
  OAI22_X1  g668(.A1(new_n868_), .A2(G162gat), .B1(new_n859_), .B2(new_n869_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(KEYINPUT122), .ZN(G1347gat));
  XOR2_X1   g670(.A(KEYINPUT22), .B(G169gat), .Z(new_n872_));
  NOR2_X1   g671(.A1(new_n503_), .A2(new_n872_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n314_), .A2(new_n386_), .A3(new_n427_), .ZN(new_n874_));
  AOI21_X1  g673(.A(KEYINPUT123), .B1(new_n829_), .B2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT123), .ZN(new_n876_));
  INV_X1    g675(.A(new_n874_), .ZN(new_n877_));
  AOI211_X1 g676(.A(new_n876_), .B(new_n877_), .C1(new_n825_), .C2(new_n828_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n873_), .B1(new_n875_), .B2(new_n878_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n877_), .B1(new_n825_), .B2(new_n828_), .ZN(new_n880_));
  AOI211_X1 g679(.A(KEYINPUT62), .B(new_n221_), .C1(new_n880_), .C2(new_n502_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT62), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n829_), .A2(new_n502_), .A3(new_n874_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n882_), .B1(new_n883_), .B2(G169gat), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n879_), .B1(new_n881_), .B2(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT124), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n879_), .B(KEYINPUT124), .C1(new_n881_), .C2(new_n884_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(G1348gat));
  INV_X1    g688(.A(G176gat), .ZN(new_n890_));
  OR2_X1    g689(.A1(new_n875_), .A2(new_n878_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n563_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  AND3_X1   g692(.A1(new_n880_), .A2(G176gat), .A3(new_n564_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT125), .ZN(new_n895_));
  OR2_X1    g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n895_), .ZN(new_n897_));
  AOI22_X1  g696(.A1(new_n890_), .A2(new_n893_), .B1(new_n896_), .B2(new_n897_), .ZN(G1349gat));
  AOI21_X1  g697(.A(G183gat), .B1(new_n880_), .B2(new_n615_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n614_), .A2(new_n204_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n899_), .B1(new_n891_), .B2(new_n900_), .ZN(G1350gat));
  NAND3_X1  g700(.A1(new_n891_), .A2(new_n205_), .A3(new_n596_), .ZN(new_n902_));
  AND2_X1   g701(.A1(new_n891_), .A2(new_n598_), .ZN(new_n903_));
  INV_X1    g702(.A(G190gat), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n902_), .B1(new_n903_), .B2(new_n904_), .ZN(G1351gat));
  NOR4_X1   g704(.A1(new_n258_), .A2(new_n436_), .A3(new_n312_), .A4(new_n427_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n906_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n907_), .B1(new_n825_), .B2(new_n828_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT126), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n908_), .B(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT127), .ZN(new_n911_));
  NAND4_X1  g710(.A1(new_n910_), .A2(new_n911_), .A3(G197gat), .A4(new_n502_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n909_), .B1(new_n829_), .B2(new_n906_), .ZN(new_n913_));
  AOI211_X1 g712(.A(KEYINPUT126), .B(new_n907_), .C1(new_n825_), .C2(new_n828_), .ZN(new_n914_));
  OAI211_X1 g713(.A(G197gat), .B(new_n502_), .C1(new_n913_), .C2(new_n914_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(KEYINPUT127), .ZN(new_n916_));
  INV_X1    g715(.A(G197gat), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n913_), .A2(new_n914_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n918_), .B2(new_n503_), .ZN(new_n919_));
  AND3_X1   g718(.A1(new_n912_), .A2(new_n916_), .A3(new_n919_), .ZN(G1352gat));
  OR3_X1    g719(.A1(new_n918_), .A2(G204gat), .A3(new_n745_), .ZN(new_n921_));
  OAI21_X1  g720(.A(G204gat), .B1(new_n918_), .B2(new_n745_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(G1353gat));
  OR2_X1    g722(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n924_), .B1(new_n910_), .B2(new_n615_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n918_), .A2(new_n614_), .ZN(new_n926_));
  XOR2_X1   g725(.A(KEYINPUT63), .B(G211gat), .Z(new_n927_));
  AOI21_X1  g726(.A(new_n925_), .B1(new_n926_), .B2(new_n927_), .ZN(G1354gat));
  OR3_X1    g727(.A1(new_n918_), .A2(G218gat), .A3(new_n651_), .ZN(new_n929_));
  OAI21_X1  g728(.A(G218gat), .B1(new_n918_), .B2(new_n599_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n929_), .A2(new_n930_), .ZN(G1355gat));
endmodule


