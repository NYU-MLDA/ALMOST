//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 0 0 0 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 0 1 0 1 0 1 0 0 0 1 0 1 0 0 1 0 0 0 0 0 1 1 0 1 1 1 0 0 1 1 0 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n741_, new_n742_, new_n743_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n851_, new_n852_, new_n854_, new_n855_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n862_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n886_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n909_, new_n910_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_;
  INV_X1    g000(.A(KEYINPUT105), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT37), .ZN(new_n203_));
  XOR2_X1   g002(.A(KEYINPUT10), .B(G99gat), .Z(new_n204_));
  INV_X1    g003(.A(G106gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT6), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT6), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n208_), .A2(G99gat), .A3(G106gat), .ZN(new_n209_));
  AOI22_X1  g008(.A1(new_n204_), .A2(new_n205_), .B1(new_n207_), .B2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G85gat), .ZN(new_n211_));
  INV_X1    g010(.A(G92gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  AND2_X1   g012(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n214_));
  NOR2_X1   g013(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n213_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G85gat), .A2(G92gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT65), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND4_X1  g019(.A1(KEYINPUT65), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n221_));
  AOI22_X1  g020(.A1(new_n216_), .A2(new_n217_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n210_), .B1(new_n222_), .B2(KEYINPUT66), .ZN(new_n223_));
  INV_X1    g022(.A(new_n217_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n224_), .B1(new_n225_), .B2(new_n213_), .ZN(new_n226_));
  AND2_X1   g025(.A1(new_n220_), .A2(new_n221_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT66), .ZN(new_n228_));
  NOR3_X1   g027(.A1(new_n226_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n213_), .A2(new_n217_), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  NOR3_X1   g031(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n207_), .A2(new_n209_), .ZN(new_n235_));
  AOI211_X1 g034(.A(KEYINPUT8), .B(new_n230_), .C1(new_n234_), .C2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT8), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT7), .ZN(new_n238_));
  INV_X1    g037(.A(G99gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n238_), .A2(new_n239_), .A3(new_n205_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n208_), .B1(G99gat), .B2(G106gat), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n206_), .A2(KEYINPUT6), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n231_), .B(new_n240_), .C1(new_n241_), .C2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n230_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n237_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  OAI22_X1  g044(.A1(new_n223_), .A2(new_n229_), .B1(new_n236_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n243_), .A2(new_n244_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT8), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n243_), .A2(new_n237_), .A3(new_n244_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n222_), .A2(KEYINPUT66), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n228_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n253_), .A2(new_n254_), .A3(new_n210_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n252_), .A2(new_n255_), .A3(KEYINPUT67), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G29gat), .B(G36gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G43gat), .B(G50gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n248_), .A2(new_n256_), .A3(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G232gat), .A2(G233gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT34), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n262_), .A2(KEYINPUT35), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n259_), .B(KEYINPUT15), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n263_), .B1(new_n264_), .B2(new_n246_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n262_), .A2(KEYINPUT35), .ZN(new_n266_));
  XOR2_X1   g065(.A(new_n266_), .B(KEYINPUT71), .Z(new_n267_));
  NAND4_X1  g066(.A1(new_n260_), .A2(KEYINPUT72), .A3(new_n265_), .A4(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n260_), .A2(new_n265_), .A3(new_n267_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT72), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n266_), .B1(new_n260_), .B2(new_n265_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n268_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G190gat), .B(G218gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G134gat), .B(G162gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n276_), .A2(KEYINPUT36), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n273_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT73), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n273_), .A2(KEYINPUT73), .A3(new_n277_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(new_n276_), .B(KEYINPUT36), .Z(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT74), .ZN(new_n284_));
  OR2_X1    g083(.A1(new_n273_), .A2(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n203_), .B1(new_n282_), .B2(new_n285_), .ZN(new_n286_));
  OAI211_X1 g085(.A(new_n268_), .B(new_n283_), .C1(new_n271_), .C2(new_n272_), .ZN(new_n287_));
  AND3_X1   g086(.A1(new_n273_), .A2(KEYINPUT73), .A3(new_n277_), .ZN(new_n288_));
  AOI21_X1  g087(.A(KEYINPUT73), .B1(new_n273_), .B2(new_n277_), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n203_), .B(new_n287_), .C1(new_n288_), .C2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT75), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n282_), .A2(KEYINPUT75), .A3(new_n203_), .A4(new_n287_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n286_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT76), .B(G15gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(G22gat), .ZN(new_n296_));
  INV_X1    g095(.A(G1gat), .ZN(new_n297_));
  INV_X1    g096(.A(G8gat), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT14), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n296_), .A2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G1gat), .B(G8gat), .ZN(new_n301_));
  OR2_X1    g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n301_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G231gat), .A2(G233gat), .ZN(new_n305_));
  XOR2_X1   g104(.A(new_n304_), .B(new_n305_), .Z(new_n306_));
  XNOR2_X1  g105(.A(G57gat), .B(G64gat), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT68), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n307_), .A2(new_n308_), .ZN(new_n311_));
  OAI21_X1  g110(.A(KEYINPUT11), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G71gat), .B(G78gat), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n307_), .A2(new_n308_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT11), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n315_), .A2(new_n316_), .A3(new_n309_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n312_), .A2(new_n314_), .A3(new_n317_), .ZN(new_n318_));
  OAI211_X1 g117(.A(KEYINPUT11), .B(new_n313_), .C1(new_n310_), .C2(new_n311_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  OR2_X1    g119(.A1(new_n306_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n306_), .A2(new_n320_), .ZN(new_n322_));
  XOR2_X1   g121(.A(G127gat), .B(G155gat), .Z(new_n323_));
  XNOR2_X1  g122(.A(G183gat), .B(G211gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  XOR2_X1   g126(.A(new_n327_), .B(KEYINPUT17), .Z(new_n328_));
  NAND3_X1  g127(.A1(new_n321_), .A2(new_n322_), .A3(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT80), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT80), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n321_), .A2(new_n331_), .A3(new_n322_), .A4(new_n328_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n321_), .A2(new_n322_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT77), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n321_), .A2(KEYINPUT77), .A3(new_n322_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n327_), .A2(KEYINPUT17), .ZN(new_n338_));
  XOR2_X1   g137(.A(new_n338_), .B(KEYINPUT79), .Z(new_n339_));
  NAND3_X1  g138(.A1(new_n336_), .A2(new_n337_), .A3(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n333_), .A2(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n294_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT81), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT27), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT98), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G226gat), .A2(G233gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT19), .ZN(new_n347_));
  XOR2_X1   g146(.A(new_n347_), .B(KEYINPUT93), .Z(new_n348_));
  NAND2_X1  g147(.A1(G183gat), .A2(G190gat), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT23), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n352_));
  OAI211_X1 g151(.A(new_n351_), .B(new_n352_), .C1(G183gat), .C2(G190gat), .ZN(new_n353_));
  OR2_X1    g152(.A1(new_n353_), .A2(KEYINPUT95), .ZN(new_n354_));
  NOR2_X1   g153(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n355_));
  INV_X1    g154(.A(G169gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n357_), .B1(new_n353_), .B2(KEYINPUT95), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT26), .B(G190gat), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT25), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(G183gat), .ZN(new_n361_));
  INV_X1    g160(.A(G183gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT25), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n361_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT94), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(KEYINPUT94), .B1(new_n361_), .B2(new_n363_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n359_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  OR2_X1    g167(.A1(G169gat), .A2(G176gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G169gat), .A2(G176gat), .ZN(new_n370_));
  AND3_X1   g169(.A1(new_n369_), .A2(KEYINPUT24), .A3(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n351_), .A2(new_n352_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n369_), .A2(KEYINPUT24), .ZN(new_n373_));
  NOR3_X1   g172(.A1(new_n371_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n374_));
  AOI22_X1  g173(.A1(new_n354_), .A2(new_n358_), .B1(new_n368_), .B2(new_n374_), .ZN(new_n375_));
  XOR2_X1   g174(.A(G211gat), .B(G218gat), .Z(new_n376_));
  INV_X1    g175(.A(KEYINPUT21), .ZN(new_n377_));
  OR2_X1    g176(.A1(G197gat), .A2(G204gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G197gat), .A2(G204gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n376_), .B1(new_n377_), .B2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n380_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(KEYINPUT21), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n381_), .A2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n382_), .A2(new_n376_), .A3(KEYINPUT21), .ZN(new_n385_));
  AND2_X1   g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(KEYINPUT20), .B1(new_n375_), .B2(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(KEYINPUT84), .B1(new_n360_), .B2(G183gat), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT84), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n389_), .A2(new_n362_), .A3(KEYINPUT25), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT85), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n392_), .B1(new_n362_), .B2(KEYINPUT25), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n360_), .A2(KEYINPUT85), .A3(G183gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n391_), .A2(new_n395_), .A3(new_n359_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT86), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n391_), .A2(new_n395_), .A3(KEYINPUT86), .A4(new_n359_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n398_), .A2(new_n374_), .A3(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n357_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(new_n353_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n384_), .A2(new_n385_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n348_), .B1(new_n387_), .B2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT20), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n407_), .B1(new_n375_), .B2(new_n386_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n347_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n403_), .A2(new_n404_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n408_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n406_), .A2(new_n411_), .ZN(new_n412_));
  XOR2_X1   g211(.A(G8gat), .B(G36gat), .Z(new_n413_));
  XNOR2_X1  g212(.A(G64gat), .B(G92gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n415_), .B(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n345_), .B1(new_n412_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n417_), .ZN(new_n419_));
  AOI211_X1 g218(.A(KEYINPUT98), .B(new_n419_), .C1(new_n406_), .C2(new_n411_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n418_), .A2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n406_), .A2(new_n419_), .A3(new_n411_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT97), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT97), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n406_), .A2(new_n424_), .A3(new_n411_), .A4(new_n419_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n423_), .A2(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n344_), .B1(new_n421_), .B2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(G155gat), .ZN(new_n428_));
  INV_X1    g227(.A(G162gat), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n428_), .A2(new_n429_), .A3(KEYINPUT89), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT89), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n431_), .B1(G155gat), .B2(G162gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n430_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G155gat), .A2(G162gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT90), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT90), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n436_), .A2(G155gat), .A3(G162gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n433_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT91), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n433_), .A2(new_n438_), .A3(KEYINPUT91), .ZN(new_n442_));
  NOR2_X1   g241(.A1(G141gat), .A2(G148gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT3), .ZN(new_n444_));
  NAND2_X1  g243(.A1(G141gat), .A2(G148gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n445_), .B(KEYINPUT2), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n444_), .A2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n441_), .A2(new_n442_), .A3(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n443_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n433_), .B1(new_n438_), .B2(KEYINPUT1), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT1), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n451_), .B1(new_n435_), .B2(new_n437_), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n449_), .B(new_n445_), .C1(new_n450_), .C2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n448_), .A2(new_n453_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n454_), .A2(KEYINPUT29), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT28), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT28), .B1(new_n454_), .B2(KEYINPUT29), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n386_), .B1(new_n454_), .B2(KEYINPUT29), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  AND2_X1   g260(.A1(KEYINPUT92), .A2(G233gat), .ZN(new_n462_));
  NOR2_X1   g261(.A1(KEYINPUT92), .A2(G233gat), .ZN(new_n463_));
  OAI21_X1  g262(.A(G228gat), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(G78gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(new_n205_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G22gat), .B(G50gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n461_), .B(new_n469_), .ZN(new_n470_));
  NOR3_X1   g269(.A1(new_n387_), .A2(new_n405_), .A3(new_n348_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n409_), .B1(new_n408_), .B2(new_n410_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  OAI211_X1 g272(.A(KEYINPUT27), .B(new_n422_), .C1(new_n473_), .C2(new_n419_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n427_), .A2(new_n470_), .A3(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT102), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT102), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n427_), .A2(new_n470_), .A3(new_n477_), .A4(new_n474_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n476_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G227gat), .A2(G233gat), .ZN(new_n480_));
  INV_X1    g279(.A(G71gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n400_), .A2(KEYINPUT30), .A3(new_n402_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(KEYINPUT30), .B1(new_n400_), .B2(new_n402_), .ZN(new_n486_));
  OAI21_X1  g285(.A(G99gat), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT30), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n403_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n489_), .A2(new_n239_), .A3(new_n484_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G15gat), .B(G43gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT87), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n487_), .A2(new_n490_), .A3(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n493_), .B1(new_n487_), .B2(new_n490_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n483_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n487_), .A2(new_n490_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(new_n492_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n487_), .A2(new_n490_), .A3(new_n493_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n498_), .A2(new_n482_), .A3(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT88), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n496_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT31), .ZN(new_n503_));
  XOR2_X1   g302(.A(G127gat), .B(G134gat), .Z(new_n504_));
  XOR2_X1   g303(.A(G113gat), .B(G120gat), .Z(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT31), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n496_), .A2(new_n500_), .A3(new_n501_), .A4(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n503_), .A2(new_n507_), .A3(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n507_), .B1(new_n503_), .B2(new_n509_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT4), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n454_), .A2(new_n514_), .A3(new_n507_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G225gat), .A2(G233gat), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT100), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n454_), .A2(new_n507_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT99), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n448_), .A2(new_n453_), .A3(new_n506_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n521_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n454_), .A2(KEYINPUT99), .A3(new_n507_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n520_), .B1(new_n526_), .B2(KEYINPUT4), .ZN(new_n527_));
  AOI211_X1 g326(.A(KEYINPUT100), .B(new_n514_), .C1(new_n524_), .C2(new_n525_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n519_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n526_), .A2(new_n516_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  XOR2_X1   g330(.A(G1gat), .B(G29gat), .Z(new_n532_));
  XNOR2_X1  g331(.A(KEYINPUT101), .B(KEYINPUT0), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G57gat), .B(G85gat), .ZN(new_n535_));
  XOR2_X1   g334(.A(new_n534_), .B(new_n535_), .Z(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n531_), .A2(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n529_), .A2(new_n530_), .A3(new_n536_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n479_), .A2(new_n513_), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n512_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(new_n510_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n470_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT33), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n539_), .A2(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n421_), .A2(new_n426_), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n529_), .A2(KEYINPUT33), .A3(new_n530_), .A4(new_n536_), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n516_), .B(new_n515_), .C1(new_n527_), .C2(new_n528_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n536_), .B1(new_n526_), .B2(new_n517_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n547_), .A2(new_n548_), .A3(new_n549_), .A4(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n419_), .A2(KEYINPUT32), .ZN(new_n554_));
  MUX2_X1   g353(.A(new_n473_), .B(new_n412_), .S(new_n554_), .Z(new_n555_));
  INV_X1    g354(.A(new_n539_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n536_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n555_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n545_), .B1(new_n553_), .B2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n427_), .A2(new_n474_), .ZN(new_n560_));
  NOR3_X1   g359(.A1(new_n560_), .A2(new_n540_), .A3(new_n470_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n544_), .B1(new_n559_), .B2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n542_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G230gat), .A2(G233gat), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n248_), .A2(new_n320_), .A3(new_n256_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n320_), .B1(new_n248_), .B2(new_n256_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n565_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n318_), .A2(new_n319_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n570_), .A2(KEYINPUT12), .A3(new_n246_), .ZN(new_n571_));
  OAI211_X1 g370(.A(new_n566_), .B(new_n571_), .C1(new_n568_), .C2(KEYINPUT12), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n569_), .B1(new_n572_), .B2(new_n565_), .ZN(new_n573_));
  XOR2_X1   g372(.A(G120gat), .B(G148gat), .Z(new_n574_));
  XNOR2_X1  g373(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G176gat), .B(G204gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n573_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT70), .ZN(new_n580_));
  INV_X1    g379(.A(new_n578_), .ZN(new_n581_));
  OAI211_X1 g380(.A(new_n569_), .B(new_n581_), .C1(new_n572_), .C2(new_n565_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n579_), .A2(new_n580_), .A3(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n573_), .A2(KEYINPUT70), .A3(new_n578_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT13), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G229gat), .A2(G233gat), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n302_), .A2(new_n303_), .A3(new_n259_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n259_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n590_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n304_), .A2(new_n264_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n595_), .A2(new_n591_), .A3(new_n589_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n594_), .A2(new_n596_), .ZN(new_n597_));
  XOR2_X1   g396(.A(G113gat), .B(G141gat), .Z(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT82), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G169gat), .B(G197gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n597_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n594_), .A2(new_n596_), .A3(new_n601_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  OR2_X1    g405(.A1(new_n606_), .A2(KEYINPUT83), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(KEYINPUT83), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n588_), .A2(new_n610_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n563_), .A2(new_n611_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n343_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT103), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n541_), .A2(G1gat), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n613_), .A2(new_n614_), .A3(KEYINPUT38), .A4(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n343_), .A2(new_n612_), .A3(new_n615_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT38), .ZN(new_n618_));
  OAI21_X1  g417(.A(KEYINPUT103), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n616_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n282_), .A2(new_n287_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n622_), .B1(new_n542_), .B2(new_n562_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n587_), .A2(new_n605_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n624_), .A2(new_n341_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n623_), .A2(new_n540_), .A3(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(G1gat), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT104), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n617_), .A2(new_n618_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n202_), .B1(new_n620_), .B2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n616_), .A2(new_n619_), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n633_), .A2(KEYINPUT105), .A3(new_n630_), .A4(new_n629_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(G1324gat));
  NAND3_X1  g434(.A1(new_n613_), .A2(new_n298_), .A3(new_n560_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT106), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n623_), .A2(new_n625_), .A3(new_n637_), .A4(new_n560_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n638_), .A2(G8gat), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT39), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n623_), .A2(new_n560_), .A3(new_n625_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(KEYINPUT106), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n639_), .A2(new_n640_), .A3(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n640_), .B1(new_n639_), .B2(new_n642_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n636_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT40), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  OAI211_X1 g446(.A(KEYINPUT40), .B(new_n636_), .C1(new_n643_), .C2(new_n644_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(G1325gat));
  AND2_X1   g448(.A1(new_n623_), .A2(new_n625_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(new_n513_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(G15gat), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n652_), .A2(KEYINPUT41), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(KEYINPUT41), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT107), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(G15gat), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n613_), .A2(new_n658_), .A3(new_n513_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT108), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n653_), .A2(KEYINPUT107), .A3(new_n654_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n657_), .A2(new_n661_), .A3(new_n662_), .ZN(G1326gat));
  INV_X1    g462(.A(G22gat), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n664_), .B1(new_n650_), .B2(new_n545_), .ZN(new_n665_));
  XOR2_X1   g464(.A(new_n665_), .B(KEYINPUT42), .Z(new_n666_));
  NAND3_X1  g465(.A1(new_n613_), .A2(new_n664_), .A3(new_n545_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1327gat));
  INV_X1    g467(.A(new_n341_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n624_), .A2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n292_), .A2(new_n293_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n286_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  AOI211_X1 g472(.A(KEYINPUT43), .B(new_n673_), .C1(new_n562_), .C2(new_n542_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT43), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n675_), .B1(new_n563_), .B2(new_n294_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n670_), .B1(new_n674_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  OAI211_X1 g478(.A(KEYINPUT44), .B(new_n670_), .C1(new_n674_), .C2(new_n676_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n679_), .A2(new_n540_), .A3(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(G29gat), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n622_), .A2(new_n341_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n612_), .A2(new_n684_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n541_), .A2(G29gat), .ZN(new_n686_));
  XOR2_X1   g485(.A(new_n686_), .B(KEYINPUT109), .Z(new_n687_));
  OAI21_X1  g486(.A(new_n682_), .B1(new_n685_), .B2(new_n687_), .ZN(G1328gat));
  INV_X1    g487(.A(new_n560_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n689_), .A2(G36gat), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n563_), .A2(new_n611_), .A3(new_n684_), .A4(new_n690_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n691_), .A2(KEYINPUT45), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n691_), .A2(KEYINPUT45), .ZN(new_n693_));
  OAI22_X1  g492(.A1(new_n692_), .A2(new_n693_), .B1(KEYINPUT110), .B2(KEYINPUT46), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n679_), .A2(new_n560_), .A3(new_n680_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n695_), .B2(G36gat), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT110), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT46), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n696_), .A2(new_n700_), .ZN(new_n701_));
  AOI211_X1 g500(.A(new_n699_), .B(new_n694_), .C1(new_n695_), .C2(G36gat), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n701_), .A2(new_n702_), .ZN(G1329gat));
  NAND3_X1  g502(.A1(new_n612_), .A2(new_n513_), .A3(new_n684_), .ZN(new_n704_));
  INV_X1    g503(.A(G43gat), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT111), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n706_), .B(new_n707_), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n679_), .A2(G43gat), .A3(new_n513_), .A4(new_n680_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(KEYINPUT47), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT47), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n708_), .A2(new_n709_), .A3(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(G1330gat));
  NAND3_X1  g513(.A1(new_n679_), .A2(new_n545_), .A3(new_n680_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(G50gat), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n470_), .A2(G50gat), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT112), .Z(new_n718_));
  OAI21_X1  g517(.A(new_n716_), .B1(new_n685_), .B2(new_n718_), .ZN(G1331gat));
  AOI211_X1 g518(.A(new_n587_), .B(new_n605_), .C1(new_n542_), .C2(new_n562_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n343_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(G57gat), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n721_), .A2(new_n722_), .A3(new_n540_), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n587_), .A2(new_n341_), .A3(new_n609_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n623_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  OAI21_X1  g525(.A(G57gat), .B1(new_n726_), .B2(new_n541_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n723_), .A2(new_n727_), .ZN(G1332gat));
  INV_X1    g527(.A(G64gat), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n721_), .A2(new_n729_), .A3(new_n560_), .ZN(new_n730_));
  AOI211_X1 g529(.A(KEYINPUT48), .B(new_n729_), .C1(new_n725_), .C2(new_n560_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT48), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n725_), .A2(new_n560_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n733_), .B2(G64gat), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n730_), .B1(new_n731_), .B2(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT113), .ZN(G1333gat));
  AOI21_X1  g535(.A(new_n481_), .B1(new_n725_), .B2(new_n513_), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n737_), .B(KEYINPUT49), .Z(new_n738_));
  NAND3_X1  g537(.A1(new_n721_), .A2(new_n481_), .A3(new_n513_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(G1334gat));
  AOI21_X1  g539(.A(new_n465_), .B1(new_n725_), .B2(new_n545_), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n741_), .B(KEYINPUT50), .Z(new_n742_));
  NAND3_X1  g541(.A1(new_n721_), .A2(new_n465_), .A3(new_n545_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(G1335gat));
  NOR3_X1   g543(.A1(new_n587_), .A2(new_n669_), .A3(new_n605_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT114), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n746_), .B1(new_n674_), .B2(new_n676_), .ZN(new_n747_));
  OAI21_X1  g546(.A(G85gat), .B1(new_n747_), .B2(new_n541_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n720_), .A2(new_n684_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n749_), .A2(new_n211_), .A3(new_n540_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n750_), .ZN(G1336gat));
  OAI21_X1  g550(.A(G92gat), .B1(new_n747_), .B2(new_n689_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n749_), .A2(new_n212_), .A3(new_n560_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(G1337gat));
  OAI21_X1  g553(.A(G99gat), .B1(new_n747_), .B2(new_n544_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n749_), .A2(new_n204_), .A3(new_n513_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g557(.A1(new_n749_), .A2(new_n205_), .A3(new_n545_), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n746_), .B(new_n545_), .C1(new_n674_), .C2(new_n676_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT52), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n760_), .A2(new_n761_), .A3(G106gat), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n760_), .B2(G106gat), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n759_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(KEYINPUT53), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT53), .ZN(new_n766_));
  OAI211_X1 g565(.A(new_n766_), .B(new_n759_), .C1(new_n762_), .C2(new_n763_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n765_), .A2(new_n767_), .ZN(G1339gat));
  AND2_X1   g567(.A1(new_n566_), .A2(new_n571_), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n252_), .A2(new_n255_), .A3(KEYINPUT67), .ZN(new_n770_));
  AOI21_X1  g569(.A(KEYINPUT67), .B1(new_n252_), .B2(new_n255_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n570_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT12), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n769_), .A2(new_n774_), .A3(KEYINPUT55), .A4(new_n564_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT115), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n248_), .A2(new_n256_), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT12), .B1(new_n777_), .B2(new_n570_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n566_), .A2(new_n571_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT115), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n780_), .A2(new_n781_), .A3(KEYINPUT55), .A4(new_n564_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n572_), .A2(new_n565_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT55), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n784_), .B1(new_n572_), .B2(new_n565_), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n776_), .A2(new_n782_), .A3(new_n783_), .A4(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(new_n578_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(KEYINPUT56), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT56), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n786_), .A2(new_n789_), .A3(new_n578_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n595_), .A2(new_n591_), .A3(new_n590_), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n791_), .A2(new_n602_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n589_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n793_));
  AOI21_X1  g592(.A(KEYINPUT117), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n793_), .A2(new_n791_), .A3(KEYINPUT117), .A4(new_n602_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n604_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n794_), .A2(new_n796_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n797_), .A2(new_n582_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n788_), .A2(new_n790_), .A3(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT58), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n788_), .A2(KEYINPUT58), .A3(new_n790_), .A4(new_n798_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n294_), .A2(new_n801_), .A3(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT57), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n583_), .A2(new_n584_), .A3(new_n797_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n605_), .A2(new_n582_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(KEYINPUT116), .A2(KEYINPUT56), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n806_), .B1(new_n787_), .B2(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n786_), .A2(new_n578_), .A3(new_n807_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n805_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n804_), .B1(new_n811_), .B2(new_n622_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n810_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n807_), .B1(new_n786_), .B2(new_n578_), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n813_), .A2(new_n814_), .A3(new_n806_), .ZN(new_n815_));
  OAI211_X1 g614(.A(KEYINPUT57), .B(new_n621_), .C1(new_n815_), .C2(new_n805_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n803_), .A2(new_n812_), .A3(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n341_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n341_), .A2(new_n609_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n587_), .A2(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(KEYINPUT54), .B1(new_n820_), .B2(new_n294_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n673_), .A2(new_n822_), .A3(new_n587_), .A4(new_n819_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n818_), .A2(new_n824_), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n479_), .A2(new_n513_), .A3(new_n540_), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT59), .B1(new_n826_), .B2(KEYINPUT119), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n825_), .B(new_n827_), .C1(KEYINPUT119), .C2(new_n826_), .ZN(new_n828_));
  AOI22_X1  g627(.A1(new_n817_), .A2(new_n341_), .B1(new_n821_), .B2(new_n823_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n826_), .ZN(new_n830_));
  OAI21_X1  g629(.A(KEYINPUT59), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n828_), .A2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(G113gat), .B1(new_n832_), .B2(new_n610_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT118), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n825_), .A2(new_n834_), .A3(new_n826_), .ZN(new_n835_));
  OAI21_X1  g634(.A(KEYINPUT118), .B1(new_n829_), .B2(new_n830_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  OR2_X1    g636(.A1(new_n606_), .A2(G113gat), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n833_), .B1(new_n837_), .B2(new_n838_), .ZN(G1340gat));
  NOR2_X1   g638(.A1(new_n587_), .A2(KEYINPUT60), .ZN(new_n840_));
  MUX2_X1   g639(.A(new_n840_), .B(KEYINPUT60), .S(G120gat), .Z(new_n841_));
  NAND3_X1  g640(.A1(new_n835_), .A2(new_n836_), .A3(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT120), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n842_), .B(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n828_), .A2(new_n588_), .A3(new_n831_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT121), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(G120gat), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n845_), .A2(new_n846_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n844_), .B1(new_n848_), .B2(new_n849_), .ZN(G1341gat));
  OAI21_X1  g649(.A(G127gat), .B1(new_n832_), .B2(new_n341_), .ZN(new_n851_));
  OR2_X1    g650(.A1(new_n341_), .A2(G127gat), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n851_), .B1(new_n837_), .B2(new_n852_), .ZN(G1342gat));
  OAI21_X1  g652(.A(G134gat), .B1(new_n832_), .B2(new_n673_), .ZN(new_n854_));
  OR2_X1    g653(.A1(new_n621_), .A2(G134gat), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n837_), .B2(new_n855_), .ZN(G1343gat));
  NOR4_X1   g655(.A1(new_n513_), .A2(new_n470_), .A3(new_n541_), .A4(new_n560_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n825_), .A2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n605_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g660(.A1(new_n859_), .A2(new_n588_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g662(.A1(new_n858_), .A2(new_n341_), .ZN(new_n864_));
  XOR2_X1   g663(.A(KEYINPUT61), .B(G155gat), .Z(new_n865_));
  XNOR2_X1  g664(.A(new_n864_), .B(new_n865_), .ZN(G1346gat));
  OAI21_X1  g665(.A(G162gat), .B1(new_n858_), .B2(new_n673_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n622_), .A2(new_n429_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n867_), .B1(new_n858_), .B2(new_n868_), .ZN(G1347gat));
  NAND4_X1  g668(.A1(new_n513_), .A2(new_n470_), .A3(new_n541_), .A4(new_n560_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n870_), .B1(new_n818_), .B2(new_n824_), .ZN(new_n871_));
  XOR2_X1   g670(.A(KEYINPUT22), .B(G169gat), .Z(new_n872_));
  NOR2_X1   g671(.A1(new_n606_), .A2(new_n872_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(KEYINPUT122), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n871_), .A2(new_n874_), .ZN(new_n875_));
  AOI211_X1 g674(.A(KEYINPUT62), .B(new_n356_), .C1(new_n871_), .C2(new_n605_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT62), .ZN(new_n877_));
  INV_X1    g676(.A(new_n870_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n825_), .A2(new_n605_), .A3(new_n878_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n877_), .B1(new_n879_), .B2(G169gat), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n875_), .B1(new_n876_), .B2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT123), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  OAI211_X1 g682(.A(KEYINPUT123), .B(new_n875_), .C1(new_n876_), .C2(new_n880_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(G1348gat));
  NAND2_X1  g684(.A1(new_n871_), .A2(new_n588_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g686(.A1(new_n871_), .A2(new_n669_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(G183gat), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n366_), .A2(new_n367_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n889_), .B1(new_n890_), .B2(new_n888_), .ZN(G1350gat));
  INV_X1    g690(.A(new_n871_), .ZN(new_n892_));
  OAI21_X1  g691(.A(G190gat), .B1(new_n892_), .B2(new_n673_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n622_), .A2(new_n359_), .ZN(new_n894_));
  XOR2_X1   g693(.A(new_n894_), .B(KEYINPUT124), .Z(new_n895_));
  OAI21_X1  g694(.A(new_n893_), .B1(new_n892_), .B2(new_n895_), .ZN(G1351gat));
  XNOR2_X1  g695(.A(KEYINPUT126), .B(G197gat), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  NOR4_X1   g697(.A1(new_n513_), .A2(new_n470_), .A3(new_n540_), .A4(new_n689_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n825_), .A2(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(KEYINPUT125), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT125), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n825_), .A2(new_n902_), .A3(new_n899_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n901_), .A2(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n898_), .B1(new_n905_), .B2(new_n606_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n904_), .A2(new_n605_), .A3(new_n897_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(G1352gat));
  OAI21_X1  g707(.A(G204gat), .B1(new_n905_), .B2(new_n587_), .ZN(new_n909_));
  INV_X1    g708(.A(G204gat), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n904_), .A2(new_n910_), .A3(new_n588_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n909_), .A2(new_n911_), .ZN(G1353gat));
  AOI21_X1  g711(.A(new_n341_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n913_));
  OAI21_X1  g712(.A(KEYINPUT127), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n914_));
  NOR3_X1   g713(.A1(KEYINPUT127), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  AOI22_X1  g715(.A1(new_n904_), .A2(new_n913_), .B1(new_n914_), .B2(new_n916_), .ZN(new_n917_));
  AND2_X1   g716(.A1(new_n904_), .A2(new_n913_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n917_), .B1(new_n918_), .B2(new_n916_), .ZN(G1354gat));
  OAI21_X1  g718(.A(G218gat), .B1(new_n905_), .B2(new_n673_), .ZN(new_n920_));
  INV_X1    g719(.A(G218gat), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n904_), .A2(new_n921_), .A3(new_n622_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n920_), .A2(new_n922_), .ZN(G1355gat));
endmodule


