//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 1 0 0 0 1 0 0 0 0 0 1 0 1 1 1 1 0 0 1 1 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 0 1 1 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n790_,
    new_n791_, new_n793_, new_n794_, new_n795_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n902_, new_n903_, new_n904_, new_n906_, new_n907_,
    new_n908_, new_n910_, new_n911_, new_n912_, new_n913_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n926_, new_n927_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n941_, new_n942_,
    new_n943_, new_n945_, new_n946_, new_n947_, new_n948_, new_n950_,
    new_n951_, new_n952_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n969_, new_n970_;
  INV_X1    g000(.A(KEYINPUT65), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT12), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT7), .ZN(new_n204_));
  INV_X1    g003(.A(G99gat), .ZN(new_n205_));
  INV_X1    g004(.A(G106gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT6), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n207_), .A2(new_n210_), .A3(new_n211_), .A4(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G85gat), .ZN(new_n214_));
  INV_X1    g013(.A(G92gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G85gat), .A2(G92gat), .ZN(new_n217_));
  AND2_X1   g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n213_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT8), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT8), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n213_), .A2(new_n221_), .A3(new_n218_), .ZN(new_n222_));
  AND2_X1   g021(.A1(new_n210_), .A2(new_n211_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n216_), .A2(KEYINPUT9), .A3(new_n217_), .ZN(new_n224_));
  AND2_X1   g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  XOR2_X1   g024(.A(KEYINPUT10), .B(G99gat), .Z(new_n226_));
  INV_X1    g025(.A(KEYINPUT9), .ZN(new_n227_));
  INV_X1    g026(.A(new_n217_), .ZN(new_n228_));
  AOI22_X1  g027(.A1(new_n226_), .A2(new_n206_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  AOI22_X1  g028(.A1(new_n220_), .A2(new_n222_), .B1(new_n225_), .B2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G57gat), .A2(G64gat), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(G57gat), .A2(G64gat), .ZN(new_n233_));
  NOR3_X1   g032(.A1(new_n232_), .A2(new_n233_), .A3(KEYINPUT64), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT64), .ZN(new_n235_));
  INV_X1    g034(.A(G57gat), .ZN(new_n236_));
  INV_X1    g035(.A(G64gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n235_), .B1(new_n238_), .B2(new_n231_), .ZN(new_n239_));
  OAI21_X1  g038(.A(KEYINPUT11), .B1(new_n234_), .B2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G71gat), .B(G78gat), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT64), .B1(new_n232_), .B2(new_n233_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n238_), .A2(new_n235_), .A3(new_n231_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT11), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n243_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n240_), .A2(new_n242_), .A3(new_n246_), .ZN(new_n247_));
  OAI211_X1 g046(.A(KEYINPUT11), .B(new_n241_), .C1(new_n234_), .C2(new_n239_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n203_), .B1(new_n230_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT67), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n226_), .A2(new_n206_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n228_), .A2(new_n227_), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n253_), .A2(new_n254_), .A3(new_n224_), .A4(new_n223_), .ZN(new_n255_));
  AND3_X1   g054(.A1(new_n213_), .A2(new_n221_), .A3(new_n218_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n221_), .B1(new_n213_), .B2(new_n218_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n255_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n258_), .A2(new_n248_), .A3(new_n247_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n259_), .A2(KEYINPUT67), .A3(new_n203_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n252_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G230gat), .A2(G233gat), .ZN(new_n262_));
  INV_X1    g061(.A(new_n249_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n263_), .A2(new_n258_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n258_), .A2(KEYINPUT12), .A3(new_n248_), .A4(new_n247_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT66), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n263_), .A2(KEYINPUT66), .A3(KEYINPUT12), .A4(new_n258_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n261_), .A2(new_n262_), .A3(new_n265_), .A4(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n265_), .A2(new_n259_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n262_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n202_), .B1(new_n271_), .B2(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(KEYINPUT65), .B1(new_n272_), .B2(new_n273_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G120gat), .B(G148gat), .ZN(new_n277_));
  INV_X1    g076(.A(G204gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  XOR2_X1   g078(.A(KEYINPUT5), .B(G176gat), .Z(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  OR3_X1    g081(.A1(new_n275_), .A2(new_n276_), .A3(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n282_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n284_));
  AND2_X1   g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT13), .ZN(new_n286_));
  OR2_X1    g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(new_n286_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G15gat), .B(G22gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G1gat), .A2(G8gat), .ZN(new_n291_));
  AND3_X1   g090(.A1(new_n291_), .A2(KEYINPUT71), .A3(KEYINPUT14), .ZN(new_n292_));
  AOI21_X1  g091(.A(KEYINPUT71), .B1(new_n291_), .B2(KEYINPUT14), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n290_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G1gat), .B(G8gat), .ZN(new_n295_));
  OR2_X1    g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n295_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G29gat), .B(G36gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G43gat), .B(G50gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n298_), .B(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n303_), .A2(G229gat), .A3(G233gat), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n298_), .A2(new_n302_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G229gat), .A2(G233gat), .ZN(new_n307_));
  INV_X1    g106(.A(new_n298_), .ZN(new_n308_));
  XOR2_X1   g107(.A(new_n301_), .B(KEYINPUT15), .Z(new_n309_));
  OAI211_X1 g108(.A(new_n306_), .B(new_n307_), .C1(new_n308_), .C2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n304_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G113gat), .B(G141gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G169gat), .B(G197gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n312_), .A2(new_n316_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n311_), .A2(new_n315_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n289_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT80), .ZN(new_n322_));
  INV_X1    g121(.A(G169gat), .ZN(new_n323_));
  INV_X1    g122(.A(G176gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G169gat), .A2(G176gat), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n325_), .A2(KEYINPUT24), .A3(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT23), .ZN(new_n328_));
  INV_X1    g127(.A(G183gat), .ZN(new_n329_));
  INV_X1    g128(.A(G190gat), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n328_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n332_));
  OR3_X1    g131(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n327_), .A2(new_n331_), .A3(new_n332_), .A4(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT25), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(G183gat), .ZN(new_n337_));
  OR2_X1    g136(.A1(new_n337_), .A2(KEYINPUT76), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT77), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(G190gat), .ZN(new_n340_));
  AOI22_X1  g139(.A1(new_n340_), .A2(KEYINPUT26), .B1(KEYINPUT25), .B2(new_n329_), .ZN(new_n341_));
  OR3_X1    g140(.A1(new_n330_), .A2(KEYINPUT77), .A3(KEYINPUT26), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n337_), .A2(KEYINPUT76), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n338_), .A2(new_n341_), .A3(new_n342_), .A4(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n335_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n326_), .ZN(new_n346_));
  AND2_X1   g145(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n347_));
  NOR2_X1   g146(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n324_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n346_), .B1(new_n349_), .B2(KEYINPUT78), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT78), .ZN(new_n351_));
  OAI211_X1 g150(.A(new_n351_), .B(new_n324_), .C1(new_n347_), .C2(new_n348_), .ZN(new_n352_));
  OAI211_X1 g151(.A(new_n331_), .B(new_n332_), .C1(G183gat), .C2(G190gat), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n350_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n345_), .A2(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT79), .B(KEYINPUT30), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n356_), .B1(new_n345_), .B2(new_n354_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n322_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n359_), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n353_), .A2(new_n352_), .ZN(new_n362_));
  AOI22_X1  g161(.A1(new_n362_), .A2(new_n350_), .B1(new_n335_), .B2(new_n344_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(new_n356_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n361_), .A2(new_n364_), .A3(KEYINPUT80), .ZN(new_n365_));
  XOR2_X1   g164(.A(G15gat), .B(G43gat), .Z(new_n366_));
  NAND2_X1  g165(.A1(G227gat), .A2(G233gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  XOR2_X1   g167(.A(G71gat), .B(G99gat), .Z(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n360_), .A2(new_n365_), .A3(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(G113gat), .A2(G120gat), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G113gat), .A2(G120gat), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n373_), .A2(KEYINPUT81), .A3(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT81), .ZN(new_n376_));
  INV_X1    g175(.A(new_n374_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n376_), .B1(new_n377_), .B2(new_n372_), .ZN(new_n378_));
  XOR2_X1   g177(.A(G127gat), .B(G134gat), .Z(new_n379_));
  AND3_X1   g178(.A1(new_n375_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n379_), .B1(new_n375_), .B2(new_n378_), .ZN(new_n381_));
  OAI21_X1  g180(.A(KEYINPUT82), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n375_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT82), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  AND2_X1   g184(.A1(new_n382_), .A2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT31), .ZN(new_n387_));
  INV_X1    g186(.A(new_n370_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n388_), .A2(KEYINPUT80), .A3(new_n364_), .A4(new_n361_), .ZN(new_n389_));
  AND3_X1   g188(.A1(new_n371_), .A2(new_n387_), .A3(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n387_), .B1(new_n371_), .B2(new_n389_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G225gat), .A2(G233gat), .ZN(new_n393_));
  XOR2_X1   g192(.A(new_n393_), .B(KEYINPUT95), .Z(new_n394_));
  INV_X1    g193(.A(KEYINPUT4), .ZN(new_n395_));
  OR2_X1    g194(.A1(G155gat), .A2(G162gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G155gat), .A2(G162gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT3), .ZN(new_n399_));
  INV_X1    g198(.A(G141gat), .ZN(new_n400_));
  INV_X1    g199(.A(G148gat), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n399_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n403_));
  OAI21_X1  g202(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n402_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G141gat), .A2(G148gat), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT2), .ZN(new_n407_));
  AND2_X1   g206(.A1(new_n407_), .A2(KEYINPUT84), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n407_), .A2(KEYINPUT84), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n406_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT85), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n405_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  OAI211_X1 g211(.A(KEYINPUT85), .B(new_n406_), .C1(new_n408_), .C2(new_n409_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n398_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT83), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n415_), .B1(new_n397_), .B2(KEYINPUT1), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n397_), .A2(KEYINPUT1), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT1), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n418_), .A2(KEYINPUT83), .A3(G155gat), .A4(G162gat), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n416_), .A2(new_n417_), .A3(new_n419_), .A4(new_n396_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n406_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(G141gat), .A2(G148gat), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n420_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n382_), .B(new_n385_), .C1(new_n414_), .C2(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(KEYINPUT84), .B(KEYINPUT2), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n411_), .B1(new_n427_), .B2(new_n421_), .ZN(new_n428_));
  AND3_X1   g227(.A1(new_n402_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n428_), .A2(new_n429_), .A3(new_n413_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n398_), .ZN(new_n431_));
  AOI22_X1  g230(.A1(new_n430_), .A2(new_n431_), .B1(new_n420_), .B2(new_n423_), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT94), .B1(new_n380_), .B2(new_n381_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n375_), .A2(new_n378_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n379_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT94), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n436_), .A2(new_n437_), .A3(new_n383_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n432_), .A2(new_n433_), .A3(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n395_), .B1(new_n426_), .B2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n430_), .A2(new_n431_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(new_n424_), .ZN(new_n442_));
  AOI21_X1  g241(.A(KEYINPUT4), .B1(new_n386_), .B2(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n394_), .B1(new_n440_), .B2(new_n443_), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n426_), .A2(new_n439_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(new_n393_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n444_), .A2(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G1gat), .B(G29gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G57gat), .B(G85gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n450_), .B(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n447_), .A2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n444_), .A2(new_n446_), .A3(new_n452_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G8gat), .B(G36gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(new_n215_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(KEYINPUT18), .B(G64gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT32), .ZN(new_n461_));
  XNOR2_X1  g260(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G226gat), .A2(G233gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(G211gat), .A2(G218gat), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT86), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G211gat), .A2(G218gat), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n466_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n468_), .ZN(new_n470_));
  OAI21_X1  g269(.A(KEYINPUT86), .B1(new_n470_), .B2(new_n465_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n278_), .A2(G197gat), .ZN(new_n472_));
  INV_X1    g271(.A(G197gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(G204gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  AOI22_X1  g274(.A1(new_n469_), .A2(new_n471_), .B1(KEYINPUT21), .B2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G197gat), .B(G204gat), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT21), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  AND2_X1   g278(.A1(new_n469_), .A2(new_n471_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n476_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n355_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT20), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n353_), .B1(KEYINPUT92), .B2(new_n326_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT92), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n346_), .B1(new_n349_), .B2(new_n485_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n484_), .A2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(KEYINPUT26), .B(G190gat), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n329_), .A2(KEYINPUT25), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(new_n337_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT90), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT90), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n490_), .A2(new_n337_), .A3(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n489_), .B1(new_n492_), .B2(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n495_), .A2(new_n334_), .ZN(new_n496_));
  NOR3_X1   g295(.A1(new_n481_), .A2(new_n487_), .A3(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n464_), .B1(new_n483_), .B2(new_n497_), .ZN(new_n498_));
  OR2_X1    g297(.A1(new_n484_), .A2(new_n486_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT91), .ZN(new_n500_));
  NOR3_X1   g299(.A1(new_n495_), .A2(new_n500_), .A3(new_n334_), .ZN(new_n501_));
  AND3_X1   g300(.A1(new_n490_), .A2(new_n337_), .A3(new_n493_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n493_), .B1(new_n490_), .B2(new_n337_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n488_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(KEYINPUT91), .B1(new_n335_), .B2(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n499_), .B1(new_n501_), .B2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(new_n481_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n464_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT20), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n477_), .A2(new_n478_), .ZN(new_n510_));
  AND3_X1   g309(.A1(new_n472_), .A2(new_n474_), .A3(new_n478_), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n471_), .B(new_n469_), .C1(new_n510_), .C2(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n512_), .B1(new_n510_), .B2(new_n480_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n509_), .B1(new_n363_), .B2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n507_), .A2(new_n508_), .A3(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n461_), .B1(new_n498_), .B2(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n508_), .B1(new_n507_), .B2(new_n514_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n464_), .A2(new_n509_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n518_), .B1(new_n363_), .B2(new_n513_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n505_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n335_), .A2(new_n504_), .A3(KEYINPUT91), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n487_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n519_), .B1(new_n522_), .B2(new_n513_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n517_), .A2(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n516_), .B1(new_n524_), .B2(new_n461_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n456_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n460_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n527_), .B1(new_n517_), .B2(new_n523_), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n482_), .B(new_n518_), .C1(new_n506_), .C2(new_n481_), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT20), .B1(new_n355_), .B2(new_n481_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n530_), .B1(new_n481_), .B2(new_n506_), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n460_), .B(new_n529_), .C1(new_n531_), .C2(new_n508_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n528_), .A2(new_n532_), .A3(KEYINPUT93), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT93), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n524_), .A2(new_n534_), .A3(new_n460_), .ZN(new_n535_));
  AND2_X1   g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT33), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n455_), .A2(new_n537_), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n444_), .A2(KEYINPUT33), .A3(new_n446_), .A4(new_n452_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n452_), .B1(new_n445_), .B2(new_n394_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n393_), .B1(new_n440_), .B2(new_n443_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n538_), .A2(new_n539_), .A3(new_n542_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n526_), .B1(new_n536_), .B2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G22gat), .B(G50gat), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT28), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT29), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n432_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n547_), .B1(new_n432_), .B2(new_n548_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n546_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n551_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n553_), .A2(new_n549_), .A3(new_n545_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n552_), .A2(new_n554_), .ZN(new_n555_));
  XOR2_X1   g354(.A(G78gat), .B(G106gat), .Z(new_n556_));
  NAND2_X1  g355(.A1(G228gat), .A2(G233gat), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n442_), .A2(KEYINPUT29), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n557_), .B1(new_n558_), .B2(new_n481_), .ZN(new_n559_));
  OAI211_X1 g358(.A(new_n557_), .B(new_n481_), .C1(new_n432_), .C2(new_n548_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n556_), .B1(new_n559_), .B2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n557_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n548_), .B1(new_n441_), .B2(new_n424_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n563_), .B1(new_n564_), .B2(new_n513_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n556_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n565_), .A2(new_n560_), .A3(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n555_), .A2(new_n562_), .A3(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n566_), .A2(KEYINPUT88), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n565_), .A2(new_n560_), .A3(new_n569_), .ZN(new_n570_));
  AND3_X1   g369(.A1(new_n570_), .A2(new_n552_), .A3(new_n554_), .ZN(new_n571_));
  OAI211_X1 g370(.A(KEYINPUT88), .B(new_n566_), .C1(new_n559_), .C2(new_n561_), .ZN(new_n572_));
  AOI22_X1  g371(.A1(new_n568_), .A2(KEYINPUT87), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT87), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n555_), .A2(new_n562_), .A3(new_n574_), .A4(new_n567_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n573_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n544_), .A2(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n456_), .B1(new_n573_), .B2(new_n575_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT27), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n533_), .A2(new_n580_), .A3(new_n535_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(KEYINPUT98), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT98), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n533_), .A2(new_n535_), .A3(new_n583_), .A4(new_n580_), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n532_), .A2(KEYINPUT97), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n532_), .A2(KEYINPUT97), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n498_), .A2(new_n515_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n580_), .B1(new_n587_), .B2(new_n527_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n585_), .A2(new_n586_), .A3(new_n588_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n579_), .A2(new_n582_), .A3(new_n584_), .A4(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n392_), .B1(new_n578_), .B2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n573_), .A2(new_n575_), .A3(new_n392_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n592_), .A2(new_n456_), .ZN(new_n593_));
  AND4_X1   g392(.A1(new_n593_), .A2(new_n584_), .A3(new_n589_), .A4(new_n582_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n591_), .A2(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n321_), .A2(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G183gat), .B(G211gat), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(G231gat), .A2(G233gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT72), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n298_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n298_), .A2(new_n601_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n249_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n604_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n606_), .A2(new_n263_), .A3(new_n602_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n598_), .B1(new_n608_), .B2(KEYINPUT74), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n608_), .A2(KEYINPUT74), .A3(new_n598_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G127gat), .B(G155gat), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n612_), .B(new_n613_), .Z(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n610_), .A2(new_n611_), .A3(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n615_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n618_));
  OAI21_X1  g417(.A(KEYINPUT17), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n618_), .ZN(new_n620_));
  AOI21_X1  g419(.A(KEYINPUT17), .B1(new_n605_), .B2(new_n607_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n620_), .A2(new_n616_), .A3(new_n621_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n619_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT36), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n230_), .A2(new_n301_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n625_), .B1(new_n309_), .B2(new_n230_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(G232gat), .A2(G233gat), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n628_), .B(KEYINPUT34), .Z(new_n629_));
  INV_X1    g428(.A(KEYINPUT35), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n632_), .A2(KEYINPUT68), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n632_), .A2(KEYINPUT68), .ZN(new_n634_));
  AOI211_X1 g433(.A(new_n633_), .B(new_n634_), .C1(new_n630_), .C2(new_n629_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n627_), .A2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(KEYINPUT69), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT69), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n627_), .A2(new_n638_), .A3(new_n635_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(new_n640_));
  XOR2_X1   g439(.A(G190gat), .B(G218gat), .Z(new_n641_));
  XOR2_X1   g440(.A(G134gat), .B(G162gat), .Z(new_n642_));
  XOR2_X1   g441(.A(new_n641_), .B(new_n642_), .Z(new_n643_));
  NOR2_X1   g442(.A1(new_n627_), .A2(new_n632_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  AND4_X1   g444(.A1(new_n624_), .A2(new_n640_), .A3(new_n643_), .A4(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n644_), .B1(new_n637_), .B2(new_n639_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n643_), .B(new_n624_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT70), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(KEYINPUT37), .B1(new_n646_), .B2(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n647_), .A2(new_n624_), .A3(new_n643_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT37), .ZN(new_n653_));
  OAI211_X1 g452(.A(new_n652_), .B(new_n653_), .C1(new_n647_), .C2(new_n648_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n651_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n623_), .A2(new_n655_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT75), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n596_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT38), .ZN(new_n659_));
  INV_X1    g458(.A(new_n456_), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n660_), .A2(G1gat), .ZN(new_n661_));
  OR3_X1    g460(.A1(new_n658_), .A2(new_n659_), .A3(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n319_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n578_), .A2(new_n590_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n392_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  AND3_X1   g465(.A1(new_n582_), .A2(new_n584_), .A3(new_n589_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(new_n593_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n623_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n652_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n670_), .A2(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n663_), .A2(new_n669_), .A3(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(G1gat), .B1(new_n674_), .B2(new_n660_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n659_), .B1(new_n658_), .B2(new_n661_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n662_), .A2(new_n675_), .A3(new_n676_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT99), .ZN(G1324gat));
  OR3_X1    g477(.A1(new_n658_), .A2(G8gat), .A3(new_n667_), .ZN(new_n679_));
  OAI21_X1  g478(.A(G8gat), .B1(new_n674_), .B2(new_n667_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(KEYINPUT100), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT100), .ZN(new_n682_));
  OAI211_X1 g481(.A(new_n682_), .B(G8gat), .C1(new_n674_), .C2(new_n667_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n681_), .A2(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n684_), .A2(KEYINPUT101), .A3(KEYINPUT39), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n685_), .B1(KEYINPUT39), .B2(new_n684_), .ZN(new_n686_));
  AOI21_X1  g485(.A(KEYINPUT101), .B1(new_n684_), .B2(KEYINPUT39), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n679_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT40), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  OAI211_X1 g489(.A(KEYINPUT40), .B(new_n679_), .C1(new_n686_), .C2(new_n687_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1325gat));
  OR2_X1    g491(.A1(new_n665_), .A2(G15gat), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n658_), .A2(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(G15gat), .B1(new_n674_), .B2(new_n665_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(KEYINPUT41), .B2(new_n695_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n696_), .B1(KEYINPUT41), .B2(new_n695_), .ZN(new_n697_));
  XOR2_X1   g496(.A(new_n697_), .B(KEYINPUT102), .Z(G1326gat));
  OAI21_X1  g497(.A(G22gat), .B1(new_n674_), .B2(new_n577_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT42), .Z(new_n700_));
  NOR3_X1   g499(.A1(new_n658_), .A2(G22gat), .A3(new_n577_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT103), .Z(G1327gat));
  INV_X1    g502(.A(KEYINPUT104), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT43), .ZN(new_n705_));
  INV_X1    g504(.A(new_n655_), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n669_), .A2(new_n704_), .A3(new_n705_), .A4(new_n706_), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n705_), .B(new_n706_), .C1(new_n591_), .C2(new_n594_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(KEYINPUT104), .ZN(new_n709_));
  OAI21_X1  g508(.A(KEYINPUT43), .B1(new_n595_), .B2(new_n655_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n707_), .A2(new_n709_), .A3(new_n710_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n321_), .A2(new_n623_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n711_), .A2(KEYINPUT44), .A3(new_n712_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n715_), .A2(new_n456_), .A3(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(KEYINPUT105), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT105), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n715_), .A2(new_n719_), .A3(new_n456_), .A4(new_n716_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n718_), .A2(G29gat), .A3(new_n720_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n623_), .A2(new_n671_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT106), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n596_), .A2(new_n723_), .ZN(new_n724_));
  OR3_X1    g523(.A1(new_n724_), .A2(G29gat), .A3(new_n660_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n721_), .A2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT107), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT107), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n721_), .A2(new_n728_), .A3(new_n725_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(G1328gat));
  INV_X1    g529(.A(new_n667_), .ZN(new_n731_));
  INV_X1    g530(.A(G36gat), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n724_), .A2(new_n733_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT45), .Z(new_n735_));
  NAND2_X1  g534(.A1(new_n715_), .A2(new_n716_), .ZN(new_n736_));
  OAI21_X1  g535(.A(G36gat), .B1(new_n736_), .B2(new_n667_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT46), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n738_), .B(new_n739_), .ZN(G1329gat));
  OAI21_X1  g539(.A(G43gat), .B1(new_n736_), .B2(new_n665_), .ZN(new_n741_));
  INV_X1    g540(.A(G43gat), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n392_), .A2(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n741_), .B1(new_n724_), .B2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n744_), .B(new_n746_), .ZN(G1330gat));
  OR3_X1    g546(.A1(new_n724_), .A2(G50gat), .A3(new_n577_), .ZN(new_n748_));
  OAI21_X1  g547(.A(G50gat), .B1(new_n736_), .B2(new_n577_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n749_), .A2(KEYINPUT109), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n749_), .A2(KEYINPUT109), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n748_), .B1(new_n750_), .B2(new_n751_), .ZN(G1331gat));
  NOR3_X1   g551(.A1(new_n595_), .A2(new_n289_), .A3(new_n320_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(new_n657_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n236_), .B1(new_n754_), .B2(new_n660_), .ZN(new_n755_));
  XOR2_X1   g554(.A(new_n755_), .B(KEYINPUT110), .Z(new_n756_));
  NAND2_X1  g555(.A1(new_n753_), .A2(new_n673_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(KEYINPUT111), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT111), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n753_), .A2(new_n759_), .A3(new_n673_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n758_), .A2(new_n760_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n660_), .A2(new_n236_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n756_), .B1(new_n761_), .B2(new_n762_), .ZN(G1332gat));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n731_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(G64gat), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n765_), .A2(KEYINPUT48), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n765_), .A2(KEYINPUT48), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n731_), .A2(new_n237_), .ZN(new_n768_));
  OAI22_X1  g567(.A1(new_n766_), .A2(new_n767_), .B1(new_n754_), .B2(new_n768_), .ZN(G1333gat));
  OR3_X1    g568(.A1(new_n754_), .A2(G71gat), .A3(new_n665_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n758_), .A2(new_n392_), .A3(new_n760_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT49), .ZN(new_n772_));
  AND3_X1   g571(.A1(new_n771_), .A2(new_n772_), .A3(G71gat), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n772_), .B1(new_n771_), .B2(G71gat), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n770_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT112), .ZN(G1334gat));
  OR3_X1    g575(.A1(new_n754_), .A2(G78gat), .A3(new_n577_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n761_), .A2(new_n576_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(G78gat), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n779_), .A2(KEYINPUT50), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n779_), .A2(KEYINPUT50), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n777_), .B1(new_n780_), .B2(new_n781_), .ZN(G1335gat));
  NOR3_X1   g581(.A1(new_n289_), .A2(new_n320_), .A3(new_n623_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n711_), .A2(new_n783_), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n784_), .A2(new_n214_), .A3(new_n660_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n723_), .A2(new_n753_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(G85gat), .B1(new_n787_), .B2(new_n456_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n785_), .A2(new_n788_), .ZN(G1336gat));
  NOR3_X1   g588(.A1(new_n784_), .A2(new_n215_), .A3(new_n667_), .ZN(new_n790_));
  AOI21_X1  g589(.A(G92gat), .B1(new_n787_), .B2(new_n731_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n790_), .A2(new_n791_), .ZN(G1337gat));
  OAI21_X1  g591(.A(G99gat), .B1(new_n784_), .B2(new_n665_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n787_), .A2(new_n226_), .A3(new_n392_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g595(.A1(new_n787_), .A2(new_n206_), .A3(new_n576_), .ZN(new_n797_));
  OAI21_X1  g596(.A(G106gat), .B1(new_n784_), .B2(new_n577_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n798_), .A2(KEYINPUT52), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n798_), .A2(KEYINPUT52), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n797_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n801_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g601(.A1(new_n275_), .A2(new_n276_), .A3(new_n282_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n318_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n316_), .B1(new_n303_), .B2(new_n307_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n306_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n805_), .B1(new_n307_), .B2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n804_), .A2(new_n807_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n803_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n264_), .B1(new_n252_), .B2(new_n260_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n811_), .A2(KEYINPUT55), .A3(new_n262_), .A4(new_n270_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n261_), .A2(new_n265_), .A3(new_n270_), .ZN(new_n813_));
  AOI22_X1  g612(.A1(new_n812_), .A2(KEYINPUT116), .B1(new_n273_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT55), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n271_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT115), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n271_), .A2(KEYINPUT115), .A3(new_n815_), .ZN(new_n819_));
  AND3_X1   g618(.A1(new_n261_), .A2(new_n265_), .A3(new_n270_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n820_), .A2(new_n821_), .A3(KEYINPUT55), .A4(new_n262_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n814_), .A2(new_n818_), .A3(new_n819_), .A4(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n282_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT56), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n823_), .A2(KEYINPUT56), .A3(new_n282_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n810_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(KEYINPUT58), .B1(new_n828_), .B2(KEYINPUT117), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n823_), .A2(KEYINPUT56), .A3(new_n282_), .ZN(new_n830_));
  AOI21_X1  g629(.A(KEYINPUT56), .B1(new_n823_), .B2(new_n282_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n809_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT117), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT58), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n832_), .A2(new_n833_), .A3(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n829_), .A2(new_n706_), .A3(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT57), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n285_), .A2(new_n808_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n826_), .A2(new_n827_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n283_), .A2(new_n320_), .A3(KEYINPUT114), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT114), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n841_), .B1(new_n803_), .B2(new_n319_), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n840_), .A2(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n838_), .B1(new_n839_), .B2(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n837_), .B1(new_n844_), .B2(new_n672_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n840_), .A2(new_n842_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n846_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n847_));
  OAI211_X1 g646(.A(KEYINPUT57), .B(new_n671_), .C1(new_n847_), .C2(new_n838_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n836_), .A2(new_n845_), .A3(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n619_), .A2(new_n622_), .A3(new_n319_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n706_), .B1(KEYINPUT113), .B2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT113), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n623_), .A2(new_n852_), .A3(new_n319_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n851_), .A2(new_n289_), .A3(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(KEYINPUT54), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT54), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n851_), .A2(new_n856_), .A3(new_n289_), .A4(new_n853_), .ZN(new_n857_));
  AOI22_X1  g656(.A1(new_n849_), .A2(new_n670_), .B1(new_n855_), .B2(new_n857_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n731_), .A2(new_n660_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  NOR3_X1   g659(.A1(new_n858_), .A2(new_n592_), .A3(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(G113gat), .B1(new_n861_), .B2(new_n320_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n849_), .A2(new_n670_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n855_), .A2(new_n857_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n860_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n592_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(KEYINPUT59), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT59), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n861_), .A2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n868_), .A2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  AND2_X1   g671(.A1(new_n320_), .A2(G113gat), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n862_), .B1(new_n872_), .B2(new_n873_), .ZN(G1340gat));
  OAI21_X1  g673(.A(G120gat), .B1(new_n871_), .B2(new_n289_), .ZN(new_n875_));
  INV_X1    g674(.A(G120gat), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n876_), .B1(new_n289_), .B2(KEYINPUT60), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n877_), .B1(KEYINPUT60), .B2(new_n876_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n875_), .B1(new_n867_), .B2(new_n878_), .ZN(G1341gat));
  AOI21_X1  g678(.A(G127gat), .B1(new_n861_), .B2(new_n623_), .ZN(new_n880_));
  AND2_X1   g679(.A1(new_n623_), .A2(G127gat), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n880_), .B1(new_n872_), .B2(new_n881_), .ZN(G1342gat));
  INV_X1    g681(.A(KEYINPUT118), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n869_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n884_));
  NOR4_X1   g683(.A1(new_n858_), .A2(KEYINPUT59), .A3(new_n592_), .A4(new_n860_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n706_), .A2(G134gat), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n884_), .A2(new_n885_), .A3(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(G134gat), .B1(new_n861_), .B2(new_n672_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n883_), .B1(new_n887_), .B2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(G134gat), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n890_), .B1(new_n867_), .B2(new_n671_), .ZN(new_n891_));
  OAI211_X1 g690(.A(KEYINPUT118), .B(new_n891_), .C1(new_n871_), .C2(new_n886_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n889_), .A2(new_n892_), .ZN(G1343gat));
  NAND2_X1  g692(.A1(new_n863_), .A2(new_n864_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n577_), .A2(new_n392_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n894_), .A2(new_n859_), .A3(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT119), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n865_), .A2(KEYINPUT119), .A3(new_n895_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n319_), .B1(new_n898_), .B2(new_n899_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(new_n400_), .ZN(G1344gat));
  AOI21_X1  g700(.A(new_n289_), .B1(new_n898_), .B2(new_n899_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(KEYINPUT120), .B(G148gat), .ZN(new_n903_));
  INV_X1    g702(.A(new_n903_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n902_), .B(new_n904_), .ZN(G1345gat));
  AOI21_X1  g704(.A(new_n670_), .B1(new_n898_), .B2(new_n899_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(KEYINPUT61), .B(G155gat), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n906_), .B(new_n908_), .ZN(G1346gat));
  NAND2_X1  g708(.A1(new_n898_), .A2(new_n899_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(new_n672_), .ZN(new_n911_));
  INV_X1    g710(.A(G162gat), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n655_), .A2(new_n912_), .ZN(new_n913_));
  AOI22_X1  g712(.A1(new_n911_), .A2(new_n912_), .B1(new_n910_), .B2(new_n913_), .ZN(G1347gat));
  NAND4_X1  g713(.A1(new_n894_), .A2(new_n320_), .A3(new_n593_), .A4(new_n731_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT121), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT62), .ZN(new_n917_));
  NAND4_X1  g716(.A1(new_n915_), .A2(new_n916_), .A3(new_n917_), .A4(G169gat), .ZN(new_n918_));
  INV_X1    g717(.A(new_n593_), .ZN(new_n919_));
  NOR3_X1   g718(.A1(new_n858_), .A2(new_n919_), .A3(new_n667_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n323_), .B1(new_n920_), .B2(new_n320_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n918_), .B1(new_n921_), .B2(new_n917_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n916_), .B1(new_n921_), .B2(new_n917_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n347_), .A2(new_n348_), .ZN(new_n924_));
  OAI22_X1  g723(.A1(new_n922_), .A2(new_n923_), .B1(new_n924_), .B2(new_n915_), .ZN(G1348gat));
  INV_X1    g724(.A(new_n289_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n920_), .A2(new_n926_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(G176gat), .ZN(G1349gat));
  INV_X1    g727(.A(KEYINPUT122), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n502_), .A2(new_n503_), .ZN(new_n930_));
  NAND4_X1  g729(.A1(new_n920_), .A2(new_n929_), .A3(new_n930_), .A4(new_n623_), .ZN(new_n931_));
  NAND4_X1  g730(.A1(new_n894_), .A2(new_n593_), .A3(new_n731_), .A4(new_n623_), .ZN(new_n932_));
  AOI21_X1  g731(.A(KEYINPUT122), .B1(new_n932_), .B2(new_n329_), .ZN(new_n933_));
  INV_X1    g732(.A(new_n930_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n932_), .A2(new_n934_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n931_), .B1(new_n933_), .B2(new_n935_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n936_), .A2(KEYINPUT123), .ZN(new_n937_));
  INV_X1    g736(.A(KEYINPUT123), .ZN(new_n938_));
  OAI211_X1 g737(.A(new_n938_), .B(new_n931_), .C1(new_n933_), .C2(new_n935_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n937_), .A2(new_n939_), .ZN(G1350gat));
  INV_X1    g739(.A(new_n920_), .ZN(new_n941_));
  OAI21_X1  g740(.A(G190gat), .B1(new_n941_), .B2(new_n655_), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n920_), .A2(new_n488_), .A3(new_n672_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n942_), .A2(new_n943_), .ZN(G1351gat));
  NAND2_X1  g743(.A1(new_n579_), .A2(new_n665_), .ZN(new_n945_));
  NOR3_X1   g744(.A1(new_n858_), .A2(new_n667_), .A3(new_n945_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n946_), .A2(new_n320_), .ZN(new_n947_));
  XNOR2_X1  g746(.A(KEYINPUT124), .B(G197gat), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n947_), .B(new_n948_), .ZN(G1352gat));
  AND2_X1   g748(.A1(new_n946_), .A2(new_n926_), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n950_), .B1(KEYINPUT125), .B2(new_n278_), .ZN(new_n951_));
  XNOR2_X1  g750(.A(KEYINPUT125), .B(G204gat), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n951_), .B1(new_n950_), .B2(new_n952_), .ZN(G1353gat));
  INV_X1    g752(.A(new_n945_), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n670_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n955_));
  NAND4_X1  g754(.A1(new_n894_), .A2(new_n731_), .A3(new_n954_), .A4(new_n955_), .ZN(new_n956_));
  INV_X1    g755(.A(KEYINPUT126), .ZN(new_n957_));
  OAI21_X1  g756(.A(KEYINPUT127), .B1(new_n956_), .B2(new_n957_), .ZN(new_n958_));
  INV_X1    g757(.A(new_n958_), .ZN(new_n959_));
  NOR3_X1   g758(.A1(new_n956_), .A2(new_n957_), .A3(KEYINPUT127), .ZN(new_n960_));
  INV_X1    g759(.A(new_n956_), .ZN(new_n961_));
  NOR2_X1   g760(.A1(new_n961_), .A2(KEYINPUT126), .ZN(new_n962_));
  NOR2_X1   g761(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n963_));
  OAI22_X1  g762(.A1(new_n959_), .A2(new_n960_), .B1(new_n962_), .B2(new_n963_), .ZN(new_n964_));
  INV_X1    g763(.A(new_n960_), .ZN(new_n965_));
  AOI21_X1  g764(.A(new_n963_), .B1(new_n956_), .B2(new_n957_), .ZN(new_n966_));
  NAND3_X1  g765(.A1(new_n965_), .A2(new_n966_), .A3(new_n958_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n964_), .A2(new_n967_), .ZN(G1354gat));
  AOI21_X1  g767(.A(G218gat), .B1(new_n946_), .B2(new_n672_), .ZN(new_n969_));
  AND2_X1   g768(.A1(new_n706_), .A2(G218gat), .ZN(new_n970_));
  AOI21_X1  g769(.A(new_n969_), .B1(new_n946_), .B2(new_n970_), .ZN(G1355gat));
endmodule


