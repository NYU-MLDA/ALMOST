//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 0 0 1 1 1 0 1 1 0 1 0 0 0 0 1 0 1 0 1 1 1 1 0 0 1 1 1 0 0 1 0 0 0 1 1 0 0 1 1 0 0 1 0 0 1 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n814_,
    new_n815_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n907_, new_n908_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n925_, new_n926_, new_n927_, new_n928_, new_n930_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n942_, new_n943_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n956_, new_n957_, new_n958_,
    new_n959_, new_n961_, new_n962_, new_n963_, new_n965_, new_n966_,
    new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n977_, new_n978_, new_n979_, new_n980_,
    new_n981_, new_n983_, new_n984_, new_n985_, new_n987_, new_n988_,
    new_n989_;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202_));
  OR2_X1    g001(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n204_));
  XOR2_X1   g003(.A(G71gat), .B(G78gat), .Z(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n204_), .A2(new_n205_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT8), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT6), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT6), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n213_), .A2(G99gat), .A3(G106gat), .ZN(new_n214_));
  AND2_X1   g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT66), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n212_), .A2(new_n214_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT66), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G99gat), .A2(G106gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(KEYINPUT7), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n217_), .A2(new_n219_), .A3(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(G85gat), .ZN(new_n223_));
  INV_X1    g022(.A(G92gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G85gat), .A2(G92gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n210_), .B1(new_n222_), .B2(new_n228_), .ZN(new_n229_));
  AOI211_X1 g028(.A(KEYINPUT8), .B(new_n227_), .C1(new_n221_), .C2(new_n218_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND4_X1  g030(.A1(KEYINPUT64), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT9), .ZN(new_n233_));
  AOI21_X1  g032(.A(KEYINPUT64), .B1(new_n226_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n233_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n232_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT65), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  OAI211_X1 g038(.A(KEYINPUT65), .B(new_n232_), .C1(new_n236_), .C2(new_n235_), .ZN(new_n240_));
  INV_X1    g039(.A(G106gat), .ZN(new_n241_));
  XOR2_X1   g040(.A(KEYINPUT10), .B(G99gat), .Z(new_n242_));
  AOI21_X1  g041(.A(new_n215_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n239_), .A2(new_n240_), .A3(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n209_), .B1(new_n231_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n230_), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n219_), .A2(new_n221_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n227_), .B1(new_n248_), .B2(new_n217_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n247_), .B1(new_n249_), .B2(new_n210_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n250_), .A2(new_n208_), .A3(new_n244_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n246_), .A2(new_n251_), .A3(KEYINPUT12), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n244_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT12), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n253_), .A2(new_n254_), .A3(new_n209_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n252_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G230gat), .A2(G233gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n246_), .A2(new_n251_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n257_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n258_), .A2(new_n261_), .ZN(new_n262_));
  XOR2_X1   g061(.A(G120gat), .B(G148gat), .Z(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G176gat), .B(G204gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n262_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n267_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n258_), .A2(new_n261_), .A3(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n268_), .A2(KEYINPUT13), .A3(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(KEYINPUT13), .B1(new_n268_), .B2(new_n270_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n274_), .A2(KEYINPUT68), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(KEYINPUT68), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT37), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G190gat), .B(G218gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G134gat), .B(G162gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  XOR2_X1   g080(.A(new_n281_), .B(KEYINPUT36), .Z(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G29gat), .B(G36gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G43gat), .B(G50gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT15), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n253_), .A2(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n250_), .A2(new_n286_), .A3(new_n244_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G232gat), .A2(G233gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT34), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT35), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n289_), .A2(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n292_), .A2(new_n293_), .ZN(new_n296_));
  NOR3_X1   g095(.A1(new_n288_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n296_), .B1(new_n288_), .B2(new_n295_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n283_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n299_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n281_), .A2(KEYINPUT36), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NOR3_X1   g102(.A1(new_n301_), .A2(new_n303_), .A3(new_n297_), .ZN(new_n304_));
  OAI211_X1 g103(.A(KEYINPUT69), .B(new_n278_), .C1(new_n300_), .C2(new_n304_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n282_), .B1(new_n301_), .B2(new_n297_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n298_), .A2(new_n302_), .A3(new_n299_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n278_), .A2(KEYINPUT69), .ZN(new_n308_));
  OR2_X1    g107(.A1(new_n278_), .A2(KEYINPUT69), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n306_), .A2(new_n307_), .A3(new_n308_), .A4(new_n309_), .ZN(new_n310_));
  AND2_X1   g109(.A1(new_n305_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G231gat), .A2(G233gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT71), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n208_), .B(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G1gat), .B(G8gat), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT70), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(G15gat), .ZN(new_n319_));
  INV_X1    g118(.A(G22gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G15gat), .A2(G22gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G1gat), .A2(G8gat), .ZN(new_n323_));
  AOI22_X1  g122(.A1(new_n321_), .A2(new_n322_), .B1(KEYINPUT14), .B2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n318_), .B(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n315_), .B(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT17), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G127gat), .B(G155gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT16), .ZN(new_n329_));
  XOR2_X1   g128(.A(G183gat), .B(G211gat), .Z(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  NOR3_X1   g130(.A1(new_n326_), .A2(new_n327_), .A3(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(KEYINPUT17), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n332_), .B1(new_n326_), .B2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n312_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n277_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT72), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT81), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G127gat), .B(G134gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G113gat), .B(G120gat), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n340_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  XOR2_X1   g142(.A(G127gat), .B(G134gat), .Z(new_n344_));
  INV_X1    g143(.A(G120gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(G113gat), .ZN(new_n346_));
  INV_X1    g145(.A(G113gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(G120gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n344_), .A2(KEYINPUT81), .A3(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT80), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n341_), .A2(new_n342_), .A3(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n351_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n354_));
  OAI211_X1 g153(.A(new_n343_), .B(new_n350_), .C1(new_n353_), .C2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G227gat), .A2(G233gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(new_n319_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G71gat), .B(G99gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(G43gat), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n359_), .A2(G43gat), .ZN(new_n362_));
  NOR3_X1   g161(.A1(new_n361_), .A2(KEYINPUT30), .A3(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT30), .ZN(new_n364_));
  OR2_X1    g163(.A1(new_n359_), .A2(G43gat), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n364_), .B1(new_n365_), .B2(new_n360_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n358_), .B1(new_n363_), .B2(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(KEYINPUT30), .B1(new_n361_), .B2(new_n362_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n365_), .A2(new_n364_), .A3(new_n360_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n368_), .A2(new_n357_), .A3(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n367_), .A2(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(G183gat), .ZN(new_n374_));
  INV_X1    g173(.A(G190gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n373_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G169gat), .A2(G176gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT79), .B(G176gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(KEYINPUT78), .A2(KEYINPUT22), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(G169gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n381_), .A2(G169gat), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n378_), .B(new_n379_), .C1(new_n383_), .C2(new_n384_), .ZN(new_n385_));
  NOR3_X1   g184(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n386_));
  AND3_X1   g185(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n387_));
  NOR3_X1   g186(.A1(new_n386_), .A2(new_n387_), .A3(new_n372_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n379_), .A2(KEYINPUT24), .ZN(new_n389_));
  NOR2_X1   g188(.A1(G169gat), .A2(G176gat), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT76), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(G169gat), .ZN(new_n392_));
  INV_X1    g191(.A(G176gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT76), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n394_), .A2(new_n395_), .A3(KEYINPUT24), .A4(new_n379_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT25), .B(G183gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT26), .B(G190gat), .ZN(new_n398_));
  AOI22_X1  g197(.A1(new_n391_), .A2(new_n396_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT77), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n388_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n391_), .A2(new_n396_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n374_), .A2(KEYINPUT25), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT25), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(G183gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n375_), .A2(KEYINPUT26), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT26), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(G190gat), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n403_), .A2(new_n405_), .A3(new_n406_), .A4(new_n408_), .ZN(new_n409_));
  AND3_X1   g208(.A1(new_n402_), .A2(new_n400_), .A3(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n385_), .B1(new_n401_), .B2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n371_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT82), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n414_), .B1(new_n371_), .B2(new_n411_), .ZN(new_n415_));
  OAI21_X1  g214(.A(KEYINPUT83), .B1(new_n413_), .B2(new_n415_), .ZN(new_n416_));
  OR2_X1    g215(.A1(new_n371_), .A2(new_n411_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT83), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n417_), .A2(new_n414_), .A3(new_n418_), .A4(new_n412_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT31), .ZN(new_n420_));
  AND3_X1   g219(.A1(new_n416_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n420_), .B1(new_n416_), .B2(new_n419_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n355_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n416_), .A2(new_n419_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(KEYINPUT31), .ZN(new_n425_));
  INV_X1    g224(.A(new_n355_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n416_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n425_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n428_));
  AND2_X1   g227(.A1(new_n423_), .A2(new_n428_), .ZN(new_n429_));
  OR2_X1    g228(.A1(G197gat), .A2(G204gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(G197gat), .A2(G204gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT21), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n430_), .A2(KEYINPUT21), .A3(new_n431_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G211gat), .B(G218gat), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n434_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  OR2_X1    g236(.A1(new_n435_), .A2(new_n436_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n411_), .A2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(KEYINPUT19), .A2(G226gat), .A3(G233gat), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(KEYINPUT19), .B1(G226gat), .B2(G233gat), .ZN(new_n443_));
  OR2_X1    g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT20), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(KEYINPUT22), .B(G169gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n380_), .A2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n449_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT90), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT24), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n452_), .B1(G169gat), .B2(G176gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n394_), .ZN(new_n454_));
  AND4_X1   g253(.A1(new_n451_), .A2(new_n388_), .A3(new_n409_), .A4(new_n454_), .ZN(new_n455_));
  AOI22_X1  g254(.A1(new_n397_), .A2(new_n398_), .B1(new_n453_), .B2(new_n394_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n451_), .B1(new_n456_), .B2(new_n388_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n450_), .B1(new_n455_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT91), .ZN(new_n459_));
  NOR3_X1   g258(.A1(new_n458_), .A2(new_n459_), .A3(new_n439_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n450_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n388_), .A2(new_n409_), .A3(new_n454_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT90), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n456_), .A2(new_n451_), .A3(new_n388_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n461_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n437_), .A2(new_n438_), .ZN(new_n466_));
  AOI21_X1  g265(.A(KEYINPUT91), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  OAI211_X1 g266(.A(new_n440_), .B(new_n447_), .C1(new_n460_), .C2(new_n467_), .ZN(new_n468_));
  XOR2_X1   g267(.A(G8gat), .B(G36gat), .Z(new_n469_));
  XNOR2_X1  g268(.A(new_n469_), .B(KEYINPUT18), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G64gat), .B(G92gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n470_), .B(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n444_), .B(KEYINPUT89), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT20), .B1(new_n465_), .B2(new_n466_), .ZN(new_n474_));
  OAI211_X1 g273(.A(new_n385_), .B(new_n466_), .C1(new_n401_), .C2(new_n410_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n473_), .B1(new_n474_), .B2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n468_), .A2(new_n472_), .A3(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT27), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n472_), .B(KEYINPUT96), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n458_), .A2(new_n439_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n473_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n482_), .A2(KEYINPUT20), .A3(new_n475_), .A4(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT95), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n446_), .B1(new_n458_), .B2(new_n439_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT95), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n486_), .A2(new_n487_), .A3(new_n475_), .A4(new_n483_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n485_), .A2(new_n488_), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n462_), .A2(new_n450_), .A3(new_n437_), .A4(new_n438_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(KEYINPUT20), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n491_), .B1(new_n411_), .B2(new_n439_), .ZN(new_n492_));
  OAI21_X1  g291(.A(KEYINPUT94), .B1(new_n492_), .B2(new_n444_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT94), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n395_), .B1(new_n453_), .B2(new_n394_), .ZN(new_n495_));
  NOR3_X1   g294(.A1(new_n389_), .A2(KEYINPUT76), .A3(new_n390_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n409_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(KEYINPUT77), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n399_), .A2(new_n400_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n498_), .A2(new_n499_), .A3(new_n388_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n466_), .B1(new_n500_), .B2(new_n385_), .ZN(new_n501_));
  OAI211_X1 g300(.A(new_n494_), .B(new_n445_), .C1(new_n501_), .C2(new_n491_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n493_), .A2(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n481_), .B1(new_n489_), .B2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT97), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n479_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  AOI22_X1  g305(.A1(new_n485_), .A2(new_n488_), .B1(new_n493_), .B2(new_n502_), .ZN(new_n507_));
  OAI21_X1  g306(.A(KEYINPUT97), .B1(new_n507_), .B2(new_n481_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT27), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n468_), .A2(new_n477_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n472_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(new_n478_), .ZN(new_n513_));
  AOI22_X1  g312(.A1(new_n506_), .A2(new_n508_), .B1(new_n509_), .B2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT84), .ZN(new_n515_));
  INV_X1    g314(.A(G155gat), .ZN(new_n516_));
  INV_X1    g315(.A(G162gat), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n515_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT84), .B1(G155gat), .B2(G162gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G155gat), .A2(G162gat), .ZN(new_n520_));
  AND3_X1   g319(.A1(new_n518_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(G141gat), .A2(G148gat), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT3), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G141gat), .A2(G148gat), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT2), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n528_));
  OAI21_X1  g327(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n524_), .A2(new_n527_), .A3(new_n528_), .A4(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n521_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n520_), .A2(KEYINPUT1), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT1), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n533_), .A2(G155gat), .A3(G162gat), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n518_), .A2(new_n532_), .A3(new_n534_), .A4(new_n519_), .ZN(new_n535_));
  XOR2_X1   g334(.A(G141gat), .B(G148gat), .Z(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n531_), .A2(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(KEYINPUT28), .B1(new_n538_), .B2(KEYINPUT29), .ZN(new_n539_));
  AOI22_X1  g338(.A1(new_n521_), .A2(new_n530_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT28), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT29), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n540_), .A2(new_n541_), .A3(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n539_), .A2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G22gat), .B(G50gat), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n544_), .B(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT88), .ZN(new_n548_));
  AND2_X1   g347(.A1(G228gat), .A2(G233gat), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n549_), .B1(new_n439_), .B2(KEYINPUT85), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n439_), .B1(new_n540_), .B2(new_n542_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  OAI221_X1 g351(.A(new_n439_), .B1(KEYINPUT85), .B2(new_n549_), .C1(new_n540_), .C2(new_n542_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G78gat), .B(G106gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT86), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n554_), .A2(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n547_), .B1(new_n548_), .B2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n552_), .A2(new_n553_), .A3(new_n555_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT87), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n557_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(KEYINPUT88), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n558_), .A2(new_n561_), .A3(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n554_), .A2(new_n556_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n547_), .B1(new_n562_), .B2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G1gat), .B(G29gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(G85gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(KEYINPUT0), .B(G57gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n344_), .A2(new_n349_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n341_), .A2(new_n342_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n540_), .A2(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n576_), .B1(new_n355_), .B2(new_n540_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(KEYINPUT4), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G225gat), .A2(G233gat), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n579_), .B(KEYINPUT92), .Z(new_n580_));
  NAND2_X1  g379(.A1(new_n574_), .A2(KEYINPUT80), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(new_n352_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n538_), .A2(new_n582_), .A3(new_n343_), .A4(new_n350_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT4), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n578_), .A2(new_n580_), .A3(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n580_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n577_), .A2(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n572_), .B1(new_n586_), .B2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n586_), .A2(new_n572_), .A3(new_n588_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n429_), .A2(new_n514_), .A3(new_n568_), .A4(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n489_), .A2(new_n503_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n595_), .A2(new_n505_), .A3(new_n480_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n479_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n508_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n513_), .A2(new_n509_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n592_), .B1(new_n564_), .B2(new_n566_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n598_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n572_), .B1(new_n577_), .B2(new_n587_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n578_), .A2(new_n585_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n602_), .B1(new_n603_), .B2(new_n587_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT93), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n605_), .A2(KEYINPUT33), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n604_), .B1(new_n589_), .B2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n588_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n584_), .B1(new_n583_), .B2(new_n576_), .ZN(new_n610_));
  AOI21_X1  g409(.A(KEYINPUT4), .B1(new_n426_), .B2(new_n538_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n609_), .B1(new_n612_), .B2(new_n580_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n606_), .B1(new_n613_), .B2(new_n572_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n608_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n472_), .A2(KEYINPUT32), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n616_), .B1(new_n489_), .B2(new_n503_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n468_), .A2(new_n616_), .A3(new_n477_), .ZN(new_n618_));
  AND3_X1   g417(.A1(new_n586_), .A2(new_n572_), .A3(new_n588_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n618_), .B1(new_n619_), .B2(new_n589_), .ZN(new_n620_));
  OAI22_X1  g419(.A1(new_n615_), .A2(new_n513_), .B1(new_n617_), .B2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(new_n568_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n429_), .B1(new_n601_), .B2(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n594_), .B1(new_n623_), .B2(KEYINPUT98), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT98), .ZN(new_n625_));
  AOI211_X1 g424(.A(new_n625_), .B(new_n429_), .C1(new_n601_), .C2(new_n622_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n624_), .A2(new_n626_), .ZN(new_n627_));
  XOR2_X1   g426(.A(G113gat), .B(G141gat), .Z(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT73), .ZN(new_n629_));
  XNOR2_X1  g428(.A(G169gat), .B(G197gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n325_), .B(new_n286_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(G229gat), .A2(G233gat), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n325_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(new_n287_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n325_), .A2(new_n286_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n638_), .A2(new_n639_), .A3(new_n634_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n636_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT74), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n632_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  AOI211_X1 g442(.A(KEYINPUT74), .B(new_n631_), .C1(new_n636_), .C2(new_n640_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(KEYINPUT75), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT75), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n645_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n627_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n277_), .A2(KEYINPUT72), .A3(new_n336_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n339_), .A2(new_n652_), .A3(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(KEYINPUT99), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT99), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n339_), .A2(new_n656_), .A3(new_n652_), .A4(new_n653_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n593_), .A2(G1gat), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n655_), .A2(new_n657_), .A3(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT38), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n300_), .A2(new_n304_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n627_), .A2(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n663_), .A2(KEYINPUT100), .ZN(new_n664_));
  AOI22_X1  g463(.A1(new_n514_), .A2(new_n600_), .B1(new_n568_), .B2(new_n621_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n625_), .B1(new_n665_), .B2(new_n429_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n623_), .A2(KEYINPUT98), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n666_), .A2(new_n667_), .A3(new_n594_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n662_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n668_), .A2(KEYINPUT100), .A3(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n664_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n277_), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n673_), .A2(new_n646_), .A3(new_n335_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n672_), .A2(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(G1gat), .B1(new_n675_), .B2(new_n593_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n659_), .A2(new_n660_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n661_), .A2(new_n676_), .A3(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT101), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n661_), .A2(KEYINPUT101), .A3(new_n676_), .A4(new_n677_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(G1324gat));
  XNOR2_X1  g481(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT39), .ZN(new_n684_));
  INV_X1    g483(.A(new_n514_), .ZN(new_n685_));
  OAI211_X1 g484(.A(new_n685_), .B(new_n674_), .C1(new_n664_), .C2(new_n671_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n684_), .B1(new_n686_), .B2(G8gat), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n686_), .A2(new_n684_), .A3(G8gat), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n514_), .A2(G8gat), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n655_), .A2(new_n657_), .A3(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n683_), .B1(new_n690_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n689_), .ZN(new_n694_));
  OAI211_X1 g493(.A(new_n692_), .B(new_n683_), .C1(new_n694_), .C2(new_n687_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n693_), .A2(new_n696_), .ZN(G1325gat));
  INV_X1    g496(.A(new_n654_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n698_), .A2(new_n319_), .A3(new_n429_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n675_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(new_n429_), .ZN(new_n701_));
  AND3_X1   g500(.A1(new_n701_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n702_));
  AOI21_X1  g501(.A(KEYINPUT41), .B1(new_n701_), .B2(G15gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n699_), .B1(new_n702_), .B2(new_n703_), .ZN(G1326gat));
  NAND3_X1  g503(.A1(new_n698_), .A2(new_n320_), .A3(new_n567_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT42), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n700_), .A2(new_n567_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n707_), .B2(G22gat), .ZN(new_n708_));
  AOI211_X1 g507(.A(KEYINPUT42), .B(new_n320_), .C1(new_n700_), .C2(new_n567_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n705_), .B1(new_n708_), .B2(new_n709_), .ZN(G1327gat));
  NOR2_X1   g509(.A1(new_n669_), .A2(new_n334_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n277_), .A2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(new_n652_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(G29gat), .B1(new_n714_), .B2(new_n592_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n673_), .A2(new_n646_), .A3(new_n334_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n312_), .B1(new_n624_), .B2(new_n626_), .ZN(new_n717_));
  XOR2_X1   g516(.A(KEYINPUT103), .B(KEYINPUT43), .Z(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n717_), .A2(KEYINPUT104), .A3(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(KEYINPUT104), .B1(new_n717_), .B2(new_n719_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT43), .ZN(new_n723_));
  OAI211_X1 g522(.A(new_n723_), .B(new_n312_), .C1(new_n624_), .C2(new_n626_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT105), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n668_), .A2(KEYINPUT105), .A3(new_n723_), .A4(new_n312_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  OAI211_X1 g527(.A(new_n716_), .B(KEYINPUT44), .C1(new_n722_), .C2(new_n728_), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n729_), .A2(G29gat), .A3(new_n592_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n717_), .A2(new_n719_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT104), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n717_), .A2(KEYINPUT104), .A3(new_n719_), .ZN(new_n735_));
  AOI22_X1  g534(.A1(new_n734_), .A2(new_n735_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n716_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n731_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n715_), .B1(new_n730_), .B2(new_n738_), .ZN(G1328gat));
  INV_X1    g538(.A(KEYINPUT107), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n740_), .A2(KEYINPUT46), .ZN(new_n741_));
  INV_X1    g540(.A(G36gat), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n734_), .A2(new_n735_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n726_), .A2(new_n727_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n737_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n514_), .B1(new_n745_), .B2(KEYINPUT44), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n742_), .B1(new_n746_), .B2(new_n738_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n714_), .A2(new_n742_), .A3(new_n685_), .ZN(new_n748_));
  XOR2_X1   g547(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n749_));
  XOR2_X1   g548(.A(new_n748_), .B(new_n749_), .Z(new_n750_));
  OAI21_X1  g549(.A(new_n741_), .B1(new_n747_), .B2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n738_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n729_), .A2(new_n685_), .ZN(new_n753_));
  OAI21_X1  g552(.A(G36gat), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n741_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n748_), .B(new_n749_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n754_), .A2(new_n755_), .A3(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n751_), .A2(new_n757_), .ZN(G1329gat));
  NAND4_X1  g557(.A1(new_n738_), .A2(G43gat), .A3(new_n729_), .A4(new_n429_), .ZN(new_n759_));
  INV_X1    g558(.A(G43gat), .ZN(new_n760_));
  INV_X1    g559(.A(new_n429_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n760_), .B1(new_n713_), .B2(new_n761_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n763_));
  AND3_X1   g562(.A1(new_n759_), .A2(new_n762_), .A3(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n759_), .B2(new_n762_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n764_), .A2(new_n765_), .ZN(G1330gat));
  OR3_X1    g565(.A1(new_n713_), .A2(G50gat), .A3(new_n568_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n738_), .A2(new_n567_), .A3(new_n729_), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n768_), .A2(KEYINPUT109), .A3(G50gat), .ZN(new_n769_));
  AOI21_X1  g568(.A(KEYINPUT109), .B1(new_n768_), .B2(G50gat), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n767_), .B1(new_n769_), .B2(new_n770_), .ZN(G1331gat));
  NAND3_X1  g570(.A1(new_n647_), .A2(new_n649_), .A3(new_n334_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n672_), .A2(KEYINPUT110), .A3(new_n673_), .A4(new_n773_), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n673_), .B(new_n773_), .C1(new_n664_), .C2(new_n671_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT110), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n592_), .A2(G57gat), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n774_), .A2(new_n777_), .A3(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT111), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n779_), .A2(new_n780_), .ZN(new_n782_));
  NOR3_X1   g581(.A1(new_n627_), .A2(new_n277_), .A3(new_n645_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n336_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(G57gat), .B1(new_n785_), .B2(new_n592_), .ZN(new_n786_));
  NOR3_X1   g585(.A1(new_n781_), .A2(new_n782_), .A3(new_n786_), .ZN(G1332gat));
  OR3_X1    g586(.A1(new_n784_), .A2(G64gat), .A3(new_n514_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n774_), .A2(new_n777_), .A3(new_n685_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT48), .ZN(new_n790_));
  AND3_X1   g589(.A1(new_n789_), .A2(new_n790_), .A3(G64gat), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n789_), .B2(G64gat), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n788_), .B1(new_n791_), .B2(new_n792_), .ZN(G1333gat));
  NAND3_X1  g592(.A1(new_n774_), .A2(new_n777_), .A3(new_n429_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT49), .ZN(new_n795_));
  AND3_X1   g594(.A1(new_n794_), .A2(new_n795_), .A3(G71gat), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n795_), .B1(new_n794_), .B2(G71gat), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n761_), .A2(G71gat), .ZN(new_n798_));
  XOR2_X1   g597(.A(new_n798_), .B(KEYINPUT112), .Z(new_n799_));
  OAI22_X1  g598(.A1(new_n796_), .A2(new_n797_), .B1(new_n784_), .B2(new_n799_), .ZN(G1334gat));
  OR3_X1    g599(.A1(new_n784_), .A2(G78gat), .A3(new_n568_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n774_), .A2(new_n777_), .A3(new_n567_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT50), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n802_), .A2(new_n803_), .A3(G78gat), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n803_), .B1(new_n802_), .B2(G78gat), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n801_), .B1(new_n804_), .B2(new_n805_), .ZN(G1335gat));
  NAND2_X1  g605(.A1(new_n783_), .A2(new_n711_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n808_), .A2(new_n223_), .A3(new_n592_), .ZN(new_n809_));
  NOR3_X1   g608(.A1(new_n277_), .A2(new_n645_), .A3(new_n334_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  NOR3_X1   g610(.A1(new_n736_), .A2(new_n593_), .A3(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n809_), .B1(new_n812_), .B2(new_n223_), .ZN(G1336gat));
  NAND3_X1  g612(.A1(new_n808_), .A2(new_n224_), .A3(new_n685_), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n736_), .A2(new_n514_), .A3(new_n811_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n814_), .B1(new_n815_), .B2(new_n224_), .ZN(G1337gat));
  INV_X1    g615(.A(KEYINPUT113), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n783_), .A2(new_n429_), .A3(new_n242_), .A4(new_n711_), .ZN(new_n818_));
  NOR3_X1   g617(.A1(new_n736_), .A2(new_n761_), .A3(new_n811_), .ZN(new_n819_));
  INV_X1    g618(.A(G99gat), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n817_), .B(new_n818_), .C1(new_n819_), .C2(new_n820_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g621(.A1(new_n808_), .A2(new_n241_), .A3(new_n567_), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n567_), .B(new_n810_), .C1(new_n722_), .C2(new_n728_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n824_), .A2(new_n825_), .A3(G106gat), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n825_), .B1(new_n824_), .B2(G106gat), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n823_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT53), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n830_), .B(new_n823_), .C1(new_n826_), .C2(new_n827_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n829_), .A2(new_n831_), .ZN(G1339gat));
  INV_X1    g631(.A(KEYINPUT114), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n772_), .A2(new_n833_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n647_), .A2(KEYINPUT114), .A3(new_n649_), .A4(new_n334_), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n836_), .A2(new_n274_), .A3(new_n311_), .A4(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n837_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n834_), .A2(new_n274_), .A3(new_n835_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n839_), .B1(new_n840_), .B2(new_n312_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n838_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT56), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n252_), .A2(new_n260_), .A3(new_n255_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n258_), .A2(KEYINPUT55), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT55), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n256_), .A2(new_n847_), .A3(new_n257_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n845_), .B1(new_n846_), .B2(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n843_), .B1(new_n849_), .B2(new_n269_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT116), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n847_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n852_));
  AOI211_X1 g651(.A(KEYINPUT55), .B(new_n260_), .C1(new_n252_), .C2(new_n255_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n844_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n854_), .A2(KEYINPUT56), .A3(new_n267_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n850_), .A2(new_n851_), .A3(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n645_), .A2(new_n270_), .ZN(new_n857_));
  AOI21_X1  g656(.A(KEYINPUT56), .B1(new_n854_), .B2(new_n267_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n857_), .B1(new_n858_), .B2(KEYINPUT116), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n856_), .A2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n268_), .A2(new_n270_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n641_), .A2(new_n631_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n633_), .A2(new_n634_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n638_), .A2(new_n639_), .A3(new_n635_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n863_), .A2(new_n631_), .A3(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT117), .ZN(new_n866_));
  OR2_X1    g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n865_), .A2(new_n866_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n862_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n861_), .A2(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n662_), .B1(new_n860_), .B2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n270_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n872_), .B1(new_n850_), .B2(new_n855_), .ZN(new_n873_));
  OR2_X1    g672(.A1(new_n873_), .A2(KEYINPUT58), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n311_), .B1(new_n873_), .B2(KEYINPUT58), .ZN(new_n875_));
  AOI22_X1  g674(.A1(new_n871_), .A2(KEYINPUT57), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n877_), .B1(new_n871_), .B2(KEYINPUT57), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT57), .ZN(new_n879_));
  AOI22_X1  g678(.A1(new_n856_), .A2(new_n859_), .B1(new_n861_), .B2(new_n869_), .ZN(new_n880_));
  OAI211_X1 g679(.A(KEYINPUT118), .B(new_n879_), .C1(new_n880_), .C2(new_n662_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n876_), .A2(new_n878_), .A3(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n842_), .B1(new_n882_), .B2(new_n335_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n761_), .A2(new_n593_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n685_), .A2(new_n567_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n883_), .A2(new_n886_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n887_), .A2(new_n347_), .A3(new_n645_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n886_), .ZN(new_n889_));
  AOI21_X1  g688(.A(KEYINPUT59), .B1(new_n889_), .B2(KEYINPUT120), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n890_), .B1(KEYINPUT120), .B2(new_n889_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n879_), .B1(new_n880_), .B2(new_n662_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n874_), .A2(new_n875_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n892_), .A2(new_n893_), .A3(KEYINPUT121), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n871_), .A2(KEYINPUT57), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(KEYINPUT121), .B1(new_n892_), .B2(new_n893_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n335_), .B1(new_n896_), .B2(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n842_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n891_), .B1(new_n898_), .B2(new_n899_), .ZN(new_n900_));
  OAI21_X1  g699(.A(KEYINPUT59), .B1(new_n883_), .B2(new_n886_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT119), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  OAI211_X1 g702(.A(KEYINPUT119), .B(KEYINPUT59), .C1(new_n883_), .C2(new_n886_), .ZN(new_n904_));
  AOI211_X1 g703(.A(new_n651_), .B(new_n900_), .C1(new_n903_), .C2(new_n904_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n888_), .B1(new_n905_), .B2(new_n347_), .ZN(G1340gat));
  OAI21_X1  g705(.A(new_n345_), .B1(new_n277_), .B2(KEYINPUT60), .ZN(new_n907_));
  OAI211_X1 g706(.A(new_n887_), .B(new_n907_), .C1(KEYINPUT60), .C2(new_n345_), .ZN(new_n908_));
  AOI211_X1 g707(.A(new_n277_), .B(new_n900_), .C1(new_n903_), .C2(new_n904_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n909_), .B2(new_n345_), .ZN(G1341gat));
  INV_X1    g709(.A(G127gat), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n887_), .A2(new_n911_), .A3(new_n334_), .ZN(new_n912_));
  AOI211_X1 g711(.A(new_n335_), .B(new_n900_), .C1(new_n903_), .C2(new_n904_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n913_), .B2(new_n911_), .ZN(G1342gat));
  NAND2_X1  g713(.A1(new_n887_), .A2(new_n662_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT122), .ZN(new_n916_));
  INV_X1    g715(.A(G134gat), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n915_), .A2(new_n916_), .A3(new_n917_), .ZN(new_n918_));
  NOR3_X1   g717(.A1(new_n883_), .A2(new_n669_), .A3(new_n886_), .ZN(new_n919_));
  OAI21_X1  g718(.A(KEYINPUT122), .B1(new_n919_), .B2(G134gat), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n918_), .A2(new_n920_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n900_), .B1(new_n903_), .B2(new_n904_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n311_), .A2(new_n917_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n921_), .B1(new_n922_), .B2(new_n923_), .ZN(G1343gat));
  NOR4_X1   g723(.A1(new_n685_), .A2(new_n429_), .A3(new_n568_), .A4(new_n593_), .ZN(new_n925_));
  INV_X1    g724(.A(new_n925_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n883_), .A2(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(new_n645_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g728(.A1(new_n927_), .A2(new_n673_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g730(.A1(new_n882_), .A2(new_n335_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(new_n899_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(new_n925_), .ZN(new_n934_));
  OAI21_X1  g733(.A(KEYINPUT123), .B1(new_n934_), .B2(new_n335_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT123), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n927_), .A2(new_n936_), .A3(new_n334_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(KEYINPUT61), .B(G155gat), .ZN(new_n938_));
  AND3_X1   g737(.A1(new_n935_), .A2(new_n937_), .A3(new_n938_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n938_), .B1(new_n935_), .B2(new_n937_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n939_), .A2(new_n940_), .ZN(G1346gat));
  OAI21_X1  g740(.A(G162gat), .B1(new_n934_), .B2(new_n311_), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n927_), .A2(new_n517_), .A3(new_n662_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n942_), .A2(new_n943_), .ZN(G1347gat));
  INV_X1    g743(.A(KEYINPUT62), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n898_), .A2(new_n899_), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n685_), .A2(new_n429_), .A3(new_n593_), .ZN(new_n947_));
  XNOR2_X1  g746(.A(new_n947_), .B(KEYINPUT124), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n948_), .A2(new_n567_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n946_), .A2(new_n949_), .ZN(new_n950_));
  NOR2_X1   g749(.A1(new_n950_), .A2(new_n646_), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n945_), .B1(new_n951_), .B2(new_n392_), .ZN(new_n952_));
  OAI211_X1 g751(.A(KEYINPUT62), .B(G169gat), .C1(new_n950_), .C2(new_n646_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n951_), .A2(new_n448_), .ZN(new_n954_));
  NAND3_X1  g753(.A1(new_n952_), .A2(new_n953_), .A3(new_n954_), .ZN(G1348gat));
  INV_X1    g754(.A(new_n950_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n956_), .A2(new_n673_), .ZN(new_n957_));
  NOR2_X1   g756(.A1(new_n883_), .A2(new_n567_), .ZN(new_n958_));
  NOR3_X1   g757(.A1(new_n948_), .A2(new_n277_), .A3(new_n393_), .ZN(new_n959_));
  AOI22_X1  g758(.A1(new_n957_), .A2(new_n380_), .B1(new_n958_), .B2(new_n959_), .ZN(G1349gat));
  NOR3_X1   g759(.A1(new_n950_), .A2(new_n397_), .A3(new_n335_), .ZN(new_n961_));
  INV_X1    g760(.A(new_n948_), .ZN(new_n962_));
  NAND3_X1  g761(.A1(new_n958_), .A2(new_n334_), .A3(new_n962_), .ZN(new_n963_));
  AOI21_X1  g762(.A(new_n961_), .B1(new_n374_), .B2(new_n963_), .ZN(G1350gat));
  OAI21_X1  g763(.A(G190gat), .B1(new_n950_), .B2(new_n311_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n662_), .A2(new_n398_), .ZN(new_n966_));
  OAI21_X1  g765(.A(new_n965_), .B1(new_n950_), .B2(new_n966_), .ZN(G1351gat));
  INV_X1    g766(.A(KEYINPUT125), .ZN(new_n968_));
  NOR3_X1   g767(.A1(new_n429_), .A2(new_n568_), .A3(new_n592_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n969_), .A2(new_n685_), .ZN(new_n970_));
  INV_X1    g769(.A(new_n970_), .ZN(new_n971_));
  NAND3_X1  g770(.A1(new_n933_), .A2(new_n968_), .A3(new_n971_), .ZN(new_n972_));
  OAI21_X1  g771(.A(KEYINPUT125), .B1(new_n883_), .B2(new_n970_), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n972_), .A2(new_n973_), .ZN(new_n974_));
  NAND2_X1  g773(.A1(new_n974_), .A2(new_n645_), .ZN(new_n975_));
  XNOR2_X1  g774(.A(new_n975_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g775(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n977_));
  NAND3_X1  g776(.A1(new_n974_), .A2(new_n673_), .A3(new_n977_), .ZN(new_n978_));
  INV_X1    g777(.A(new_n974_), .ZN(new_n979_));
  NOR2_X1   g778(.A1(new_n979_), .A2(new_n277_), .ZN(new_n980_));
  XOR2_X1   g779(.A(KEYINPUT126), .B(G204gat), .Z(new_n981_));
  OAI21_X1  g780(.A(new_n978_), .B1(new_n980_), .B2(new_n981_), .ZN(G1353gat));
  AOI211_X1 g781(.A(KEYINPUT63), .B(G211gat), .C1(new_n974_), .C2(new_n334_), .ZN(new_n983_));
  XNOR2_X1  g782(.A(KEYINPUT63), .B(G211gat), .ZN(new_n984_));
  AOI211_X1 g783(.A(new_n335_), .B(new_n984_), .C1(new_n972_), .C2(new_n973_), .ZN(new_n985_));
  NOR2_X1   g784(.A1(new_n983_), .A2(new_n985_), .ZN(G1354gat));
  OAI21_X1  g785(.A(G218gat), .B1(new_n979_), .B2(new_n311_), .ZN(new_n987_));
  INV_X1    g786(.A(G218gat), .ZN(new_n988_));
  NAND3_X1  g787(.A1(new_n974_), .A2(new_n988_), .A3(new_n662_), .ZN(new_n989_));
  NAND2_X1  g788(.A1(new_n987_), .A2(new_n989_), .ZN(G1355gat));
endmodule


