//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 1 0 1 1 0 1 1 0 1 0 0 0 0 1 1 1 1 0 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 0 1 1 1 0 0 0 0 1 0 1 0 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n754_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n774_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n791_, new_n792_, new_n793_, new_n795_, new_n796_, new_n797_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n903_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n910_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n926_, new_n927_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n934_, new_n935_, new_n936_,
    new_n937_, new_n938_, new_n940_, new_n941_, new_n943_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n950_, new_n951_;
  OR2_X1    g000(.A1(G211gat), .A2(G218gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G211gat), .A2(G218gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  OR2_X1    g003(.A1(new_n204_), .A2(KEYINPUT86), .ZN(new_n205_));
  INV_X1    g004(.A(G204gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(G197gat), .ZN(new_n207_));
  INV_X1    g006(.A(G197gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(G204gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n207_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n204_), .A2(KEYINPUT86), .ZN(new_n211_));
  NAND4_X1  g010(.A1(new_n205_), .A2(KEYINPUT21), .A3(new_n210_), .A4(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT85), .ZN(new_n213_));
  AOI22_X1  g012(.A1(new_n210_), .A2(KEYINPUT21), .B1(new_n202_), .B2(new_n203_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT21), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n207_), .A2(new_n209_), .A3(new_n215_), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n213_), .B1(new_n214_), .B2(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n208_), .A2(G204gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n206_), .A2(G197gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT21), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  AND4_X1   g019(.A1(new_n213_), .A2(new_n220_), .A3(new_n204_), .A4(new_n216_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n212_), .B1(new_n217_), .B2(new_n221_), .ZN(new_n222_));
  OR2_X1    g021(.A1(G155gat), .A2(G162gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G155gat), .A2(G162gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n225_));
  INV_X1    g024(.A(G141gat), .ZN(new_n226_));
  INV_X1    g025(.A(G148gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT2), .ZN(new_n230_));
  AOI21_X1  g029(.A(KEYINPUT82), .B1(G141gat), .B2(G148gat), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n228_), .B(new_n229_), .C1(new_n230_), .C2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n230_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n223_), .B(new_n224_), .C1(new_n232_), .C2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n224_), .A2(KEYINPUT1), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n236_), .A2(new_n223_), .A3(KEYINPUT81), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(KEYINPUT81), .B1(new_n236_), .B2(new_n223_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n224_), .A2(KEYINPUT1), .ZN(new_n240_));
  NOR3_X1   g039(.A1(new_n238_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G141gat), .B(G148gat), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n235_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT29), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n222_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G228gat), .A2(G233gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT84), .ZN(new_n248_));
  OR2_X1    g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n246_), .A2(G228gat), .A3(G233gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT87), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT87), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n249_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n244_), .A2(new_n245_), .ZN(new_n255_));
  XOR2_X1   g054(.A(G22gat), .B(G50gat), .Z(new_n256_));
  XNOR2_X1  g055(.A(new_n255_), .B(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  AND3_X1   g057(.A1(new_n252_), .A2(new_n254_), .A3(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n258_), .B1(new_n252_), .B2(new_n254_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G78gat), .B(G106gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT88), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT83), .B(KEYINPUT28), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  OR3_X1    g064(.A1(new_n259_), .A2(new_n260_), .A3(new_n265_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n265_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G127gat), .A2(G134gat), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(G127gat), .A2(G134gat), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  AND2_X1   g072(.A1(G113gat), .A2(G120gat), .ZN(new_n274_));
  NOR2_X1   g073(.A1(G113gat), .A2(G120gat), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(KEYINPUT80), .B1(new_n273_), .B2(new_n276_), .ZN(new_n277_));
  OAI22_X1  g076(.A1(new_n272_), .A2(new_n271_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n275_), .ZN(new_n279_));
  INV_X1    g078(.A(G127gat), .ZN(new_n280_));
  INV_X1    g079(.A(G134gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G113gat), .A2(G120gat), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n279_), .A2(new_n282_), .A3(new_n270_), .A4(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n278_), .A2(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n277_), .B1(new_n285_), .B2(KEYINPUT80), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT31), .ZN(new_n287_));
  OR2_X1    g086(.A1(new_n287_), .A2(KEYINPUT79), .ZN(new_n288_));
  AND2_X1   g087(.A1(new_n288_), .A2(G43gat), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n288_), .A2(G43gat), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G227gat), .A2(G233gat), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n291_), .B(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT23), .ZN(new_n295_));
  AND3_X1   g094(.A1(KEYINPUT76), .A2(G183gat), .A3(G190gat), .ZN(new_n296_));
  AOI21_X1  g095(.A(KEYINPUT76), .B1(G183gat), .B2(G190gat), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n295_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G183gat), .A2(G190gat), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n299_), .A2(new_n295_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT24), .ZN(new_n302_));
  INV_X1    g101(.A(G169gat), .ZN(new_n303_));
  INV_X1    g102(.A(G176gat), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n302_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n298_), .A2(new_n301_), .A3(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT77), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G169gat), .A2(G176gat), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(G190gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT75), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT75), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(G190gat), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n313_), .A2(new_n315_), .A3(KEYINPUT26), .ZN(new_n316_));
  OR2_X1    g115(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(KEYINPUT25), .B(G183gat), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n311_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT77), .ZN(new_n321_));
  NAND4_X1  g120(.A1(new_n298_), .A2(new_n321_), .A3(new_n301_), .A4(new_n305_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n307_), .A2(new_n320_), .A3(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(KEYINPUT78), .B(G176gat), .ZN(new_n324_));
  XOR2_X1   g123(.A(KEYINPUT22), .B(G169gat), .Z(new_n325_));
  NOR2_X1   g124(.A1(new_n299_), .A2(KEYINPUT23), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT76), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n299_), .A2(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(KEYINPUT76), .A2(G183gat), .A3(G190gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n326_), .B1(new_n330_), .B2(KEYINPUT23), .ZN(new_n331_));
  AOI21_X1  g130(.A(G183gat), .B1(new_n313_), .B2(new_n315_), .ZN(new_n332_));
  OAI221_X1 g131(.A(new_n308_), .B1(new_n324_), .B2(new_n325_), .C1(new_n331_), .C2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n323_), .A2(new_n333_), .ZN(new_n334_));
  XOR2_X1   g133(.A(KEYINPUT30), .B(G15gat), .Z(new_n335_));
  XNOR2_X1  g134(.A(G71gat), .B(G99gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n334_), .B(new_n337_), .ZN(new_n338_));
  AND2_X1   g137(.A1(new_n294_), .A2(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n294_), .A2(new_n338_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G8gat), .B(G36gat), .ZN(new_n342_));
  INV_X1    g141(.A(G92gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT18), .B(G64gat), .ZN(new_n345_));
  XOR2_X1   g144(.A(new_n344_), .B(new_n345_), .Z(new_n346_));
  INV_X1    g145(.A(new_n222_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n305_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n348_));
  OAI21_X1  g147(.A(KEYINPUT23), .B1(new_n296_), .B2(new_n297_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n326_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n348_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n352_));
  AND3_X1   g151(.A1(new_n317_), .A2(KEYINPUT89), .A3(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(KEYINPUT89), .B1(new_n317_), .B2(new_n352_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n319_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT90), .ZN(new_n356_));
  AND3_X1   g155(.A1(new_n351_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n356_), .B1(new_n351_), .B2(new_n355_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(G183gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(new_n312_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n298_), .A2(new_n361_), .A3(new_n301_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT92), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n298_), .A2(KEYINPUT92), .A3(new_n361_), .A4(new_n301_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n308_), .B(KEYINPUT91), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n367_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(KEYINPUT93), .B1(new_n366_), .B2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT93), .ZN(new_n371_));
  AOI211_X1 g170(.A(new_n371_), .B(new_n368_), .C1(new_n364_), .C2(new_n365_), .ZN(new_n372_));
  OAI211_X1 g171(.A(new_n347_), .B(new_n359_), .C1(new_n370_), .C2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT94), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n300_), .B1(new_n330_), .B2(new_n295_), .ZN(new_n376_));
  AOI21_X1  g175(.A(KEYINPUT92), .B1(new_n376_), .B2(new_n361_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n365_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n369_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(new_n371_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n368_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(KEYINPUT93), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n383_), .A2(KEYINPUT94), .A3(new_n347_), .A4(new_n359_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n334_), .A2(new_n222_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G226gat), .A2(G233gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT19), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT20), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n385_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n375_), .A2(new_n384_), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n387_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n359_), .B1(new_n370_), .B2(new_n372_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(new_n222_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n323_), .A2(new_n333_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n388_), .B1(new_n396_), .B2(new_n347_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n393_), .B1(new_n395_), .B2(new_n397_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n346_), .B1(new_n392_), .B2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n351_), .A2(new_n355_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(KEYINPUT90), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n351_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n403_), .B1(new_n380_), .B2(new_n382_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n397_), .B1(new_n404_), .B2(new_n347_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(new_n387_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n375_), .A2(new_n384_), .A3(new_n391_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n346_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n406_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(KEYINPUT27), .B1(new_n399_), .B2(new_n409_), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n400_), .B(new_n212_), .C1(new_n217_), .C2(new_n221_), .ZN(new_n411_));
  OAI21_X1  g210(.A(KEYINPUT20), .B1(new_n411_), .B2(new_n381_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT99), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT99), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n414_), .B(KEYINPUT20), .C1(new_n411_), .C2(new_n381_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n413_), .A2(new_n385_), .A3(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(new_n387_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n395_), .A2(new_n393_), .A3(new_n397_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n417_), .A2(KEYINPUT100), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT100), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n416_), .A2(new_n420_), .A3(new_n387_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n419_), .A2(new_n346_), .A3(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n390_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n423_));
  AOI22_X1  g222(.A1(new_n384_), .A2(new_n423_), .B1(new_n405_), .B2(new_n387_), .ZN(new_n424_));
  AOI21_X1  g223(.A(KEYINPUT103), .B1(new_n424_), .B2(new_n408_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n422_), .A2(new_n425_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n419_), .A2(KEYINPUT103), .A3(new_n346_), .A4(new_n421_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n410_), .B1(new_n428_), .B2(KEYINPUT27), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G225gat), .A2(G233gat), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT4), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n236_), .A2(new_n223_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT81), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n240_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n242_), .B1(new_n435_), .B2(new_n237_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n223_), .A2(new_n224_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n228_), .A2(new_n229_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n231_), .A2(new_n230_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n437_), .B1(new_n440_), .B2(new_n233_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n286_), .B1(new_n436_), .B2(new_n441_), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n235_), .B(new_n285_), .C1(new_n241_), .C2(new_n242_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n432_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(KEYINPUT4), .B1(new_n243_), .B2(new_n286_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n431_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n442_), .A2(new_n443_), .A3(new_n430_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G1gat), .B(G29gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  XOR2_X1   g249(.A(G57gat), .B(G85gat), .Z(new_n451_));
  XNOR2_X1  g250(.A(new_n450_), .B(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n446_), .A2(new_n447_), .A3(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT101), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n452_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  AOI211_X1 g255(.A(KEYINPUT101), .B(new_n452_), .C1(new_n446_), .C2(new_n447_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n269_), .A2(new_n341_), .A3(new_n429_), .A4(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n408_), .A2(KEYINPUT32), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n419_), .A2(new_n462_), .A3(new_n421_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT98), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n464_), .B1(new_n424_), .B2(new_n461_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n406_), .A2(new_n407_), .A3(new_n461_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n466_), .A2(KEYINPUT98), .ZN(new_n467_));
  OAI211_X1 g266(.A(new_n458_), .B(new_n463_), .C1(new_n465_), .C2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT102), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n399_), .A2(new_n409_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT33), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n453_), .A2(new_n472_), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n446_), .A2(KEYINPUT33), .A3(new_n447_), .A4(new_n452_), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n442_), .A2(new_n443_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n452_), .B1(new_n475_), .B2(new_n431_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n430_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n477_));
  AND3_X1   g276(.A1(new_n476_), .A2(new_n477_), .A3(KEYINPUT96), .ZN(new_n478_));
  AOI21_X1  g277(.A(KEYINPUT96), .B1(new_n476_), .B2(new_n477_), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n473_), .B(new_n474_), .C1(new_n478_), .C2(new_n479_), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT97), .B1(new_n471_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n480_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT97), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n482_), .A2(new_n483_), .A3(new_n409_), .A4(new_n399_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n481_), .A2(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n424_), .A2(new_n464_), .A3(new_n461_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n466_), .A2(KEYINPUT98), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n488_), .A2(KEYINPUT102), .A3(new_n458_), .A4(new_n463_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n470_), .A2(new_n485_), .A3(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n458_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n491_));
  AOI22_X1  g290(.A1(new_n490_), .A2(new_n269_), .B1(new_n491_), .B2(new_n429_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n460_), .B1(new_n492_), .B2(new_n341_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT13), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G230gat), .A2(G233gat), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT65), .ZN(new_n496_));
  INV_X1    g295(.A(G99gat), .ZN(new_n497_));
  INV_X1    g296(.A(G106gat), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n496_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n499_), .A2(KEYINPUT64), .A3(KEYINPUT7), .ZN(new_n500_));
  AND3_X1   g299(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n501_));
  AOI21_X1  g300(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT64), .ZN(new_n504_));
  NOR2_X1   g303(.A1(G99gat), .A2(G106gat), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n504_), .B1(new_n505_), .B2(new_n496_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT7), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n507_), .B1(new_n505_), .B2(new_n504_), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n500_), .B(new_n503_), .C1(new_n506_), .C2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT8), .ZN(new_n510_));
  XOR2_X1   g309(.A(G85gat), .B(G92gat), .Z(new_n511_));
  NAND3_X1  g310(.A1(new_n509_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n510_), .B1(new_n509_), .B2(new_n511_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(KEYINPUT10), .B(G99gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G85gat), .A2(G92gat), .ZN(new_n516_));
  OAI22_X1  g315(.A1(new_n515_), .A2(G106gat), .B1(KEYINPUT9), .B2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n511_), .A2(KEYINPUT9), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(new_n503_), .ZN(new_n519_));
  OAI22_X1  g318(.A1(new_n513_), .A2(new_n514_), .B1(new_n517_), .B2(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G71gat), .B(G78gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G57gat), .B(G64gat), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n521_), .B1(KEYINPUT11), .B2(new_n522_), .ZN(new_n523_));
  XOR2_X1   g322(.A(G57gat), .B(G64gat), .Z(new_n524_));
  INV_X1    g323(.A(KEYINPUT11), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n523_), .A2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n522_), .A2(new_n521_), .A3(KEYINPUT11), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n520_), .A2(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n519_), .A2(new_n517_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n509_), .A2(new_n511_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT8), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n532_), .B1(new_n534_), .B2(new_n512_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(new_n529_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n495_), .B1(new_n531_), .B2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT66), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(KEYINPUT12), .B1(new_n535_), .B2(KEYINPUT67), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(new_n531_), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n520_), .A2(KEYINPUT67), .A3(KEYINPUT12), .A4(new_n530_), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n541_), .A2(new_n495_), .A3(new_n542_), .A4(new_n536_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G120gat), .B(G148gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(new_n206_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(KEYINPUT5), .B(G176gat), .ZN(new_n547_));
  XOR2_X1   g346(.A(new_n546_), .B(new_n547_), .Z(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NOR3_X1   g348(.A1(new_n539_), .A2(new_n544_), .A3(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n537_), .B(KEYINPUT66), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n548_), .B1(new_n551_), .B2(new_n543_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n494_), .B1(new_n550_), .B2(new_n552_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n549_), .B1(new_n539_), .B2(new_n544_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n551_), .A2(new_n543_), .A3(new_n548_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n554_), .A2(KEYINPUT13), .A3(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n553_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT15), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G29gat), .B(G36gat), .ZN(new_n559_));
  INV_X1    g358(.A(G50gat), .ZN(new_n560_));
  OR2_X1    g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n559_), .A2(new_n560_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(KEYINPUT68), .B(G43gat), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n561_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n563_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n558_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n561_), .A2(new_n562_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n563_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n570_), .A2(KEYINPUT15), .A3(new_n564_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n567_), .A2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(KEYINPUT69), .B(G15gat), .ZN(new_n573_));
  INV_X1    g372(.A(G22gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  XOR2_X1   g374(.A(KEYINPUT70), .B(G1gat), .Z(new_n576_));
  INV_X1    g375(.A(G8gat), .ZN(new_n577_));
  OAI21_X1  g376(.A(KEYINPUT14), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G1gat), .B(G8gat), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n575_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n579_), .B1(new_n575_), .B2(new_n578_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n572_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n570_), .A2(new_n564_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n582_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n585_), .B1(new_n580_), .B2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G229gat), .A2(G233gat), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n584_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n589_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n586_), .A2(new_n580_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n585_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n591_), .B1(new_n594_), .B2(new_n587_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n590_), .A2(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G113gat), .B(G141gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G169gat), .B(G197gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n596_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT73), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n596_), .A2(KEYINPUT73), .A3(new_n599_), .ZN(new_n603_));
  OAI21_X1  g402(.A(KEYINPUT74), .B1(new_n596_), .B2(new_n599_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT74), .ZN(new_n605_));
  INV_X1    g404(.A(new_n599_), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n590_), .A2(new_n595_), .A3(new_n605_), .A4(new_n606_), .ZN(new_n607_));
  AOI22_X1  g406(.A1(new_n602_), .A2(new_n603_), .B1(new_n604_), .B2(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n557_), .A2(new_n608_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n493_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n572_), .A2(new_n520_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n535_), .A2(new_n593_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(G232gat), .A2(G233gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT34), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT35), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n611_), .A2(new_n612_), .A3(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n615_), .A2(new_n616_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  AOI22_X1  g419(.A1(new_n572_), .A2(new_n520_), .B1(new_n616_), .B2(new_n615_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n619_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n621_), .A2(new_n622_), .A3(new_n612_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n620_), .A2(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G190gat), .B(G218gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(G134gat), .B(G162gat), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n625_), .B(new_n626_), .Z(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT36), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n624_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT37), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT36), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n620_), .A2(new_n631_), .A3(new_n627_), .A4(new_n623_), .ZN(new_n632_));
  AND3_X1   g431(.A1(new_n629_), .A2(new_n630_), .A3(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n630_), .B1(new_n629_), .B2(new_n632_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n527_), .A2(KEYINPUT71), .A3(new_n528_), .ZN(new_n636_));
  AOI21_X1  g435(.A(KEYINPUT71), .B1(new_n527_), .B2(new_n528_), .ZN(new_n637_));
  OAI211_X1 g436(.A(G231gat), .B(G233gat), .C1(new_n636_), .C2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT71), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n529_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(G231gat), .A2(G233gat), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n527_), .A2(KEYINPUT71), .A3(new_n528_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n640_), .A2(new_n641_), .A3(new_n642_), .ZN(new_n643_));
  AND3_X1   g442(.A1(new_n638_), .A2(new_n583_), .A3(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n583_), .B1(new_n638_), .B2(new_n643_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(G127gat), .B(G155gat), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(G211gat), .ZN(new_n647_));
  XNOR2_X1  g446(.A(KEYINPUT16), .B(G183gat), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n647_), .B(new_n648_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n649_), .A2(KEYINPUT17), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n649_), .A2(KEYINPUT17), .ZN(new_n651_));
  NOR4_X1   g450(.A1(new_n644_), .A2(new_n645_), .A3(new_n650_), .A4(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT67), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n653_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n643_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n641_), .B1(new_n640_), .B2(new_n642_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n592_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n638_), .A2(new_n583_), .A3(new_n643_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n657_), .A2(KEYINPUT67), .A3(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n654_), .A2(new_n659_), .A3(new_n650_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(KEYINPUT72), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT72), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n654_), .A2(new_n659_), .A3(new_n662_), .A4(new_n650_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n652_), .B1(new_n661_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n635_), .A2(new_n665_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n610_), .A2(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n458_), .B(KEYINPUT104), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n667_), .A2(new_n576_), .A3(new_n669_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT105), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT38), .ZN(new_n672_));
  OR2_X1    g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n671_), .A2(new_n672_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n629_), .A2(new_n632_), .ZN(new_n675_));
  XOR2_X1   g474(.A(new_n675_), .B(KEYINPUT106), .Z(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n677_), .A2(new_n665_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n610_), .A2(new_n678_), .ZN(new_n679_));
  OAI21_X1  g478(.A(G1gat), .B1(new_n679_), .B2(new_n459_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n673_), .A2(new_n674_), .A3(new_n680_), .ZN(G1324gat));
  INV_X1    g480(.A(new_n429_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n667_), .A2(new_n577_), .A3(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT39), .ZN(new_n684_));
  INV_X1    g483(.A(new_n679_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(new_n682_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n684_), .B1(new_n686_), .B2(G8gat), .ZN(new_n687_));
  AOI211_X1 g486(.A(KEYINPUT39), .B(new_n577_), .C1(new_n685_), .C2(new_n682_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n683_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT40), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n689_), .B(new_n690_), .ZN(G1325gat));
  INV_X1    g490(.A(new_n667_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n341_), .ZN(new_n693_));
  OR3_X1    g492(.A1(new_n692_), .A2(G15gat), .A3(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(G15gat), .B1(new_n679_), .B2(new_n693_), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n695_), .A2(KEYINPUT41), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(KEYINPUT41), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n694_), .A2(new_n696_), .A3(new_n697_), .ZN(G1326gat));
  OAI21_X1  g497(.A(G22gat), .B1(new_n679_), .B2(new_n269_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT42), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n268_), .A2(new_n574_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT107), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n700_), .B1(new_n692_), .B2(new_n702_), .ZN(G1327gat));
  NOR2_X1   g502(.A1(new_n664_), .A2(new_n675_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT111), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n610_), .A2(new_n705_), .ZN(new_n706_));
  OR3_X1    g505(.A1(new_n706_), .A2(G29gat), .A3(new_n459_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n609_), .A2(new_n665_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT43), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n635_), .A2(KEYINPUT108), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n635_), .A2(KEYINPUT108), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n710_), .B1(new_n493_), .B2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n635_), .A2(new_n710_), .ZN(new_n715_));
  AOI22_X1  g514(.A1(new_n469_), .A2(new_n468_), .B1(new_n481_), .B2(new_n484_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n268_), .B1(new_n716_), .B2(new_n489_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n491_), .A2(new_n429_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n693_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n715_), .B1(new_n719_), .B2(new_n460_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n709_), .B1(new_n714_), .B2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(KEYINPUT109), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT44), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n721_), .A2(KEYINPUT109), .A3(KEYINPUT44), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n668_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n726_), .A2(KEYINPUT110), .ZN(new_n727_));
  OAI21_X1  g526(.A(G29gat), .B1(new_n726_), .B2(KEYINPUT110), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n707_), .B1(new_n727_), .B2(new_n728_), .ZN(G1328gat));
  INV_X1    g528(.A(KEYINPUT46), .ZN(new_n730_));
  INV_X1    g529(.A(G36gat), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n724_), .A2(new_n725_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n731_), .B1(new_n732_), .B2(new_n682_), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n610_), .A2(new_n731_), .A3(new_n682_), .A4(new_n705_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT45), .Z(new_n735_));
  OAI21_X1  g534(.A(new_n730_), .B1(new_n733_), .B2(new_n735_), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n721_), .A2(KEYINPUT109), .A3(KEYINPUT44), .ZN(new_n737_));
  AOI21_X1  g536(.A(KEYINPUT44), .B1(new_n721_), .B2(KEYINPUT109), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  OAI21_X1  g538(.A(G36gat), .B1(new_n739_), .B2(new_n429_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n735_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n740_), .A2(KEYINPUT46), .A3(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n736_), .A2(new_n742_), .ZN(G1329gat));
  INV_X1    g542(.A(KEYINPUT47), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n341_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(G43gat), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n706_), .A2(G43gat), .A3(new_n693_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n744_), .B1(new_n746_), .B2(new_n748_), .ZN(new_n749_));
  AOI211_X1 g548(.A(KEYINPUT47), .B(new_n747_), .C1(new_n745_), .C2(G43gat), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1330gat));
  OAI21_X1  g550(.A(G50gat), .B1(new_n739_), .B2(new_n269_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n268_), .A2(new_n560_), .ZN(new_n753_));
  XOR2_X1   g552(.A(new_n753_), .B(KEYINPUT112), .Z(new_n754_));
  OAI21_X1  g553(.A(new_n752_), .B1(new_n706_), .B2(new_n754_), .ZN(G1331gat));
  INV_X1    g554(.A(new_n557_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n608_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n493_), .A2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(new_n666_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(G57gat), .B1(new_n761_), .B2(new_n669_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n759_), .A2(new_n678_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n458_), .A2(G57gat), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n762_), .B1(new_n763_), .B2(new_n764_), .ZN(G1332gat));
  INV_X1    g564(.A(G64gat), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n766_), .B1(new_n763_), .B2(new_n682_), .ZN(new_n767_));
  XOR2_X1   g566(.A(new_n767_), .B(KEYINPUT48), .Z(new_n768_));
  NAND3_X1  g567(.A1(new_n761_), .A2(new_n766_), .A3(new_n682_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(G1333gat));
  NAND2_X1  g569(.A1(new_n763_), .A2(new_n341_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(G71gat), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT49), .ZN(new_n773_));
  OR2_X1    g572(.A1(new_n693_), .A2(G71gat), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n773_), .B1(new_n760_), .B2(new_n774_), .ZN(G1334gat));
  INV_X1    g574(.A(G78gat), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n776_), .B1(new_n763_), .B2(new_n268_), .ZN(new_n777_));
  XOR2_X1   g576(.A(new_n777_), .B(KEYINPUT50), .Z(new_n778_));
  NAND3_X1  g577(.A1(new_n761_), .A2(new_n776_), .A3(new_n268_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(G1335gat));
  INV_X1    g579(.A(G85gat), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n759_), .A2(new_n705_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n781_), .B1(new_n782_), .B2(new_n668_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT113), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n714_), .A2(new_n720_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n758_), .A2(new_n665_), .ZN(new_n786_));
  XOR2_X1   g585(.A(new_n786_), .B(KEYINPUT114), .Z(new_n787_));
  NOR2_X1   g586(.A1(new_n785_), .A2(new_n787_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n459_), .A2(new_n781_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n784_), .B1(new_n788_), .B2(new_n789_), .ZN(G1336gat));
  INV_X1    g589(.A(new_n782_), .ZN(new_n791_));
  AOI21_X1  g590(.A(G92gat), .B1(new_n791_), .B2(new_n682_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n429_), .A2(new_n343_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n792_), .B1(new_n788_), .B2(new_n793_), .ZN(G1337gat));
  NOR3_X1   g593(.A1(new_n782_), .A2(new_n515_), .A3(new_n693_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n788_), .A2(new_n341_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n795_), .B1(new_n796_), .B2(G99gat), .ZN(new_n797_));
  XOR2_X1   g596(.A(new_n797_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g597(.A1(new_n791_), .A2(new_n498_), .A3(new_n268_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT52), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n788_), .A2(new_n268_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n800_), .B1(new_n801_), .B2(G106gat), .ZN(new_n802_));
  AOI211_X1 g601(.A(KEYINPUT52), .B(new_n498_), .C1(new_n788_), .C2(new_n268_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n799_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(KEYINPUT53), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n806_), .B(new_n799_), .C1(new_n802_), .C2(new_n803_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n805_), .A2(new_n807_), .ZN(G1339gat));
  OAI211_X1 g607(.A(new_n664_), .B(new_n608_), .C1(new_n633_), .C2(new_n634_), .ZN(new_n809_));
  OR4_X1    g608(.A1(KEYINPUT115), .A2(new_n557_), .A3(new_n809_), .A4(KEYINPUT54), .ZN(new_n810_));
  INV_X1    g609(.A(new_n809_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n756_), .A2(new_n811_), .A3(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT115), .ZN(new_n814_));
  OAI21_X1  g613(.A(KEYINPUT54), .B1(new_n557_), .B2(new_n809_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT116), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  OAI211_X1 g616(.A(KEYINPUT116), .B(KEYINPUT54), .C1(new_n557_), .C2(new_n809_), .ZN(new_n818_));
  AND4_X1   g617(.A1(new_n810_), .A2(new_n814_), .A3(new_n817_), .A4(new_n818_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n541_), .A2(KEYINPUT55), .A3(new_n542_), .A4(new_n536_), .ZN(new_n820_));
  OAI21_X1  g619(.A(KEYINPUT55), .B1(new_n495_), .B2(KEYINPUT117), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n543_), .A2(new_n820_), .A3(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n821_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n541_), .A2(new_n542_), .A3(new_n536_), .A4(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n822_), .A2(KEYINPUT118), .A3(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n549_), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT118), .B1(new_n822_), .B2(new_n824_), .ZN(new_n827_));
  OAI21_X1  g626(.A(KEYINPUT56), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n822_), .A2(new_n824_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT118), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT56), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n831_), .A2(new_n832_), .A3(new_n549_), .A4(new_n825_), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n828_), .A2(new_n833_), .A3(new_n555_), .A4(new_n757_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n584_), .A2(new_n588_), .A3(new_n591_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n589_), .B1(new_n594_), .B2(new_n587_), .ZN(new_n836_));
  AND3_X1   g635(.A1(new_n835_), .A2(new_n836_), .A3(new_n599_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n837_), .B1(new_n604_), .B2(new_n607_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n838_), .B1(new_n550_), .B2(new_n552_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n834_), .A2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n675_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT57), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n635_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n828_), .A2(new_n833_), .A3(new_n555_), .A4(new_n838_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT58), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n844_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n847_), .B1(new_n846_), .B2(new_n845_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n840_), .A2(KEYINPUT57), .A3(new_n675_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n843_), .A2(new_n848_), .A3(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n819_), .B1(new_n850_), .B2(new_n665_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n269_), .A2(new_n429_), .A3(new_n341_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n852_), .A2(new_n668_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n851_), .A2(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(G113gat), .B1(new_n855_), .B2(new_n757_), .ZN(new_n856_));
  OAI21_X1  g655(.A(KEYINPUT59), .B1(new_n851_), .B2(new_n854_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT59), .ZN(new_n858_));
  AOI21_X1  g657(.A(KEYINPUT57), .B1(new_n840_), .B2(new_n675_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n675_), .ZN(new_n860_));
  AOI211_X1 g659(.A(new_n842_), .B(new_n860_), .C1(new_n834_), .C2(new_n839_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n859_), .A2(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n664_), .B1(new_n862_), .B2(new_n848_), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n858_), .B(new_n853_), .C1(new_n863_), .C2(new_n819_), .ZN(new_n864_));
  AND3_X1   g663(.A1(new_n857_), .A2(KEYINPUT119), .A3(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(KEYINPUT119), .B1(new_n857_), .B2(new_n864_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  AND2_X1   g666(.A1(new_n757_), .A2(G113gat), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n856_), .B1(new_n867_), .B2(new_n868_), .ZN(G1340gat));
  NAND2_X1  g668(.A1(new_n857_), .A2(new_n864_), .ZN(new_n870_));
  OAI21_X1  g669(.A(G120gat), .B1(new_n870_), .B2(new_n756_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n756_), .A2(KEYINPUT60), .ZN(new_n872_));
  MUX2_X1   g671(.A(new_n872_), .B(KEYINPUT60), .S(G120gat), .Z(new_n873_));
  NAND2_X1  g672(.A1(new_n855_), .A2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n871_), .A2(new_n874_), .ZN(G1341gat));
  NOR2_X1   g674(.A1(new_n665_), .A2(new_n280_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n865_), .A2(new_n866_), .A3(new_n877_), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n851_), .A2(new_n665_), .A3(new_n854_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n880_), .A2(KEYINPUT120), .A3(new_n280_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT120), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n882_), .B1(new_n879_), .B2(G127gat), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n881_), .A2(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(KEYINPUT121), .B1(new_n878_), .B2(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT119), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n870_), .A2(new_n886_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n857_), .A2(KEYINPUT119), .A3(new_n864_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n887_), .A2(new_n888_), .A3(new_n876_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT121), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n889_), .A2(new_n890_), .A3(new_n883_), .A4(new_n881_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n885_), .A2(new_n891_), .ZN(G1342gat));
  AOI21_X1  g691(.A(G134gat), .B1(new_n855_), .B2(new_n677_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n844_), .A2(new_n281_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n893_), .B1(new_n867_), .B2(new_n894_), .ZN(G1343gat));
  NAND2_X1  g694(.A1(new_n850_), .A2(new_n665_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n819_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  NOR4_X1   g697(.A1(new_n682_), .A2(new_n269_), .A3(new_n341_), .A4(new_n668_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n900_), .A2(new_n608_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(new_n226_), .ZN(G1344gat));
  NOR2_X1   g701(.A1(new_n900_), .A2(new_n756_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(new_n227_), .ZN(G1345gat));
  OR3_X1    g703(.A1(new_n900_), .A2(KEYINPUT122), .A3(new_n665_), .ZN(new_n905_));
  OAI21_X1  g704(.A(KEYINPUT122), .B1(new_n900_), .B2(new_n665_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(KEYINPUT61), .B(G155gat), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n907_), .B(new_n908_), .ZN(G1346gat));
  INV_X1    g708(.A(new_n900_), .ZN(new_n910_));
  AOI21_X1  g709(.A(G162gat), .B1(new_n910_), .B2(new_n677_), .ZN(new_n911_));
  AND2_X1   g710(.A1(new_n713_), .A2(G162gat), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n911_), .B1(new_n910_), .B2(new_n912_), .ZN(G1347gat));
  NAND3_X1  g712(.A1(new_n682_), .A2(new_n668_), .A3(new_n341_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(KEYINPUT123), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(new_n757_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(KEYINPUT124), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n851_), .A2(new_n268_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(G169gat), .ZN(new_n920_));
  AND2_X1   g719(.A1(new_n920_), .A2(KEYINPUT62), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n920_), .A2(KEYINPUT62), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n918_), .A2(new_n915_), .ZN(new_n923_));
  OR2_X1    g722(.A1(new_n608_), .A2(new_n325_), .ZN(new_n924_));
  OAI22_X1  g723(.A1(new_n921_), .A2(new_n922_), .B1(new_n923_), .B2(new_n924_), .ZN(G1348gat));
  NOR2_X1   g724(.A1(new_n923_), .A2(new_n756_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n926_), .A2(new_n324_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n927_), .B1(G176gat), .B2(new_n926_), .ZN(G1349gat));
  NAND3_X1  g727(.A1(new_n918_), .A2(new_n664_), .A3(new_n915_), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT125), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n929_), .B1(new_n930_), .B2(G183gat), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n319_), .B1(KEYINPUT125), .B2(G183gat), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n931_), .B1(new_n929_), .B2(new_n932_), .ZN(G1350gat));
  NOR2_X1   g732(.A1(new_n353_), .A2(new_n354_), .ZN(new_n934_));
  OR3_X1    g733(.A1(new_n923_), .A2(new_n934_), .A3(new_n676_), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n918_), .A2(new_n635_), .A3(new_n915_), .ZN(new_n936_));
  AND3_X1   g735(.A1(new_n936_), .A2(KEYINPUT126), .A3(G190gat), .ZN(new_n937_));
  AOI21_X1  g736(.A(KEYINPUT126), .B1(new_n936_), .B2(G190gat), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n935_), .B1(new_n937_), .B2(new_n938_), .ZN(G1351gat));
  AND4_X1   g738(.A1(new_n491_), .A2(new_n898_), .A3(new_n682_), .A4(new_n693_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n940_), .A2(new_n757_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g741(.A1(new_n940_), .A2(new_n557_), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n943_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g743(.A(new_n665_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n945_));
  XNOR2_X1  g744(.A(new_n945_), .B(KEYINPUT127), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n940_), .A2(new_n946_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n948_));
  XOR2_X1   g747(.A(new_n947_), .B(new_n948_), .Z(G1354gat));
  AOI21_X1  g748(.A(G218gat), .B1(new_n940_), .B2(new_n677_), .ZN(new_n950_));
  AND2_X1   g749(.A1(new_n635_), .A2(G218gat), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n950_), .B1(new_n940_), .B2(new_n951_), .ZN(G1355gat));
endmodule


