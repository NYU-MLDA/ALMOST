//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 0 0 0 1 0 1 0 0 1 0 0 1 0 0 0 0 1 1 1 1 0 0 1 1 0 0 1 0 0 1 1 0 0 0 0 1 1 1 1 1 0 1 1 0 0 1 1 1 1 0 1 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n761_, new_n762_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n798_, new_n799_, new_n800_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n907_, new_n909_, new_n910_, new_n912_, new_n913_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n926_, new_n927_, new_n928_,
    new_n930_, new_n931_, new_n933_, new_n934_, new_n936_, new_n937_,
    new_n938_, new_n940_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n956_, new_n957_;
  XOR2_X1   g000(.A(G134gat), .B(G162gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G190gat), .B(G218gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT36), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n204_), .A2(new_n205_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G232gat), .A2(G233gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT34), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT35), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT8), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT68), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT7), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NOR2_X1   g013(.A1(KEYINPUT68), .A2(KEYINPUT7), .ZN(new_n215_));
  OAI22_X1  g014(.A1(new_n214_), .A2(new_n215_), .B1(G99gat), .B2(G106gat), .ZN(new_n216_));
  INV_X1    g015(.A(G99gat), .ZN(new_n217_));
  INV_X1    g016(.A(G106gat), .ZN(new_n218_));
  OAI211_X1 g017(.A(new_n217_), .B(new_n218_), .C1(new_n212_), .C2(new_n213_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n216_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G99gat), .A2(G106gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n221_), .B(KEYINPUT6), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n220_), .B1(KEYINPUT70), .B2(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n223_), .B1(KEYINPUT70), .B2(new_n222_), .ZN(new_n224_));
  XOR2_X1   g023(.A(G85gat), .B(G92gat), .Z(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(KEYINPUT69), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n211_), .B1(new_n224_), .B2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n216_), .A2(new_n222_), .A3(new_n219_), .ZN(new_n228_));
  AND3_X1   g027(.A1(new_n226_), .A2(new_n211_), .A3(new_n228_), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n227_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT66), .ZN(new_n231_));
  OAI211_X1 g030(.A(G85gat), .B(G92gat), .C1(new_n231_), .C2(KEYINPUT9), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n231_), .B(KEYINPUT9), .C1(G85gat), .C2(G92gat), .ZN(new_n233_));
  AND2_X1   g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n232_), .A2(new_n233_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT10), .B(G99gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT65), .ZN(new_n237_));
  OAI221_X1 g036(.A(new_n222_), .B1(new_n234_), .B2(new_n235_), .C1(new_n237_), .C2(G106gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT67), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n230_), .A2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G29gat), .B(G36gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G43gat), .B(G50gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT15), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n240_), .A2(KEYINPUT73), .A3(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT73), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n227_), .A2(new_n229_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT67), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n238_), .B(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n244_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n246_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n245_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT74), .ZN(new_n255_));
  INV_X1    g054(.A(new_n243_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n255_), .B1(new_n240_), .B2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n250_), .A2(KEYINPUT74), .A3(new_n243_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n210_), .B1(new_n254_), .B2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n240_), .A2(new_n244_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n210_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n209_), .A2(KEYINPUT35), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n259_), .A2(new_n261_), .A3(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n206_), .B(new_n207_), .C1(new_n260_), .C2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n259_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n262_), .B1(new_n268_), .B2(new_n253_), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n269_), .A2(new_n205_), .A3(new_n204_), .A4(new_n265_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n267_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT37), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n267_), .A2(KEYINPUT37), .A3(new_n270_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G57gat), .B(G64gat), .ZN(new_n277_));
  OR2_X1    g076(.A1(new_n277_), .A2(KEYINPUT11), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(KEYINPUT11), .ZN(new_n279_));
  XOR2_X1   g078(.A(G71gat), .B(G78gat), .Z(new_n280_));
  NAND3_X1  g079(.A1(new_n278_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n281_));
  OR2_X1    g080(.A1(new_n279_), .A2(new_n280_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G15gat), .B(G22gat), .ZN(new_n284_));
  INV_X1    g083(.A(G1gat), .ZN(new_n285_));
  INV_X1    g084(.A(G8gat), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT14), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n284_), .A2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G1gat), .B(G8gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n283_), .B(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G231gat), .A2(G233gat), .ZN(new_n292_));
  XOR2_X1   g091(.A(new_n291_), .B(new_n292_), .Z(new_n293_));
  XOR2_X1   g092(.A(G127gat), .B(G155gat), .Z(new_n294_));
  XNOR2_X1  g093(.A(G183gat), .B(G211gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  XOR2_X1   g095(.A(KEYINPUT75), .B(KEYINPUT16), .Z(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT17), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n293_), .A2(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n293_), .A2(KEYINPUT17), .A3(new_n298_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n276_), .A2(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G226gat), .A2(G233gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT21), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT90), .ZN(new_n310_));
  INV_X1    g109(.A(G204gat), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n310_), .B1(new_n311_), .B2(G197gat), .ZN(new_n312_));
  INV_X1    g111(.A(G197gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n313_), .A2(KEYINPUT90), .A3(G204gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT89), .ZN(new_n316_));
  AND2_X1   g115(.A1(KEYINPUT88), .A2(G204gat), .ZN(new_n317_));
  NOR2_X1   g116(.A1(KEYINPUT88), .A2(G204gat), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n316_), .B1(new_n319_), .B2(G197gat), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT88), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(new_n311_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(KEYINPUT88), .A2(G204gat), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n322_), .A2(new_n316_), .A3(G197gat), .A4(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n309_), .B(new_n315_), .C1(new_n320_), .C2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G211gat), .B(G218gat), .ZN(new_n327_));
  NOR3_X1   g126(.A1(new_n317_), .A2(new_n318_), .A3(G197gat), .ZN(new_n328_));
  OAI21_X1  g127(.A(KEYINPUT21), .B1(new_n313_), .B2(new_n311_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n327_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n326_), .A2(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n327_), .A2(new_n309_), .ZN(new_n333_));
  AND2_X1   g132(.A1(new_n312_), .A2(new_n314_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n322_), .A2(G197gat), .A3(new_n323_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(KEYINPUT89), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n334_), .B1(new_n336_), .B2(new_n324_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT91), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n333_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  AOI211_X1 g138(.A(KEYINPUT91), .B(new_n334_), .C1(new_n336_), .C2(new_n324_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n332_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT22), .B(G169gat), .ZN(new_n342_));
  INV_X1    g141(.A(G176gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT78), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G169gat), .A2(G176gat), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G183gat), .A2(G190gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT23), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT23), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n351_), .A2(G183gat), .A3(G190gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(G183gat), .A2(G190gat), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n348_), .B1(new_n353_), .B2(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n342_), .A2(KEYINPUT78), .A3(new_n343_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n346_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  AND3_X1   g157(.A1(new_n349_), .A2(KEYINPUT77), .A3(KEYINPUT23), .ZN(new_n359_));
  AOI21_X1  g158(.A(KEYINPUT77), .B1(new_n349_), .B2(KEYINPUT23), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n352_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT76), .ZN(new_n362_));
  INV_X1    g161(.A(G169gat), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n362_), .A2(new_n363_), .A3(new_n343_), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT76), .B1(G169gat), .B2(G176gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT24), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n364_), .A2(KEYINPUT24), .A3(new_n365_), .A4(new_n347_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(KEYINPUT26), .B(G190gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(KEYINPUT25), .B(G183gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n361_), .A2(new_n368_), .A3(new_n369_), .A4(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n358_), .A2(new_n373_), .ZN(new_n374_));
  OAI211_X1 g173(.A(KEYINPUT95), .B(KEYINPUT20), .C1(new_n341_), .C2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n361_), .A2(new_n355_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n348_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(G169gat), .A2(G176gat), .ZN(new_n378_));
  AOI22_X1  g177(.A1(new_n350_), .A2(new_n352_), .B1(new_n367_), .B2(new_n378_), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n379_), .A2(new_n369_), .ZN(new_n380_));
  INV_X1    g179(.A(G183gat), .ZN(new_n381_));
  AND2_X1   g180(.A1(new_n381_), .A2(KEYINPUT25), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n381_), .A2(KEYINPUT25), .ZN(new_n383_));
  OAI21_X1  g182(.A(KEYINPUT96), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT96), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n371_), .A2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n384_), .A2(new_n386_), .A3(new_n370_), .ZN(new_n387_));
  AOI22_X1  g186(.A1(new_n376_), .A2(new_n377_), .B1(new_n380_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n341_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n375_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n374_), .ZN(new_n392_));
  OAI211_X1 g191(.A(new_n392_), .B(new_n332_), .C1(new_n340_), .C2(new_n339_), .ZN(new_n393_));
  AOI21_X1  g192(.A(KEYINPUT95), .B1(new_n393_), .B2(KEYINPUT20), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n308_), .B1(new_n391_), .B2(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n330_), .B1(new_n337_), .B2(new_n309_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n333_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n315_), .B1(new_n320_), .B2(new_n325_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n397_), .B1(new_n398_), .B2(KEYINPUT91), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n337_), .A2(new_n338_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n396_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n401_), .A2(new_n392_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n388_), .B(new_n332_), .C1(new_n339_), .C2(new_n340_), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n403_), .A2(KEYINPUT20), .A3(new_n307_), .A4(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n395_), .A2(new_n405_), .ZN(new_n406_));
  XOR2_X1   g205(.A(G8gat), .B(G36gat), .Z(new_n407_));
  XNOR2_X1  g206(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G64gat), .B(G92gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n406_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n411_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n395_), .A2(new_n405_), .A3(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT27), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NOR4_X1   g216(.A1(new_n391_), .A2(new_n394_), .A3(KEYINPUT102), .A4(new_n308_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT102), .ZN(new_n419_));
  AND3_X1   g218(.A1(new_n404_), .A2(KEYINPUT101), .A3(KEYINPUT20), .ZN(new_n420_));
  AOI21_X1  g219(.A(KEYINPUT101), .B1(new_n404_), .B2(KEYINPUT20), .ZN(new_n421_));
  NOR3_X1   g220(.A1(new_n420_), .A2(new_n421_), .A3(new_n402_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n419_), .B1(new_n422_), .B2(new_n307_), .ZN(new_n423_));
  NOR3_X1   g222(.A1(new_n391_), .A2(new_n308_), .A3(new_n394_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n418_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n426_), .A2(new_n413_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n414_), .A2(KEYINPUT27), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n417_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G225gat), .A2(G233gat), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT4), .ZN(new_n432_));
  NOR2_X1   g231(.A1(G141gat), .A2(G148gat), .ZN(new_n433_));
  NOR2_X1   g232(.A1(KEYINPUT84), .A2(KEYINPUT3), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  OAI22_X1  g234(.A1(KEYINPUT84), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G141gat), .A2(G148gat), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT2), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n435_), .A2(new_n436_), .A3(new_n439_), .A4(new_n440_), .ZN(new_n441_));
  XOR2_X1   g240(.A(G155gat), .B(G162gat), .Z(new_n442_));
  INV_X1    g241(.A(G155gat), .ZN(new_n443_));
  INV_X1    g242(.A(G162gat), .ZN(new_n444_));
  OAI21_X1  g243(.A(KEYINPUT1), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT1), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n446_), .A2(G155gat), .A3(G162gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n443_), .A2(new_n444_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n445_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  XOR2_X1   g248(.A(G141gat), .B(G148gat), .Z(new_n450_));
  AOI22_X1  g249(.A1(new_n441_), .A2(new_n442_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(G134gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(G127gat), .ZN(new_n453_));
  INV_X1    g252(.A(G127gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(G134gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(G120gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(G113gat), .ZN(new_n458_));
  INV_X1    g257(.A(G113gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(G120gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n458_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n456_), .A2(new_n461_), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n453_), .A2(new_n455_), .A3(new_n458_), .A4(new_n460_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(KEYINPUT98), .B1(new_n451_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n441_), .A2(new_n442_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n449_), .A2(new_n450_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n464_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n465_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n468_), .A2(KEYINPUT98), .A3(new_n469_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n432_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(KEYINPUT99), .B(KEYINPUT4), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n470_), .A2(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n431_), .B1(new_n473_), .B2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n471_), .A2(new_n430_), .A3(new_n472_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G1gat), .B(G29gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(G85gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(KEYINPUT0), .B(G57gat), .ZN(new_n481_));
  XOR2_X1   g280(.A(new_n480_), .B(new_n481_), .Z(new_n482_));
  NAND2_X1  g281(.A1(new_n478_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n482_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n476_), .A2(new_n484_), .A3(new_n477_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(KEYINPUT93), .B(KEYINPUT29), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n468_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  OAI211_X1 g288(.A(G228gat), .B(G233gat), .C1(new_n401_), .C2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G78gat), .B(G106gat), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT92), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G228gat), .A2(G233gat), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT29), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n493_), .B1(new_n451_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n341_), .A2(new_n492_), .A3(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n492_), .B1(new_n341_), .B2(new_n496_), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n490_), .B(new_n491_), .C1(new_n498_), .C2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT87), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT92), .B1(new_n401_), .B2(new_n495_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(new_n497_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n491_), .B1(new_n503_), .B2(new_n490_), .ZN(new_n504_));
  XOR2_X1   g303(.A(KEYINPUT86), .B(KEYINPUT28), .Z(new_n505_));
  INV_X1    g304(.A(KEYINPUT85), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n451_), .A2(new_n506_), .A3(new_n494_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n506_), .B1(new_n451_), .B2(new_n494_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n505_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT85), .B1(new_n468_), .B2(KEYINPUT29), .ZN(new_n511_));
  INV_X1    g310(.A(new_n505_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n511_), .A2(new_n507_), .A3(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n510_), .A2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G22gat), .B(G50gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  NOR3_X1   g315(.A1(new_n501_), .A2(new_n504_), .A3(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n515_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n514_), .B(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT87), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n493_), .B1(new_n341_), .B2(new_n488_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n521_), .B1(new_n502_), .B2(new_n497_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n520_), .B1(new_n522_), .B2(new_n491_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n490_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n491_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n519_), .B1(new_n523_), .B2(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n517_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  AND3_X1   g328(.A1(new_n358_), .A2(new_n373_), .A3(KEYINPUT30), .ZN(new_n530_));
  AOI21_X1  g329(.A(KEYINPUT30), .B1(new_n358_), .B2(new_n373_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G71gat), .B(G99gat), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT80), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(G15gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n533_), .B(KEYINPUT80), .ZN(new_n537_));
  INV_X1    g336(.A(G15gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n536_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G227gat), .A2(G233gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n536_), .A2(new_n539_), .A3(G227gat), .A4(G233gat), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n532_), .A2(new_n544_), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n542_), .B(new_n543_), .C1(new_n530_), .C2(new_n531_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT79), .B(G43gat), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n545_), .A2(new_n546_), .A3(new_n548_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT81), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n464_), .B(KEYINPUT31), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT82), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n553_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  OR2_X1    g356(.A1(new_n552_), .A2(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(KEYINPUT82), .B1(new_n552_), .B2(KEYINPUT81), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n558_), .B1(new_n559_), .B2(new_n555_), .ZN(new_n560_));
  NOR4_X1   g359(.A1(new_n429_), .A2(new_n486_), .A3(new_n529_), .A4(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT83), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n558_), .B(new_n562_), .C1(new_n559_), .C2(new_n555_), .ZN(new_n563_));
  AND3_X1   g362(.A1(new_n545_), .A2(new_n548_), .A3(new_n546_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n548_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n565_));
  OAI21_X1  g364(.A(KEYINPUT81), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n555_), .B1(new_n566_), .B2(new_n556_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n552_), .A2(new_n557_), .ZN(new_n568_));
  OAI21_X1  g367(.A(KEYINPUT83), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n563_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT33), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n483_), .A2(KEYINPUT100), .A3(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n484_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n574_));
  OR3_X1    g373(.A1(new_n473_), .A2(new_n431_), .A3(new_n475_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n471_), .A2(new_n472_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n482_), .B1(new_n576_), .B2(new_n431_), .ZN(new_n577_));
  AOI22_X1  g376(.A1(new_n574_), .A2(KEYINPUT33), .B1(new_n575_), .B2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT100), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n579_), .B1(new_n574_), .B2(KEYINPUT33), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n573_), .A2(new_n578_), .A3(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n414_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n413_), .B1(new_n395_), .B2(new_n405_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n581_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n413_), .A2(KEYINPUT32), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n395_), .A2(new_n405_), .A3(new_n586_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n486_), .A2(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n588_), .B1(new_n426_), .B2(new_n586_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n529_), .B1(new_n585_), .B2(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n391_), .A2(new_n394_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n591_), .A2(new_n419_), .A3(new_n307_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n404_), .A2(KEYINPUT20), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT101), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n404_), .A2(KEYINPUT101), .A3(KEYINPUT20), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n595_), .A2(new_n403_), .A3(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(KEYINPUT102), .B1(new_n597_), .B2(new_n308_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n592_), .B1(new_n598_), .B2(new_n424_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n428_), .B1(new_n599_), .B2(new_n411_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n486_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n601_), .B1(new_n517_), .B2(new_n527_), .ZN(new_n602_));
  AOI21_X1  g401(.A(KEYINPUT27), .B1(new_n412_), .B2(new_n414_), .ZN(new_n603_));
  NOR3_X1   g402(.A1(new_n600_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n571_), .B1(new_n590_), .B2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT103), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n573_), .A2(new_n578_), .A3(new_n580_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n415_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n486_), .A2(new_n587_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n586_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n610_), .B1(new_n599_), .B2(new_n611_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n528_), .B1(new_n609_), .B2(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n516_), .B1(new_n501_), .B2(new_n504_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n523_), .A2(new_n526_), .A3(new_n519_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n486_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  OAI211_X1 g415(.A(new_n616_), .B(new_n417_), .C1(new_n427_), .C2(new_n428_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n613_), .A2(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n618_), .A2(KEYINPUT103), .A3(new_n571_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n561_), .B1(new_n607_), .B2(new_n619_), .ZN(new_n620_));
  OR2_X1    g419(.A1(new_n290_), .A2(new_n256_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(G229gat), .A2(G233gat), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n244_), .A2(new_n290_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n290_), .B(new_n256_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n622_), .ZN(new_n626_));
  AOI22_X1  g425(.A1(new_n623_), .A2(new_n624_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  XOR2_X1   g426(.A(G113gat), .B(G141gat), .Z(new_n628_));
  XNOR2_X1  g427(.A(G169gat), .B(G197gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n628_), .B(new_n629_), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n627_), .A2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n627_), .A2(new_n630_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT13), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n230_), .A2(new_n239_), .A3(new_n283_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n283_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n637_), .B1(new_n247_), .B2(new_n249_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n636_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(G230gat), .A2(G233gat), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT64), .Z(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n639_), .A2(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n636_), .A2(KEYINPUT12), .A3(new_n638_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT12), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n240_), .A2(new_n645_), .A3(new_n637_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n644_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(new_n642_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n643_), .A2(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(G120gat), .B(G148gat), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT5), .ZN(new_n651_));
  XOR2_X1   g450(.A(G176gat), .B(G204gat), .Z(new_n652_));
  XNOR2_X1  g451(.A(new_n651_), .B(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  OR2_X1    g453(.A1(new_n654_), .A2(KEYINPUT71), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n655_), .B(KEYINPUT72), .Z(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n649_), .A2(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n639_), .A2(new_n642_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n641_), .B1(new_n644_), .B2(new_n646_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n661_), .A2(new_n656_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n635_), .B1(new_n658_), .B2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n649_), .A2(new_n657_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n661_), .A2(new_n656_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n664_), .A2(new_n665_), .A3(KEYINPUT13), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n663_), .A2(new_n666_), .ZN(new_n667_));
  NOR4_X1   g466(.A1(new_n304_), .A2(new_n620_), .A3(new_n634_), .A4(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n486_), .B(KEYINPUT104), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n668_), .A2(new_n285_), .A3(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT38), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT105), .Z(new_n674_));
  INV_X1    g473(.A(new_n561_), .ZN(new_n675_));
  AOI21_X1  g474(.A(KEYINPUT103), .B1(new_n618_), .B2(new_n571_), .ZN(new_n676_));
  AOI211_X1 g475(.A(new_n606_), .B(new_n570_), .C1(new_n613_), .C2(new_n617_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n675_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(new_n271_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n667_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(new_n633_), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n679_), .A2(new_n302_), .A3(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n285_), .B1(new_n682_), .B2(new_n486_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n683_), .B1(new_n672_), .B2(new_n671_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n674_), .A2(new_n684_), .ZN(G1324gat));
  AOI21_X1  g484(.A(new_n286_), .B1(new_n682_), .B2(new_n429_), .ZN(new_n686_));
  XOR2_X1   g485(.A(new_n686_), .B(KEYINPUT39), .Z(new_n687_));
  NAND3_X1  g486(.A1(new_n668_), .A2(new_n286_), .A3(new_n429_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n689_), .B(KEYINPUT40), .Z(G1325gat));
  AOI21_X1  g489(.A(new_n538_), .B1(new_n682_), .B2(new_n570_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT41), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n668_), .A2(new_n538_), .A3(new_n570_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1326gat));
  INV_X1    g493(.A(G22gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n695_), .B1(new_n682_), .B2(new_n529_), .ZN(new_n696_));
  XOR2_X1   g495(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n697_));
  XNOR2_X1  g496(.A(new_n696_), .B(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n668_), .A2(new_n695_), .A3(new_n529_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1327gat));
  NOR2_X1   g499(.A1(new_n620_), .A2(new_n634_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n271_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(new_n302_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n703_), .A2(new_n667_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n701_), .A2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(G29gat), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n706_), .A2(new_n707_), .A3(new_n486_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT108), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n680_), .A2(new_n633_), .A3(new_n302_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n620_), .A2(new_n276_), .A3(KEYINPUT43), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT43), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n713_), .B1(new_n678_), .B2(new_n275_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n711_), .B1(new_n712_), .B2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT107), .ZN(new_n716_));
  AOI21_X1  g515(.A(KEYINPUT44), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(KEYINPUT43), .B1(new_n620_), .B2(new_n276_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n678_), .A2(new_n713_), .A3(new_n275_), .ZN(new_n719_));
  AOI211_X1 g518(.A(new_n716_), .B(new_n710_), .C1(new_n718_), .C2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n710_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n722_));
  AOI22_X1  g521(.A1(new_n717_), .A2(new_n721_), .B1(KEYINPUT44), .B2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(new_n670_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n709_), .B1(new_n724_), .B2(G29gat), .ZN(new_n725_));
  AOI211_X1 g524(.A(KEYINPUT108), .B(new_n707_), .C1(new_n723_), .C2(new_n670_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n708_), .B1(new_n725_), .B2(new_n726_), .ZN(G1328gat));
  INV_X1    g526(.A(G36gat), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n429_), .A2(new_n728_), .ZN(new_n729_));
  OR3_X1    g528(.A1(new_n705_), .A2(KEYINPUT110), .A3(new_n729_), .ZN(new_n730_));
  OAI21_X1  g529(.A(KEYINPUT110), .B1(new_n705_), .B2(new_n729_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  XOR2_X1   g531(.A(KEYINPUT111), .B(KEYINPUT45), .Z(new_n733_));
  XNOR2_X1  g532(.A(new_n732_), .B(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n722_), .A2(KEYINPUT44), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT44), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n736_), .B1(new_n722_), .B2(KEYINPUT107), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n429_), .B(new_n735_), .C1(new_n737_), .C2(new_n720_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT109), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n738_), .A2(new_n739_), .A3(G36gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n738_), .B2(G36gat), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n734_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT46), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  OAI211_X1 g543(.A(KEYINPUT46), .B(new_n734_), .C1(new_n740_), .C2(new_n741_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1329gat));
  INV_X1    g545(.A(G43gat), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n747_), .B1(new_n705_), .B2(new_n571_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT112), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n560_), .A2(new_n747_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n723_), .B2(new_n750_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n735_), .B1(new_n737_), .B2(new_n720_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n750_), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n752_), .A2(KEYINPUT112), .A3(new_n753_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n748_), .B1(new_n751_), .B2(new_n754_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(KEYINPUT113), .B(KEYINPUT47), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n748_), .B(new_n756_), .C1(new_n751_), .C2(new_n754_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(G1330gat));
  AOI21_X1  g559(.A(G50gat), .B1(new_n706_), .B2(new_n529_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n529_), .A2(G50gat), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n723_), .B2(new_n762_), .ZN(G1331gat));
  NOR2_X1   g562(.A1(new_n302_), .A2(new_n633_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  NOR3_X1   g564(.A1(new_n679_), .A2(new_n680_), .A3(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(G57gat), .B1(new_n767_), .B2(new_n601_), .ZN(new_n768_));
  NOR4_X1   g567(.A1(new_n304_), .A2(new_n620_), .A3(new_n633_), .A4(new_n680_), .ZN(new_n769_));
  INV_X1    g568(.A(G57gat), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n769_), .A2(new_n770_), .A3(new_n670_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n768_), .A2(new_n771_), .ZN(G1332gat));
  INV_X1    g571(.A(G64gat), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n773_), .B1(new_n766_), .B2(new_n429_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(KEYINPUT114), .B(KEYINPUT48), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n774_), .B(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n769_), .A2(new_n773_), .A3(new_n429_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(G1333gat));
  INV_X1    g577(.A(G71gat), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n779_), .B1(new_n766_), .B2(new_n570_), .ZN(new_n780_));
  XOR2_X1   g579(.A(new_n780_), .B(KEYINPUT49), .Z(new_n781_));
  NAND3_X1  g580(.A1(new_n769_), .A2(new_n779_), .A3(new_n570_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(G1334gat));
  INV_X1    g582(.A(G78gat), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n784_), .B1(new_n766_), .B2(new_n529_), .ZN(new_n785_));
  XOR2_X1   g584(.A(new_n785_), .B(KEYINPUT50), .Z(new_n786_));
  NAND3_X1  g585(.A1(new_n769_), .A2(new_n784_), .A3(new_n529_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT115), .ZN(G1335gat));
  NOR4_X1   g588(.A1(new_n620_), .A2(new_n633_), .A3(new_n680_), .A4(new_n703_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT116), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n669_), .A2(G85gat), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n667_), .A2(new_n634_), .A3(new_n302_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n793_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(new_n486_), .ZN(new_n795_));
  AOI22_X1  g594(.A1(new_n791_), .A2(new_n792_), .B1(G85gat), .B2(new_n795_), .ZN(new_n796_));
  XOR2_X1   g595(.A(new_n796_), .B(KEYINPUT117), .Z(G1336gat));
  INV_X1    g596(.A(G92gat), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n791_), .A2(new_n798_), .A3(new_n429_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n794_), .A2(new_n429_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n799_), .B1(new_n800_), .B2(new_n798_), .ZN(G1337gat));
  INV_X1    g600(.A(new_n560_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n237_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n791_), .A2(new_n802_), .A3(new_n803_), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n794_), .A2(new_n570_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n804_), .B1(new_n805_), .B2(new_n217_), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n806_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g606(.A1(new_n791_), .A2(new_n218_), .A3(new_n529_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n794_), .A2(new_n529_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(G106gat), .ZN(new_n810_));
  AND2_X1   g609(.A1(new_n810_), .A2(KEYINPUT52), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n810_), .A2(KEYINPUT52), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n808_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n813_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g613(.A1(new_n661_), .A2(new_n654_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n644_), .A2(new_n641_), .A3(new_n646_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n648_), .A2(KEYINPUT55), .A3(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n654_), .B1(new_n660_), .B2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n817_), .A2(KEYINPUT56), .A3(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(KEYINPUT56), .B1(new_n817_), .B2(new_n819_), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n633_), .B(new_n815_), .C1(new_n821_), .C2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n624_), .A2(new_n621_), .A3(new_n626_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n630_), .B1(new_n625_), .B2(new_n622_), .ZN(new_n825_));
  AOI22_X1  g624(.A1(new_n627_), .A2(new_n630_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(new_n658_), .B2(new_n662_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n702_), .B1(new_n823_), .B2(new_n827_), .ZN(new_n828_));
  OR2_X1    g627(.A1(new_n828_), .A2(KEYINPUT57), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n817_), .A2(new_n819_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT56), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  AOI22_X1  g631(.A1(new_n832_), .A2(new_n820_), .B1(new_n661_), .B2(new_n654_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n826_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT58), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n833_), .A2(KEYINPUT58), .A3(new_n826_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n836_), .A2(new_n837_), .A3(new_n275_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n828_), .A2(KEYINPUT57), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n829_), .A2(new_n838_), .A3(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n303_), .B1(new_n840_), .B2(KEYINPUT119), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT119), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n829_), .A2(new_n838_), .A3(new_n842_), .A4(new_n839_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT118), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n844_), .B1(new_n667_), .B2(new_n765_), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n663_), .A2(KEYINPUT118), .A3(new_n666_), .A4(new_n764_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n276_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(KEYINPUT54), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT54), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n847_), .A2(new_n850_), .A3(new_n276_), .ZN(new_n851_));
  AOI22_X1  g650(.A1(new_n841_), .A2(new_n843_), .B1(new_n849_), .B2(new_n851_), .ZN(new_n852_));
  OR4_X1    g651(.A1(new_n529_), .A2(new_n429_), .A3(new_n560_), .A4(new_n669_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(KEYINPUT120), .ZN(new_n854_));
  OAI21_X1  g653(.A(KEYINPUT121), .B1(new_n852_), .B2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n837_), .A2(new_n275_), .ZN(new_n856_));
  AOI21_X1  g655(.A(KEYINPUT58), .B1(new_n833_), .B2(new_n826_), .ZN(new_n857_));
  OAI22_X1  g656(.A1(new_n856_), .A2(new_n857_), .B1(new_n828_), .B2(KEYINPUT57), .ZN(new_n858_));
  INV_X1    g657(.A(new_n839_), .ZN(new_n859_));
  OAI21_X1  g658(.A(KEYINPUT119), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n860_), .A2(new_n302_), .A3(new_n843_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n849_), .A2(new_n851_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n854_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT121), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  AND2_X1   g664(.A1(new_n855_), .A2(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n866_), .A2(new_n459_), .A3(new_n633_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n863_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT123), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n869_), .B(new_n302_), .C1(new_n858_), .C2(new_n859_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n862_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n869_), .B1(new_n840_), .B2(new_n302_), .ZN(new_n872_));
  OR2_X1    g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT59), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(KEYINPUT122), .ZN(new_n875_));
  OR2_X1    g674(.A1(new_n874_), .A2(KEYINPUT122), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n854_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n877_));
  AOI22_X1  g676(.A1(new_n868_), .A2(KEYINPUT59), .B1(new_n873_), .B2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n633_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n867_), .B1(new_n880_), .B2(new_n459_), .ZN(G1340gat));
  OAI21_X1  g680(.A(new_n457_), .B1(new_n680_), .B2(KEYINPUT60), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n866_), .B(new_n882_), .C1(KEYINPUT60), .C2(new_n457_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n878_), .A2(new_n667_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n883_), .B1(new_n885_), .B2(new_n457_), .ZN(G1341gat));
  OAI21_X1  g685(.A(new_n877_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n303_), .B(new_n887_), .C1(new_n863_), .C2(new_n874_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(G127gat), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n302_), .A2(G127gat), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n855_), .A2(new_n865_), .A3(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT124), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n889_), .A2(new_n891_), .A3(KEYINPUT124), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1342gat));
  NAND3_X1  g695(.A1(new_n866_), .A2(new_n452_), .A3(new_n702_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n878_), .A2(new_n275_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n897_), .B1(new_n899_), .B2(new_n452_), .ZN(G1343gat));
  NAND2_X1  g699(.A1(new_n861_), .A2(new_n862_), .ZN(new_n901_));
  NOR4_X1   g700(.A1(new_n429_), .A2(new_n570_), .A3(new_n528_), .A4(new_n669_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n903_), .A2(new_n634_), .ZN(new_n904_));
  XOR2_X1   g703(.A(KEYINPUT125), .B(G141gat), .Z(new_n905_));
  XNOR2_X1  g704(.A(new_n904_), .B(new_n905_), .ZN(G1344gat));
  NOR2_X1   g705(.A1(new_n903_), .A2(new_n680_), .ZN(new_n907_));
  XOR2_X1   g706(.A(new_n907_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g707(.A1(new_n903_), .A2(new_n302_), .ZN(new_n909_));
  XOR2_X1   g708(.A(KEYINPUT61), .B(G155gat), .Z(new_n910_));
  XNOR2_X1  g709(.A(new_n909_), .B(new_n910_), .ZN(G1346gat));
  OAI21_X1  g710(.A(G162gat), .B1(new_n903_), .B2(new_n276_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n702_), .A2(new_n444_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n903_), .B2(new_n913_), .ZN(G1347gat));
  NOR2_X1   g713(.A1(new_n571_), .A2(new_n670_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(new_n429_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n916_), .A2(new_n529_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n873_), .A2(new_n917_), .ZN(new_n918_));
  OAI21_X1  g717(.A(G169gat), .B1(new_n918_), .B2(new_n634_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n918_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n922_), .A2(new_n633_), .A3(new_n342_), .ZN(new_n923_));
  OAI211_X1 g722(.A(KEYINPUT62), .B(G169gat), .C1(new_n918_), .C2(new_n634_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n921_), .A2(new_n923_), .A3(new_n924_), .ZN(G1348gat));
  AOI21_X1  g724(.A(G176gat), .B1(new_n922_), .B2(new_n667_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n852_), .A2(new_n529_), .ZN(new_n927_));
  NOR3_X1   g726(.A1(new_n680_), .A2(new_n916_), .A3(new_n343_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n926_), .B1(new_n927_), .B2(new_n928_), .ZN(G1349gat));
  NAND4_X1  g728(.A1(new_n927_), .A2(new_n429_), .A3(new_n303_), .A4(new_n915_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n302_), .B1(new_n384_), .B2(new_n386_), .ZN(new_n931_));
  AOI22_X1  g730(.A1(new_n930_), .A2(new_n381_), .B1(new_n922_), .B2(new_n931_), .ZN(G1350gat));
  OAI21_X1  g731(.A(G190gat), .B1(new_n918_), .B2(new_n276_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n702_), .A2(new_n370_), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n933_), .B1(new_n918_), .B2(new_n934_), .ZN(G1351gat));
  AND3_X1   g734(.A1(new_n571_), .A2(new_n616_), .A3(new_n429_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n901_), .A2(new_n936_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n937_), .A2(new_n634_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(new_n313_), .ZN(G1352gat));
  NOR2_X1   g738(.A1(new_n937_), .A2(new_n680_), .ZN(new_n940_));
  MUX2_X1   g739(.A(G204gat), .B(new_n319_), .S(new_n940_), .Z(G1353gat));
  AND2_X1   g740(.A1(new_n901_), .A2(new_n936_), .ZN(new_n942_));
  INV_X1    g741(.A(KEYINPUT63), .ZN(new_n943_));
  INV_X1    g742(.A(G211gat), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n303_), .B1(new_n943_), .B2(new_n944_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(new_n945_), .B(KEYINPUT126), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n942_), .A2(new_n946_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n947_), .A2(KEYINPUT127), .ZN(new_n948_));
  INV_X1    g747(.A(KEYINPUT127), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n942_), .A2(new_n949_), .A3(new_n946_), .ZN(new_n950_));
  NAND4_X1  g749(.A1(new_n948_), .A2(new_n943_), .A3(new_n944_), .A4(new_n950_), .ZN(new_n951_));
  AND3_X1   g750(.A1(new_n942_), .A2(new_n949_), .A3(new_n946_), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n949_), .B1(new_n942_), .B2(new_n946_), .ZN(new_n953_));
  OAI22_X1  g752(.A1(new_n952_), .A2(new_n953_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n951_), .A2(new_n954_), .ZN(G1354gat));
  OR3_X1    g754(.A1(new_n937_), .A2(G218gat), .A3(new_n271_), .ZN(new_n956_));
  OAI21_X1  g755(.A(G218gat), .B1(new_n937_), .B2(new_n276_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n956_), .A2(new_n957_), .ZN(G1355gat));
endmodule


