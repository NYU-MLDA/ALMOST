//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 1 1 0 1 0 0 1 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 1 1 1 1 1 0 0 0 0 0 1 1 1 0 1 0 1 1 0 0 1 1 0 1 1 0 1 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n699_, new_n700_, new_n701_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n756_, new_n757_, new_n758_, new_n759_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n777_, new_n778_, new_n779_, new_n780_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n796_,
    new_n797_, new_n799_, new_n800_, new_n801_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n890_, new_n892_, new_n893_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n907_, new_n908_, new_n909_, new_n911_,
    new_n912_, new_n914_, new_n915_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n922_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n930_, new_n931_;
  INV_X1    g000(.A(KEYINPUT75), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT35), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT70), .ZN(new_n204_));
  INV_X1    g003(.A(G85gat), .ZN(new_n205_));
  INV_X1    g004(.A(G92gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G85gat), .A2(G92gat), .ZN(new_n208_));
  AND2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT8), .ZN(new_n210_));
  AND2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT6), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT6), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(G99gat), .A3(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT64), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n213_), .A2(new_n215_), .A3(KEYINPUT64), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT7), .ZN(new_n221_));
  INV_X1    g020(.A(G99gat), .ZN(new_n222_));
  INV_X1    g021(.A(G106gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n221_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n211_), .B1(new_n220_), .B2(new_n226_), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n213_), .A2(new_n215_), .ZN(new_n228_));
  OAI211_X1 g027(.A(KEYINPUT66), .B(new_n209_), .C1(new_n228_), .C2(new_n226_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT8), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n216_), .A2(new_n225_), .A3(new_n224_), .ZN(new_n231_));
  AOI21_X1  g030(.A(KEYINPUT66), .B1(new_n231_), .B2(new_n209_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n227_), .B1(new_n230_), .B2(new_n232_), .ZN(new_n233_));
  OR2_X1    g032(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n234_), .A2(new_n223_), .A3(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n207_), .A2(KEYINPUT9), .A3(new_n208_), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n208_), .A2(KEYINPUT9), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n236_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n240_), .A2(KEYINPUT65), .A3(new_n219_), .A4(new_n218_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT65), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n242_), .B1(new_n220_), .B2(new_n239_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n233_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G29gat), .B(G36gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G43gat), .B(G50gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT15), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n245_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n209_), .B1(new_n228_), .B2(new_n226_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT66), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n256_), .A2(KEYINPUT8), .A3(new_n229_), .ZN(new_n257_));
  AOI22_X1  g056(.A1(new_n257_), .A2(new_n227_), .B1(new_n243_), .B2(new_n241_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n253_), .B1(new_n258_), .B2(new_n248_), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n233_), .A2(new_n244_), .A3(new_n253_), .A4(new_n248_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n204_), .B(new_n252_), .C1(new_n259_), .C2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G232gat), .A2(G233gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT34), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n262_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n264_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n250_), .B1(new_n244_), .B2(new_n233_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n233_), .A2(new_n244_), .A3(new_n248_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT69), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n267_), .B1(new_n269_), .B2(new_n260_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n266_), .B1(new_n270_), .B2(new_n204_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n203_), .B1(new_n265_), .B2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n262_), .A2(new_n264_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n270_), .A2(new_n203_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n270_), .A2(new_n204_), .A3(new_n266_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n273_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  XOR2_X1   g075(.A(G190gat), .B(G218gat), .Z(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT71), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G134gat), .B(G162gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT36), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n272_), .A2(KEYINPUT73), .A3(new_n276_), .A4(new_n281_), .ZN(new_n282_));
  AND2_X1   g081(.A1(new_n282_), .A2(KEYINPUT37), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT36), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n280_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(KEYINPUT72), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  AND3_X1   g086(.A1(new_n273_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n288_));
  AOI21_X1  g087(.A(KEYINPUT35), .B1(new_n273_), .B2(new_n275_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n287_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT73), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n272_), .A2(new_n276_), .A3(new_n281_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n290_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n283_), .A2(new_n293_), .A3(KEYINPUT74), .ZN(new_n294_));
  INV_X1    g093(.A(new_n292_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n286_), .B1(new_n272_), .B2(new_n276_), .ZN(new_n296_));
  OR3_X1    g095(.A1(new_n295_), .A2(new_n296_), .A3(KEYINPUT37), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n294_), .A2(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(KEYINPUT74), .B1(new_n283_), .B2(new_n293_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n202_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n283_), .A2(new_n293_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT74), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n303_), .A2(KEYINPUT75), .A3(new_n294_), .A4(new_n297_), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n300_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(G1gat), .ZN(new_n306_));
  INV_X1    g105(.A(G8gat), .ZN(new_n307_));
  OAI21_X1  g106(.A(KEYINPUT14), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  AND2_X1   g107(.A1(new_n308_), .A2(KEYINPUT76), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n308_), .A2(KEYINPUT76), .ZN(new_n310_));
  XOR2_X1   g109(.A(G15gat), .B(G22gat), .Z(new_n311_));
  NOR3_X1   g110(.A1(new_n309_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(G1gat), .B(G8gat), .Z(new_n313_));
  OR2_X1    g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n312_), .A2(new_n313_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G57gat), .B(G64gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT11), .ZN(new_n318_));
  XOR2_X1   g117(.A(G71gat), .B(G78gat), .Z(new_n319_));
  NOR2_X1   g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  AND2_X1   g119(.A1(new_n318_), .A2(new_n319_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n317_), .A2(KEYINPUT11), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n320_), .B1(new_n321_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n316_), .B(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G231gat), .A2(G233gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT17), .ZN(new_n329_));
  XOR2_X1   g128(.A(G127gat), .B(G155gat), .Z(new_n330_));
  XNOR2_X1  g129(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G183gat), .B(G211gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  OR3_X1    g133(.A1(new_n328_), .A2(new_n329_), .A3(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(KEYINPUT17), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n328_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n335_), .A2(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n305_), .A2(new_n338_), .ZN(new_n339_));
  XOR2_X1   g138(.A(KEYINPUT104), .B(KEYINPUT27), .Z(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  XOR2_X1   g140(.A(G8gat), .B(G36gat), .Z(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT18), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G64gat), .B(G92gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT20), .ZN(new_n347_));
  INV_X1    g146(.A(G197gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(KEYINPUT88), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT88), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(G197gat), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n349_), .A2(new_n351_), .A3(G204gat), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT90), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT21), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n349_), .A2(new_n351_), .A3(KEYINPUT90), .A4(G204gat), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT89), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n357_), .B1(new_n348_), .B2(G204gat), .ZN(new_n358_));
  INV_X1    g157(.A(G204gat), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n359_), .A2(KEYINPUT89), .A3(G197gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n354_), .A2(new_n355_), .A3(new_n356_), .A4(new_n361_), .ZN(new_n362_));
  XOR2_X1   g161(.A(G211gat), .B(G218gat), .Z(new_n363_));
  NAND3_X1  g162(.A1(new_n349_), .A2(new_n351_), .A3(new_n359_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n355_), .B1(G197gat), .B2(G204gat), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n363_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n354_), .A2(new_n356_), .A3(new_n361_), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n363_), .A2(KEYINPUT21), .ZN(new_n368_));
  AOI22_X1  g167(.A1(new_n362_), .A2(new_n366_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  AND2_X1   g168(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n370_));
  NOR2_X1   g169(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n371_));
  OAI21_X1  g170(.A(G183gat), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT79), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  OAI211_X1 g173(.A(KEYINPUT79), .B(G183gat), .C1(new_n370_), .C2(new_n371_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT80), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(G190gat), .ZN(new_n377_));
  OR2_X1    g176(.A1(new_n377_), .A2(KEYINPUT26), .ZN(new_n378_));
  INV_X1    g177(.A(G183gat), .ZN(new_n379_));
  AOI22_X1  g178(.A1(new_n377_), .A2(KEYINPUT26), .B1(KEYINPUT25), .B2(new_n379_), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n374_), .A2(new_n375_), .A3(new_n378_), .A4(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT24), .ZN(new_n382_));
  INV_X1    g181(.A(G169gat), .ZN(new_n383_));
  INV_X1    g182(.A(G176gat), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n382_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G169gat), .A2(G176gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(KEYINPUT24), .ZN(new_n387_));
  NOR2_X1   g186(.A1(G169gat), .A2(G176gat), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n385_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT23), .ZN(new_n390_));
  NAND3_X1  g189(.A1(KEYINPUT81), .A2(G183gat), .A3(G190gat), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(KEYINPUT81), .B1(G183gat), .B2(G190gat), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n390_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G183gat), .A2(G190gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(KEYINPUT23), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n389_), .B1(new_n394_), .B2(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(KEYINPUT23), .B1(new_n392_), .B2(new_n393_), .ZN(new_n398_));
  OR2_X1    g197(.A1(G183gat), .A2(G190gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n395_), .A2(new_n390_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n398_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT82), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(G169gat), .ZN(new_n403_));
  AOI21_X1  g202(.A(G176gat), .B1(new_n403_), .B2(KEYINPUT22), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n383_), .A2(KEYINPUT22), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(new_n402_), .ZN(new_n406_));
  AOI22_X1  g205(.A1(new_n404_), .A2(new_n406_), .B1(G169gat), .B2(G176gat), .ZN(new_n407_));
  AOI22_X1  g206(.A1(new_n381_), .A2(new_n397_), .B1(new_n401_), .B2(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n347_), .B1(new_n369_), .B2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n362_), .A2(new_n366_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n367_), .A2(new_n368_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT22), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(G169gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n383_), .A2(KEYINPUT22), .ZN(new_n415_));
  AND3_X1   g214(.A1(new_n414_), .A2(new_n415_), .A3(KEYINPUT96), .ZN(new_n416_));
  AOI21_X1  g215(.A(KEYINPUT96), .B1(new_n414_), .B2(new_n415_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n384_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT81), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n395_), .A2(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(KEYINPUT23), .B1(new_n420_), .B2(new_n391_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n396_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n399_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  XOR2_X1   g222(.A(new_n386_), .B(KEYINPUT95), .Z(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n418_), .A2(new_n423_), .A3(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n389_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(KEYINPUT25), .B(G183gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(KEYINPUT26), .B(G190gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n427_), .A2(new_n400_), .A3(new_n398_), .A4(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n426_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n412_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n409_), .A2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n435_));
  AND2_X1   g234(.A1(G226gat), .A2(G233gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(KEYINPUT94), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n434_), .A2(KEYINPUT97), .A3(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT96), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n413_), .A2(G169gat), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n441_), .B1(new_n405_), .B2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n414_), .A2(new_n415_), .A3(KEYINPUT96), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n424_), .B1(new_n445_), .B2(new_n384_), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n398_), .A2(new_n400_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n389_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n448_));
  AOI22_X1  g247(.A1(new_n446_), .A2(new_n423_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n347_), .B1(new_n449_), .B2(new_n369_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n408_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(new_n412_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n450_), .A2(new_n437_), .A3(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n440_), .A2(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(KEYINPUT97), .B1(new_n434_), .B2(new_n439_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n346_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n434_), .A2(new_n439_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT97), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n459_), .A2(new_n345_), .A3(new_n440_), .A4(new_n453_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n341_), .B1(new_n456_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT27), .ZN(new_n462_));
  INV_X1    g261(.A(new_n437_), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n410_), .A2(new_n426_), .A3(new_n411_), .A4(new_n431_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT20), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n369_), .A2(new_n408_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n463_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n409_), .A2(new_n433_), .A3(new_n438_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n345_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT102), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n462_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n437_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n409_), .A2(new_n433_), .A3(new_n438_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n346_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(KEYINPUT102), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n471_), .A2(new_n475_), .A3(new_n460_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT103), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT103), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n471_), .A2(new_n475_), .A3(new_n460_), .A4(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n461_), .B1(new_n477_), .B2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT85), .ZN(new_n481_));
  INV_X1    g280(.A(G141gat), .ZN(new_n482_));
  INV_X1    g281(.A(G148gat), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n481_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT85), .B1(G141gat), .B2(G148gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  OR2_X1    g285(.A1(G155gat), .A2(G162gat), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT1), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G155gat), .A2(G162gat), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n487_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G141gat), .A2(G148gat), .ZN(new_n491_));
  NAND3_X1  g290(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n486_), .A2(new_n490_), .A3(new_n491_), .A4(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT3), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n494_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT2), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n491_), .A2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n495_), .A2(new_n497_), .A3(new_n498_), .A4(new_n499_), .ZN(new_n500_));
  AND2_X1   g299(.A1(new_n487_), .A2(new_n489_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n493_), .A2(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(KEYINPUT87), .B1(new_n503_), .B2(KEYINPUT29), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n412_), .A2(new_n504_), .ZN(new_n505_));
  AND2_X1   g304(.A1(KEYINPUT86), .A2(G228gat), .ZN(new_n506_));
  NOR2_X1   g305(.A1(KEYINPUT86), .A2(G228gat), .ZN(new_n507_));
  OAI21_X1  g306(.A(G233gat), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n505_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n492_), .A2(new_n491_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n510_), .B1(new_n485_), .B2(new_n484_), .ZN(new_n511_));
  AOI22_X1  g310(.A1(new_n511_), .A2(new_n490_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT29), .ZN(new_n513_));
  NOR3_X1   g312(.A1(new_n512_), .A2(KEYINPUT91), .A3(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT91), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n508_), .B1(new_n503_), .B2(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n514_), .B1(new_n504_), .B2(new_n516_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n509_), .B1(new_n517_), .B2(new_n369_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G78gat), .B(G106gat), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n509_), .B(new_n519_), .C1(new_n369_), .C2(new_n517_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(KEYINPUT92), .B1(new_n518_), .B2(new_n520_), .ZN(new_n524_));
  INV_X1    g323(.A(G50gat), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT28), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n526_), .B1(new_n503_), .B2(KEYINPUT29), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n512_), .A2(KEYINPUT28), .A3(new_n513_), .ZN(new_n528_));
  INV_X1    g327(.A(G22gat), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n527_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n529_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n525_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n532_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n534_), .A2(G50gat), .A3(new_n530_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n523_), .B1(new_n524_), .B2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n536_), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n538_), .A2(new_n521_), .A3(KEYINPUT92), .A4(new_n522_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n537_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G1gat), .B(G29gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(G85gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(KEYINPUT0), .B(G57gat), .ZN(new_n543_));
  XOR2_X1   g342(.A(new_n542_), .B(new_n543_), .Z(new_n544_));
  INV_X1    g343(.A(KEYINPUT4), .ZN(new_n545_));
  INV_X1    g344(.A(G134gat), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(G127gat), .ZN(new_n547_));
  INV_X1    g346(.A(G127gat), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(G134gat), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G113gat), .B(G120gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n503_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT99), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n551_), .A2(new_n547_), .A3(new_n549_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n551_), .B1(new_n547_), .B2(new_n549_), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n493_), .B(new_n502_), .C1(new_n555_), .C2(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n553_), .A2(new_n554_), .A3(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n503_), .A2(KEYINPUT99), .A3(new_n552_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n545_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n503_), .A2(new_n545_), .A3(new_n552_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n561_), .A2(G225gat), .A3(G233gat), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n560_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT100), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n558_), .A2(new_n559_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G225gat), .A2(G233gat), .ZN(new_n566_));
  AOI22_X1  g365(.A1(new_n563_), .A2(new_n564_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(KEYINPUT100), .B1(new_n560_), .B2(new_n562_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n544_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n565_), .A2(KEYINPUT4), .ZN(new_n570_));
  INV_X1    g369(.A(new_n562_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n570_), .A2(new_n564_), .A3(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n565_), .A2(new_n566_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n572_), .A2(new_n568_), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n544_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(KEYINPUT101), .B1(new_n569_), .B2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n567_), .A2(new_n544_), .A3(new_n568_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n574_), .A2(new_n575_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT101), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n578_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n540_), .B1(new_n577_), .B2(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(KEYINPUT105), .B1(new_n480_), .B2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n480_), .A2(KEYINPUT105), .A3(new_n582_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n540_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n456_), .A2(new_n460_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT98), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT33), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n570_), .A2(new_n566_), .A3(new_n561_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n566_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n544_), .B1(new_n565_), .B2(new_n592_), .ZN(new_n593_));
  AOI22_X1  g392(.A1(new_n578_), .A2(new_n590_), .B1(new_n591_), .B2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n456_), .A2(KEYINPUT98), .A3(new_n460_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n576_), .A2(KEYINPUT33), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n589_), .A2(new_n594_), .A3(new_n595_), .A4(new_n596_), .ZN(new_n597_));
  AND2_X1   g396(.A1(new_n345_), .A2(KEYINPUT32), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n598_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n459_), .A2(new_n440_), .A3(new_n453_), .ZN(new_n600_));
  OAI221_X1 g399(.A(new_n599_), .B1(new_n600_), .B2(new_n598_), .C1(new_n569_), .C2(new_n576_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n586_), .B1(new_n597_), .B2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n584_), .A2(new_n585_), .A3(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT84), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n408_), .B(KEYINPUT30), .Z(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(G227gat), .A2(G233gat), .ZN(new_n608_));
  INV_X1    g407(.A(G15gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(G71gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(new_n222_), .ZN(new_n612_));
  OR2_X1    g411(.A1(new_n607_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n607_), .A2(new_n612_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(KEYINPUT83), .B(G43gat), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n613_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n615_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n605_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n618_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n620_), .A2(KEYINPUT84), .A3(new_n616_), .ZN(new_n621_));
  XOR2_X1   g420(.A(new_n552_), .B(KEYINPUT31), .Z(new_n622_));
  NAND3_X1  g421(.A1(new_n619_), .A2(new_n621_), .A3(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n622_), .ZN(new_n624_));
  OAI211_X1 g423(.A(new_n605_), .B(new_n624_), .C1(new_n617_), .C2(new_n618_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n480_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n627_), .A2(new_n586_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n577_), .A2(new_n581_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n626_), .A2(new_n630_), .ZN(new_n631_));
  AOI22_X1  g430(.A1(new_n604_), .A2(new_n626_), .B1(new_n628_), .B2(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n258_), .A2(new_n325_), .ZN(new_n633_));
  OR2_X1    g432(.A1(new_n633_), .A2(KEYINPUT12), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n245_), .A2(new_n324_), .ZN(new_n635_));
  OAI21_X1  g434(.A(KEYINPUT12), .B1(new_n633_), .B2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(G230gat), .A2(G233gat), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n634_), .A2(new_n636_), .A3(new_n637_), .ZN(new_n638_));
  OAI211_X1 g437(.A(G230gat), .B(G233gat), .C1(new_n633_), .C2(new_n635_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(G120gat), .B(G148gat), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT5), .ZN(new_n641_));
  XNOR2_X1  g440(.A(G176gat), .B(G204gat), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n641_), .B(new_n642_), .Z(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n638_), .A2(new_n639_), .A3(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT67), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n644_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n647_), .A2(new_n648_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  XOR2_X1   g450(.A(KEYINPUT68), .B(KEYINPUT13), .Z(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT13), .ZN(new_n654_));
  OAI22_X1  g453(.A1(new_n649_), .A2(new_n650_), .B1(KEYINPUT68), .B2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n653_), .A2(new_n655_), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n316_), .B(new_n248_), .Z(new_n657_));
  AND3_X1   g456(.A1(new_n314_), .A2(new_n248_), .A3(new_n315_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n658_), .B1(new_n251_), .B2(new_n316_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(G229gat), .A2(G233gat), .ZN(new_n660_));
  MUX2_X1   g459(.A(new_n657_), .B(new_n659_), .S(new_n660_), .Z(new_n661_));
  XNOR2_X1  g460(.A(G113gat), .B(G141gat), .ZN(new_n662_));
  XNOR2_X1  g461(.A(G169gat), .B(G197gat), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n662_), .B(new_n663_), .Z(new_n664_));
  XNOR2_X1  g463(.A(new_n661_), .B(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n656_), .A2(new_n666_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n632_), .A2(new_n667_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n339_), .A2(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n669_), .A2(new_n306_), .A3(new_n630_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT38), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n631_), .A2(new_n628_), .ZN(new_n672_));
  AND3_X1   g471(.A1(new_n480_), .A2(KEYINPUT105), .A3(new_n582_), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n673_), .A2(new_n583_), .A3(new_n602_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n626_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n672_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n295_), .A2(new_n296_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n678_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT107), .ZN(new_n680_));
  INV_X1    g479(.A(new_n338_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT106), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n682_), .B1(new_n656_), .B2(new_n666_), .ZN(new_n683_));
  AOI211_X1 g482(.A(KEYINPUT106), .B(new_n665_), .C1(new_n653_), .C2(new_n655_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n681_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  NOR3_X1   g484(.A1(new_n680_), .A2(new_n629_), .A3(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n671_), .B1(new_n306_), .B2(new_n686_), .ZN(G1324gat));
  NOR2_X1   g486(.A1(new_n680_), .A2(new_n685_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n307_), .B1(new_n688_), .B2(new_n627_), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n689_), .B(KEYINPUT39), .Z(new_n690_));
  NAND3_X1  g489(.A1(new_n669_), .A2(new_n307_), .A3(new_n627_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT40), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n692_), .B(new_n693_), .ZN(G1325gat));
  AOI21_X1  g493(.A(new_n609_), .B1(new_n688_), .B2(new_n675_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT41), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n669_), .A2(new_n609_), .A3(new_n675_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(G1326gat));
  AOI21_X1  g497(.A(new_n529_), .B1(new_n688_), .B2(new_n586_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT42), .Z(new_n700_));
  NAND3_X1  g499(.A1(new_n669_), .A2(new_n529_), .A3(new_n586_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(G1327gat));
  NOR2_X1   g501(.A1(new_n678_), .A2(new_n681_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n668_), .A2(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(G29gat), .B1(new_n704_), .B2(new_n630_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT43), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n305_), .A2(KEYINPUT109), .A3(new_n706_), .A4(new_n676_), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n676_), .A2(new_n706_), .A3(new_n300_), .A4(new_n304_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT109), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n300_), .A2(new_n304_), .ZN(new_n711_));
  OAI21_X1  g510(.A(KEYINPUT43), .B1(new_n711_), .B2(new_n632_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n707_), .A2(new_n710_), .A3(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n338_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(KEYINPUT108), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT108), .ZN(new_n716_));
  OAI211_X1 g515(.A(new_n716_), .B(new_n338_), .C1(new_n683_), .C2(new_n684_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n713_), .A2(KEYINPUT44), .A3(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(KEYINPUT44), .B1(new_n713_), .B2(new_n718_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n630_), .A2(G29gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n705_), .B1(new_n721_), .B2(new_n722_), .ZN(G1328gat));
  INV_X1    g522(.A(G36gat), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n704_), .A2(new_n724_), .A3(new_n627_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT45), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n725_), .B(new_n726_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n712_), .B1(new_n709_), .B2(new_n708_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n708_), .A2(new_n709_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n718_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n713_), .A2(KEYINPUT44), .A3(new_n718_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n732_), .A2(new_n627_), .A3(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n727_), .B1(new_n734_), .B2(G36gat), .ZN(new_n735_));
  AOI21_X1  g534(.A(KEYINPUT111), .B1(new_n735_), .B2(KEYINPUT46), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT46), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n737_), .B1(new_n735_), .B2(KEYINPUT110), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT110), .ZN(new_n739_));
  AOI211_X1 g538(.A(new_n739_), .B(new_n727_), .C1(new_n734_), .C2(G36gat), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n736_), .B1(new_n738_), .B2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n727_), .ZN(new_n742_));
  NOR3_X1   g541(.A1(new_n719_), .A2(new_n720_), .A3(new_n480_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n742_), .B1(new_n743_), .B2(new_n724_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(new_n739_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n735_), .A2(KEYINPUT110), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n745_), .A2(KEYINPUT111), .A3(new_n737_), .A4(new_n746_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n741_), .A2(new_n747_), .ZN(G1329gat));
  AOI21_X1  g547(.A(G43gat), .B1(new_n704_), .B2(new_n675_), .ZN(new_n749_));
  XOR2_X1   g548(.A(new_n749_), .B(KEYINPUT113), .Z(new_n750_));
  AND2_X1   g549(.A1(new_n675_), .A2(G43gat), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n721_), .A2(KEYINPUT112), .A3(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(KEYINPUT112), .B1(new_n721_), .B2(new_n751_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n750_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g554(.A1(new_n704_), .A2(new_n525_), .A3(new_n586_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n721_), .A2(KEYINPUT114), .A3(new_n586_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(G50gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(KEYINPUT114), .B1(new_n721_), .B2(new_n586_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n756_), .B1(new_n758_), .B2(new_n759_), .ZN(G1331gat));
  NOR2_X1   g559(.A1(new_n656_), .A2(new_n666_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n632_), .A2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n339_), .A2(new_n763_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT115), .ZN(new_n765_));
  AOI21_X1  g564(.A(G57gat), .B1(new_n765_), .B2(new_n630_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT116), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n680_), .A2(new_n338_), .A3(new_n762_), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n630_), .A2(G57gat), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n767_), .B1(new_n768_), .B2(new_n769_), .ZN(G1332gat));
  INV_X1    g569(.A(G64gat), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n771_), .B1(new_n768_), .B2(new_n627_), .ZN(new_n772_));
  XOR2_X1   g571(.A(KEYINPUT117), .B(KEYINPUT48), .Z(new_n773_));
  XNOR2_X1  g572(.A(new_n772_), .B(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n765_), .A2(new_n771_), .A3(new_n627_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(G1333gat));
  INV_X1    g575(.A(G71gat), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n777_), .B1(new_n768_), .B2(new_n675_), .ZN(new_n778_));
  XOR2_X1   g577(.A(new_n778_), .B(KEYINPUT49), .Z(new_n779_));
  NAND3_X1  g578(.A1(new_n765_), .A2(new_n777_), .A3(new_n675_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(G1334gat));
  INV_X1    g580(.A(G78gat), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n782_), .B1(new_n768_), .B2(new_n586_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(KEYINPUT118), .B(KEYINPUT50), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n783_), .B(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n765_), .A2(new_n782_), .A3(new_n586_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(G1335gat));
  INV_X1    g586(.A(new_n713_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n761_), .A2(new_n338_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n205_), .B1(new_n790_), .B2(new_n630_), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n763_), .A2(new_n703_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n629_), .A2(G85gat), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n791_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  XOR2_X1   g593(.A(new_n794_), .B(KEYINPUT119), .Z(G1336gat));
  NAND3_X1  g594(.A1(new_n792_), .A2(new_n206_), .A3(new_n627_), .ZN(new_n796_));
  NOR3_X1   g595(.A1(new_n788_), .A2(new_n480_), .A3(new_n789_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n796_), .B1(new_n797_), .B2(new_n206_), .ZN(G1337gat));
  NAND4_X1  g597(.A1(new_n792_), .A2(new_n234_), .A3(new_n235_), .A4(new_n675_), .ZN(new_n799_));
  NOR3_X1   g598(.A1(new_n788_), .A2(new_n626_), .A3(new_n789_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n799_), .B1(new_n800_), .B2(new_n222_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n801_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND2_X1  g601(.A1(new_n790_), .A2(new_n586_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(G106gat), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(KEYINPUT120), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n223_), .B1(new_n790_), .B2(new_n586_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT120), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n806_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n805_), .A2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n804_), .A2(KEYINPUT120), .A3(new_n806_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n792_), .A2(new_n223_), .A3(new_n586_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(KEYINPUT53), .B1(new_n810_), .B2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n805_), .A2(new_n809_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n815_), .A2(new_n816_), .A3(new_n811_), .A4(new_n812_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n814_), .A2(new_n817_), .ZN(G1339gat));
  INV_X1    g617(.A(KEYINPUT122), .ZN(new_n819_));
  INV_X1    g618(.A(G113gat), .ZN(new_n820_));
  INV_X1    g619(.A(new_n656_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n821_), .A2(new_n666_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n711_), .A2(new_n681_), .A3(new_n822_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n823_), .B(KEYINPUT54), .ZN(new_n824_));
  INV_X1    g623(.A(new_n664_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n661_), .A2(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n659_), .A2(G229gat), .A3(G233gat), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n664_), .B1(new_n657_), .B2(new_n660_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n826_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n637_), .B1(new_n634_), .B2(new_n636_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT55), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n638_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n634_), .A2(new_n636_), .A3(KEYINPUT55), .A4(new_n637_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  AND3_X1   g633(.A1(new_n834_), .A2(KEYINPUT56), .A3(new_n643_), .ZN(new_n835_));
  AOI21_X1  g634(.A(KEYINPUT56), .B1(new_n834_), .B2(new_n643_), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n645_), .B(new_n829_), .C1(new_n835_), .C2(new_n836_), .ZN(new_n837_));
  XOR2_X1   g636(.A(new_n837_), .B(KEYINPUT58), .Z(new_n838_));
  NOR2_X1   g637(.A1(new_n711_), .A2(new_n838_), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n666_), .B(new_n645_), .C1(new_n835_), .C2(new_n836_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n651_), .A2(new_n829_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n677_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(KEYINPUT57), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n338_), .B1(new_n839_), .B2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n824_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT59), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n626_), .A2(new_n629_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n628_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n845_), .A2(new_n846_), .A3(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  AND3_X1   g650(.A1(new_n824_), .A2(KEYINPUT121), .A3(new_n844_), .ZN(new_n852_));
  AOI21_X1  g651(.A(KEYINPUT121), .B1(new_n824_), .B2(new_n844_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n849_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n851_), .B1(new_n854_), .B2(KEYINPUT59), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n820_), .B1(new_n855_), .B2(new_n666_), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n854_), .A2(G113gat), .A3(new_n665_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n819_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT121), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n845_), .A2(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n824_), .A2(KEYINPUT121), .A3(new_n844_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n848_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n666_), .B(new_n850_), .C1(new_n862_), .C2(new_n846_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(G113gat), .ZN(new_n864_));
  INV_X1    g663(.A(new_n857_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n864_), .A2(KEYINPUT122), .A3(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n858_), .A2(new_n866_), .ZN(G1340gat));
  INV_X1    g666(.A(G120gat), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n868_), .B1(new_n656_), .B2(KEYINPUT60), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(KEYINPUT123), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n870_), .B1(KEYINPUT60), .B2(new_n868_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n854_), .A2(new_n871_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(KEYINPUT124), .ZN(new_n873_));
  INV_X1    g672(.A(new_n855_), .ZN(new_n874_));
  OAI21_X1  g673(.A(G120gat), .B1(new_n874_), .B2(new_n656_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n875_), .ZN(G1341gat));
  OAI21_X1  g675(.A(new_n548_), .B1(new_n854_), .B2(new_n338_), .ZN(new_n877_));
  OR2_X1    g676(.A1(new_n877_), .A2(KEYINPUT125), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(KEYINPUT125), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n855_), .A2(G127gat), .A3(new_n681_), .ZN(new_n880_));
  AND3_X1   g679(.A1(new_n878_), .A2(new_n879_), .A3(new_n880_), .ZN(G1342gat));
  OAI21_X1  g680(.A(G134gat), .B1(new_n874_), .B2(new_n711_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n862_), .A2(new_n546_), .A3(new_n677_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(G1343gat));
  NAND2_X1  g683(.A1(new_n860_), .A2(new_n861_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n675_), .A2(new_n629_), .A3(new_n540_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n885_), .A2(new_n480_), .A3(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n887_), .A2(new_n665_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(new_n482_), .ZN(G1344gat));
  NOR2_X1   g688(.A1(new_n887_), .A2(new_n656_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(new_n483_), .ZN(G1345gat));
  NOR2_X1   g690(.A1(new_n887_), .A2(new_n338_), .ZN(new_n892_));
  XOR2_X1   g691(.A(KEYINPUT61), .B(G155gat), .Z(new_n893_));
  XNOR2_X1  g692(.A(new_n892_), .B(new_n893_), .ZN(G1346gat));
  OAI21_X1  g693(.A(G162gat), .B1(new_n887_), .B2(new_n711_), .ZN(new_n895_));
  OR2_X1    g694(.A1(new_n678_), .A2(G162gat), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n887_), .B2(new_n896_), .ZN(G1347gat));
  NAND2_X1  g696(.A1(new_n631_), .A2(new_n627_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(new_n586_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n845_), .A2(new_n899_), .ZN(new_n900_));
  OAI21_X1  g699(.A(G169gat), .B1(new_n900_), .B2(new_n665_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n901_), .A2(KEYINPUT62), .ZN(new_n902_));
  AND2_X1   g701(.A1(new_n901_), .A2(KEYINPUT62), .ZN(new_n903_));
  INV_X1    g702(.A(new_n900_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n904_), .A2(new_n445_), .A3(new_n666_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n902_), .B1(new_n903_), .B2(new_n905_), .ZN(G1348gat));
  AOI21_X1  g705(.A(G176gat), .B1(new_n904_), .B2(new_n821_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n586_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n908_));
  NOR3_X1   g707(.A1(new_n898_), .A2(new_n384_), .A3(new_n656_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n907_), .B1(new_n908_), .B2(new_n909_), .ZN(G1349gat));
  NOR3_X1   g709(.A1(new_n900_), .A2(new_n428_), .A3(new_n338_), .ZN(new_n911_));
  NAND4_X1  g710(.A1(new_n908_), .A2(new_n627_), .A3(new_n631_), .A4(new_n681_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n911_), .B1(new_n912_), .B2(new_n379_), .ZN(G1350gat));
  OAI21_X1  g712(.A(G190gat), .B1(new_n900_), .B2(new_n711_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n677_), .A2(new_n429_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n914_), .B1(new_n900_), .B2(new_n915_), .ZN(G1351gat));
  NAND3_X1  g715(.A1(new_n627_), .A2(new_n626_), .A3(new_n582_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n917_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n918_));
  AOI22_X1  g717(.A1(new_n918_), .A2(new_n666_), .B1(KEYINPUT126), .B2(G197gat), .ZN(new_n919_));
  NOR2_X1   g718(.A1(KEYINPUT126), .A2(G197gat), .ZN(new_n920_));
  XOR2_X1   g719(.A(new_n919_), .B(new_n920_), .Z(G1352gat));
  NAND2_X1  g720(.A1(new_n918_), .A2(new_n821_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(G204gat), .ZN(G1353gat));
  AND2_X1   g722(.A1(new_n918_), .A2(new_n681_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n925_));
  AND2_X1   g724(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n924_), .B1(new_n925_), .B2(new_n926_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n927_), .B1(new_n924_), .B2(new_n925_), .ZN(G1354gat));
  AOI21_X1  g727(.A(G218gat), .B1(new_n918_), .B2(new_n677_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n305_), .A2(G218gat), .ZN(new_n930_));
  XOR2_X1   g729(.A(new_n930_), .B(KEYINPUT127), .Z(new_n931_));
  AOI21_X1  g730(.A(new_n929_), .B1(new_n918_), .B2(new_n931_), .ZN(G1355gat));
endmodule


