//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 0 1 1 0 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 0 0 0 1 0 0 0 1 0 1 1 1 0 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n699_,
    new_n700_, new_n701_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n719_, new_n720_,
    new_n721_, new_n723_, new_n724_, new_n725_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n739_, new_n740_, new_n741_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n857_, new_n859_,
    new_n860_, new_n861_, new_n863_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n909_, new_n910_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n917_, new_n918_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_;
  AND2_X1   g000(.A1(G57gat), .A2(G64gat), .ZN(new_n202_));
  NOR2_X1   g001(.A1(G57gat), .A2(G64gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT68), .B1(new_n202_), .B2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G57gat), .ZN(new_n205_));
  INV_X1    g004(.A(G64gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT68), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G57gat), .A2(G64gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT11), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n204_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G71gat), .ZN(new_n213_));
  INV_X1    g012(.A(G78gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G71gat), .A2(G78gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n212_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT69), .ZN(new_n218_));
  AND2_X1   g017(.A1(new_n204_), .A2(new_n210_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n219_), .A2(new_n211_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT69), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n212_), .A2(new_n221_), .A3(new_n215_), .A4(new_n216_), .ZN(new_n222_));
  AND3_X1   g021(.A1(new_n218_), .A2(new_n220_), .A3(new_n222_), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n220_), .B1(new_n218_), .B2(new_n222_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NOR3_X1   g026(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT6), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT65), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT65), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT6), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G99gat), .A2(G106gat), .ZN(new_n234_));
  AND3_X1   g033(.A1(new_n231_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n234_), .B1(new_n231_), .B2(new_n233_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n229_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  OR2_X1    g036(.A1(G85gat), .A2(G92gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G85gat), .A2(G92gat), .ZN(new_n239_));
  AND2_X1   g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT66), .B(KEYINPUT8), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n237_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT67), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n237_), .A2(new_n240_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT8), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT67), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n237_), .A2(new_n246_), .A3(new_n240_), .A4(new_n241_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n243_), .A2(new_n245_), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n236_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n231_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n252_));
  OR2_X1    g051(.A1(new_n252_), .A2(KEYINPUT64), .ZN(new_n253_));
  NAND3_X1  g052(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(KEYINPUT64), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n253_), .A2(new_n238_), .A3(new_n254_), .A4(new_n255_), .ZN(new_n256_));
  XOR2_X1   g055(.A(KEYINPUT10), .B(G99gat), .Z(new_n257_));
  INV_X1    g056(.A(G106gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n251_), .A2(new_n256_), .A3(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT71), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT71), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n251_), .A2(new_n256_), .A3(new_n262_), .A4(new_n259_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n248_), .A2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n225_), .A2(new_n265_), .A3(KEYINPUT12), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n248_), .B(new_n260_), .C1(new_n223_), .C2(new_n224_), .ZN(new_n267_));
  AND2_X1   g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G230gat), .A2(G233gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n248_), .A2(new_n260_), .ZN(new_n270_));
  AOI21_X1  g069(.A(KEYINPUT12), .B1(new_n225_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT72), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  AOI211_X1 g072(.A(KEYINPUT72), .B(KEYINPUT12), .C1(new_n225_), .C2(new_n270_), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n268_), .B(new_n269_), .C1(new_n273_), .C2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n225_), .A2(new_n270_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(new_n267_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n269_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT70), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n277_), .A2(new_n281_), .A3(new_n278_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n275_), .A2(new_n280_), .A3(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G120gat), .B(G148gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G176gat), .B(G204gat), .ZN(new_n287_));
  XOR2_X1   g086(.A(new_n286_), .B(new_n287_), .Z(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n283_), .A2(new_n289_), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n275_), .A2(new_n280_), .A3(new_n282_), .A4(new_n288_), .ZN(new_n291_));
  AND3_X1   g090(.A1(new_n290_), .A2(KEYINPUT13), .A3(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(KEYINPUT13), .B1(new_n290_), .B2(new_n291_), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G29gat), .A2(G36gat), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(G29gat), .A2(G36gat), .ZN(new_n297_));
  OAI21_X1  g096(.A(G43gat), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(G29gat), .ZN(new_n299_));
  INV_X1    g098(.A(G36gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(G43gat), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n301_), .A2(new_n302_), .A3(new_n295_), .ZN(new_n303_));
  AND3_X1   g102(.A1(new_n298_), .A2(new_n303_), .A3(G50gat), .ZN(new_n304_));
  AOI21_X1  g103(.A(G50gat), .B1(new_n298_), .B2(new_n303_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT15), .ZN(new_n306_));
  NOR3_X1   g105(.A1(new_n304_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(G50gat), .ZN(new_n308_));
  NOR3_X1   g107(.A1(new_n296_), .A2(new_n297_), .A3(G43gat), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n302_), .B1(new_n301_), .B2(new_n295_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n308_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n298_), .A2(new_n303_), .A3(G50gat), .ZN(new_n312_));
  AOI21_X1  g111(.A(KEYINPUT15), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n307_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G15gat), .B(G22gat), .ZN(new_n316_));
  INV_X1    g115(.A(G1gat), .ZN(new_n317_));
  INV_X1    g116(.A(G8gat), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT14), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n316_), .A2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G1gat), .B(G8gat), .ZN(new_n321_));
  OR2_X1    g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n321_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n315_), .A2(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n304_), .A2(new_n305_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n326_), .A2(new_n323_), .A3(new_n322_), .ZN(new_n327_));
  AND2_X1   g126(.A1(new_n325_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G229gat), .A2(G233gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  XOR2_X1   g129(.A(new_n324_), .B(new_n326_), .Z(new_n331_));
  NAND3_X1  g130(.A1(new_n331_), .A2(G229gat), .A3(G233gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G113gat), .B(G141gat), .ZN(new_n334_));
  INV_X1    g133(.A(G169gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(G197gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n333_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n338_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n330_), .A2(new_n332_), .A3(new_n340_), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n294_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G183gat), .A2(G190gat), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT23), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n346_), .B(new_n347_), .C1(G183gat), .C2(G190gat), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT83), .ZN(new_n349_));
  OR2_X1    g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n349_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(G169gat), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n350_), .A2(new_n351_), .A3(new_n353_), .ZN(new_n354_));
  XOR2_X1   g153(.A(G169gat), .B(G176gat), .Z(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT25), .B(G183gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT26), .B(G190gat), .ZN(new_n357_));
  AOI22_X1  g156(.A1(new_n355_), .A2(KEYINPUT24), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT24), .ZN(new_n359_));
  INV_X1    g158(.A(G176gat), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n359_), .A2(new_n335_), .A3(new_n360_), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n358_), .A2(new_n346_), .A3(new_n347_), .A4(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n354_), .A2(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(KEYINPUT85), .B(KEYINPUT31), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G127gat), .B(G134gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G113gat), .B(G120gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT84), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  OR2_X1    g169(.A1(new_n366_), .A2(new_n367_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(new_n368_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT84), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n370_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  XOR2_X1   g173(.A(G15gat), .B(G43gat), .Z(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  OR2_X1    g175(.A1(new_n365_), .A2(new_n376_), .ZN(new_n377_));
  XOR2_X1   g176(.A(G71gat), .B(G99gat), .Z(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT30), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G227gat), .A2(G233gat), .ZN(new_n380_));
  XOR2_X1   g179(.A(new_n379_), .B(new_n380_), .Z(new_n381_));
  NAND2_X1  g180(.A1(new_n365_), .A2(new_n376_), .ZN(new_n382_));
  AND3_X1   g181(.A1(new_n377_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n381_), .B1(new_n377_), .B2(new_n382_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(G155gat), .A2(G162gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT86), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G155gat), .A2(G162gat), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT1), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n387_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(G141gat), .ZN(new_n392_));
  INV_X1    g191(.A(G148gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G141gat), .A2(G148gat), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n391_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n394_), .B1(KEYINPUT87), .B2(KEYINPUT3), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n395_), .A2(KEYINPUT88), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT2), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT2), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n395_), .A2(KEYINPUT88), .A3(new_n400_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(KEYINPUT87), .A2(KEYINPUT3), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n402_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n397_), .A2(new_n399_), .A3(new_n401_), .A4(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n404_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n396_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(KEYINPUT29), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G197gat), .B(G204gat), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT21), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  XOR2_X1   g209(.A(G211gat), .B(G218gat), .Z(new_n411_));
  NOR2_X1   g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n408_), .A2(new_n409_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n408_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n415_), .A2(new_n411_), .A3(KEYINPUT21), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n416_), .A2(KEYINPUT91), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT91), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n418_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n414_), .B1(new_n417_), .B2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G228gat), .A2(G233gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(KEYINPUT90), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n407_), .A2(new_n420_), .A3(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT92), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n420_), .A2(new_n424_), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n414_), .B(KEYINPUT92), .C1(new_n417_), .C2(new_n419_), .ZN(new_n426_));
  AOI22_X1  g225(.A1(new_n425_), .A2(new_n426_), .B1(KEYINPUT29), .B2(new_n406_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n423_), .B1(new_n427_), .B2(new_n422_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G22gat), .B(G50gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  OR2_X1    g229(.A1(new_n406_), .A2(KEYINPUT29), .ZN(new_n431_));
  XOR2_X1   g230(.A(G78gat), .B(G106gat), .Z(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT89), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT28), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n431_), .B(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n429_), .ZN(new_n436_));
  OAI211_X1 g235(.A(new_n436_), .B(new_n423_), .C1(new_n427_), .C2(new_n422_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n430_), .A2(new_n435_), .A3(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n435_), .B1(new_n430_), .B2(new_n437_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(KEYINPUT4), .B1(new_n374_), .B2(new_n406_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n374_), .A2(new_n406_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT95), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n372_), .A2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n371_), .A2(KEYINPUT95), .A3(new_n368_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n445_), .A2(new_n396_), .A3(new_n405_), .A4(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n443_), .A2(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n442_), .B1(new_n448_), .B2(KEYINPUT4), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G225gat), .A2(G233gat), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n449_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n448_), .A2(new_n450_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G1gat), .B(G29gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G57gat), .B(G85gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n452_), .A2(new_n453_), .A3(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT99), .ZN(new_n460_));
  INV_X1    g259(.A(new_n453_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n461_), .B1(new_n451_), .B2(new_n449_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT99), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n462_), .A2(new_n463_), .A3(new_n458_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n458_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n452_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n465_), .B1(new_n466_), .B2(new_n461_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n460_), .A2(new_n464_), .A3(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(G226gat), .A2(G233gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n469_), .B(KEYINPUT19), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n361_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n471_));
  OR2_X1    g270(.A1(new_n471_), .A2(KEYINPUT93), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(KEYINPUT93), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n472_), .A2(new_n358_), .A3(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n353_), .A2(new_n348_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n420_), .A2(new_n476_), .ZN(new_n477_));
  AND2_X1   g276(.A1(KEYINPUT98), .A2(KEYINPUT20), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n479_), .B1(KEYINPUT98), .B2(KEYINPUT20), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n425_), .A2(new_n426_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(new_n363_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n470_), .B1(new_n480_), .B2(new_n483_), .ZN(new_n484_));
  AND2_X1   g283(.A1(new_n354_), .A2(new_n362_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n425_), .A2(new_n426_), .A3(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n420_), .A2(new_n476_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n486_), .A2(KEYINPUT20), .A3(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n484_), .B1(new_n470_), .B2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G8gat), .B(G36gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT18), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(G64gat), .ZN(new_n492_));
  INV_X1    g291(.A(G92gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  AND2_X1   g293(.A1(new_n494_), .A2(KEYINPUT32), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n489_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n488_), .A2(new_n470_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT20), .ZN(new_n498_));
  NOR3_X1   g297(.A1(new_n477_), .A2(new_n498_), .A3(new_n470_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(new_n482_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n497_), .A2(new_n500_), .ZN(new_n501_));
  OR2_X1    g300(.A1(new_n501_), .A2(new_n495_), .ZN(new_n502_));
  AND3_X1   g301(.A1(new_n468_), .A2(new_n496_), .A3(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n494_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n501_), .A2(KEYINPUT94), .A3(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT94), .ZN(new_n506_));
  AOI22_X1  g305(.A1(new_n488_), .A2(new_n470_), .B1(new_n499_), .B2(new_n482_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n506_), .B1(new_n507_), .B2(new_n494_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n494_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n458_), .B1(new_n448_), .B2(new_n450_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT97), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT97), .ZN(new_n512_));
  OAI211_X1 g311(.A(new_n512_), .B(new_n458_), .C1(new_n448_), .C2(new_n450_), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n511_), .B(new_n513_), .C1(new_n451_), .C2(new_n449_), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n505_), .A2(new_n508_), .A3(new_n509_), .A4(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT33), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n516_), .B1(new_n462_), .B2(new_n458_), .ZN(new_n517_));
  OAI211_X1 g316(.A(KEYINPUT33), .B(new_n465_), .C1(new_n466_), .C2(new_n461_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n515_), .A2(new_n519_), .ZN(new_n520_));
  OAI211_X1 g319(.A(new_n385_), .B(new_n441_), .C1(new_n503_), .C2(new_n520_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n385_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n377_), .A2(new_n382_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n381_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n377_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n440_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n527_), .A2(new_n528_), .A3(new_n438_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n522_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n468_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n505_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT27), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n504_), .A2(KEYINPUT100), .ZN(new_n535_));
  OR2_X1    g334(.A1(new_n504_), .A2(KEYINPUT100), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n489_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n509_), .A2(KEYINPUT101), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n533_), .B1(new_n509_), .B2(KEYINPUT101), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n537_), .A2(new_n538_), .A3(new_n539_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n530_), .A2(new_n531_), .A3(new_n534_), .A4(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n521_), .A2(new_n541_), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n343_), .A2(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n314_), .B1(new_n248_), .B2(new_n264_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT75), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G232gat), .A2(G233gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(KEYINPUT34), .ZN(new_n548_));
  XNOR2_X1  g347(.A(KEYINPUT74), .B(KEYINPUT35), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n548_), .A2(new_n549_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n248_), .A2(new_n326_), .A3(new_n260_), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n546_), .A2(new_n550_), .A3(new_n551_), .A4(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n545_), .B1(new_n265_), .B2(new_n315_), .ZN(new_n554_));
  AOI211_X1 g353(.A(KEYINPUT75), .B(new_n314_), .C1(new_n248_), .C2(new_n264_), .ZN(new_n555_));
  OAI211_X1 g354(.A(new_n551_), .B(new_n552_), .C1(new_n554_), .C2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n550_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G190gat), .B(G218gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT76), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(G134gat), .ZN(new_n561_));
  INV_X1    g360(.A(G162gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT36), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT77), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n563_), .A2(KEYINPUT77), .A3(new_n564_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n553_), .A2(new_n558_), .A3(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT78), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n553_), .A2(new_n558_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n563_), .B(new_n564_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n573_), .A2(new_n575_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n553_), .A2(new_n558_), .A3(KEYINPUT78), .A4(new_n569_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n572_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(KEYINPUT37), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT37), .ZN(new_n580_));
  AOI21_X1  g379(.A(KEYINPUT79), .B1(new_n573_), .B2(new_n575_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT79), .ZN(new_n582_));
  AOI211_X1 g381(.A(new_n582_), .B(new_n574_), .C1(new_n553_), .C2(new_n558_), .ZN(new_n583_));
  OAI211_X1 g382(.A(new_n580_), .B(new_n570_), .C1(new_n581_), .C2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n579_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(G231gat), .ZN(new_n587_));
  INV_X1    g386(.A(G233gat), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n324_), .A2(new_n589_), .ZN(new_n590_));
  OAI211_X1 g389(.A(new_n322_), .B(new_n323_), .C1(new_n587_), .C2(new_n588_), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n224_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n218_), .A2(new_n220_), .A3(new_n222_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n592_), .A2(new_n593_), .A3(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n590_), .A2(new_n591_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n596_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  XOR2_X1   g397(.A(G183gat), .B(G211gat), .Z(new_n599_));
  XNOR2_X1  g398(.A(G127gat), .B(G155gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(KEYINPUT17), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n598_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(KEYINPUT81), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT81), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n598_), .A2(new_n608_), .A3(new_n605_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n607_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n603_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT17), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n595_), .A2(new_n613_), .A3(new_n597_), .A4(new_n604_), .ZN(new_n614_));
  AOI21_X1  g413(.A(KEYINPUT82), .B1(new_n610_), .B2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT82), .ZN(new_n616_));
  INV_X1    g415(.A(new_n614_), .ZN(new_n617_));
  AOI211_X1 g416(.A(new_n616_), .B(new_n617_), .C1(new_n607_), .C2(new_n609_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n615_), .A2(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n586_), .A2(new_n619_), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n543_), .A2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n621_), .A2(new_n317_), .A3(new_n468_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT38), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n610_), .A2(new_n614_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n581_), .A2(new_n583_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n626_), .A2(new_n570_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT102), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n543_), .A2(new_n625_), .A3(new_n628_), .ZN(new_n629_));
  OAI21_X1  g428(.A(G1gat), .B1(new_n629_), .B2(new_n531_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n623_), .A2(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT103), .ZN(G1324gat));
  NAND2_X1  g431(.A1(new_n540_), .A2(new_n534_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  OAI21_X1  g433(.A(G8gat), .B1(new_n629_), .B2(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n635_), .B1(KEYINPUT104), .B2(KEYINPUT39), .ZN(new_n636_));
  NOR2_X1   g435(.A1(KEYINPUT104), .A2(KEYINPUT39), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n621_), .A2(new_n318_), .A3(new_n633_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT40), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n640_), .B(new_n641_), .ZN(G1325gat));
  OAI21_X1  g441(.A(G15gat), .B1(new_n629_), .B2(new_n385_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(KEYINPUT105), .B(KEYINPUT41), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n643_), .B(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(G15gat), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n621_), .A2(new_n646_), .A3(new_n527_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(G1326gat));
  XNOR2_X1  g447(.A(new_n441_), .B(KEYINPUT106), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n543_), .A2(new_n628_), .A3(new_n625_), .A4(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(G22gat), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT42), .ZN(new_n652_));
  INV_X1    g451(.A(G22gat), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n621_), .A2(new_n653_), .A3(new_n649_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n652_), .A2(new_n654_), .ZN(G1327gat));
  NAND2_X1  g454(.A1(new_n627_), .A2(new_n619_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n543_), .A2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n658_), .A2(new_n299_), .A3(new_n468_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n585_), .B(KEYINPUT109), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT108), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n521_), .A2(new_n662_), .A3(new_n541_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n662_), .B1(new_n521_), .B2(new_n541_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n660_), .B1(new_n661_), .B2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT43), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n586_), .A2(new_n542_), .A3(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  OAI211_X1 g468(.A(new_n343_), .B(new_n619_), .C1(new_n666_), .C2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n660_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT109), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n585_), .B(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n542_), .A2(KEYINPUT108), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n521_), .A2(new_n662_), .A3(new_n541_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n673_), .B1(new_n675_), .B2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(new_n668_), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n680_), .A2(KEYINPUT44), .A3(new_n343_), .A4(new_n619_), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n672_), .A2(new_n468_), .A3(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n659_), .B1(new_n682_), .B2(new_n299_), .ZN(G1328gat));
  XNOR2_X1  g482(.A(KEYINPUT111), .B(KEYINPUT46), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n672_), .A2(new_n633_), .A3(new_n681_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(G36gat), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(KEYINPUT110), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT110), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n685_), .A2(new_n688_), .A3(G36gat), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n689_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n658_), .A2(new_n300_), .A3(new_n633_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT45), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n684_), .B1(new_n690_), .B2(new_n692_), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n685_), .A2(new_n688_), .A3(G36gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n688_), .B1(new_n685_), .B2(G36gat), .ZN(new_n695_));
  OAI211_X1 g494(.A(new_n684_), .B(new_n692_), .C1(new_n694_), .C2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n693_), .A2(new_n697_), .ZN(G1329gat));
  NAND3_X1  g497(.A1(new_n658_), .A2(new_n302_), .A3(new_n527_), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n672_), .A2(new_n527_), .A3(new_n681_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n699_), .B1(new_n700_), .B2(new_n302_), .ZN(new_n701_));
  XOR2_X1   g500(.A(new_n701_), .B(KEYINPUT47), .Z(G1330gat));
  NAND3_X1  g501(.A1(new_n658_), .A2(new_n308_), .A3(new_n649_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n441_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n672_), .A2(new_n704_), .A3(new_n681_), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n705_), .A2(KEYINPUT112), .A3(G50gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(KEYINPUT112), .B1(new_n705_), .B2(G50gat), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n703_), .B1(new_n706_), .B2(new_n707_), .ZN(G1331gat));
  NOR2_X1   g507(.A1(new_n292_), .A2(new_n293_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n342_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n711_), .A2(new_n542_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n712_), .A2(new_n620_), .ZN(new_n713_));
  AOI21_X1  g512(.A(G57gat), .B1(new_n713_), .B2(new_n468_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n619_), .ZN(new_n715_));
  AND3_X1   g514(.A1(new_n628_), .A2(new_n715_), .A3(new_n712_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n531_), .A2(new_n205_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n714_), .B1(new_n716_), .B2(new_n717_), .ZN(G1332gat));
  AOI21_X1  g517(.A(new_n206_), .B1(new_n716_), .B2(new_n633_), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT48), .Z(new_n720_));
  NAND3_X1  g519(.A1(new_n713_), .A2(new_n206_), .A3(new_n633_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1333gat));
  AOI21_X1  g521(.A(new_n213_), .B1(new_n716_), .B2(new_n527_), .ZN(new_n723_));
  XOR2_X1   g522(.A(new_n723_), .B(KEYINPUT49), .Z(new_n724_));
  NAND3_X1  g523(.A1(new_n713_), .A2(new_n213_), .A3(new_n527_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(G1334gat));
  AOI21_X1  g525(.A(new_n214_), .B1(new_n716_), .B2(new_n649_), .ZN(new_n727_));
  XOR2_X1   g526(.A(new_n727_), .B(KEYINPUT50), .Z(new_n728_));
  NAND3_X1  g527(.A1(new_n713_), .A2(new_n214_), .A3(new_n649_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(G1335gat));
  AOI21_X1  g529(.A(new_n715_), .B1(new_n679_), .B2(new_n668_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(new_n711_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n468_), .A2(G85gat), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n733_), .B(KEYINPUT113), .Z(new_n734_));
  AND2_X1   g533(.A1(new_n712_), .A2(new_n657_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n735_), .A2(new_n468_), .ZN(new_n736_));
  OAI22_X1  g535(.A1(new_n732_), .A2(new_n734_), .B1(G85gat), .B2(new_n736_), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n737_), .B(KEYINPUT114), .Z(G1336gat));
  AOI21_X1  g537(.A(G92gat), .B1(new_n735_), .B2(new_n633_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n732_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n634_), .A2(new_n493_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n739_), .B1(new_n740_), .B2(new_n741_), .ZN(G1337gat));
  OAI21_X1  g541(.A(G99gat), .B1(new_n732_), .B2(new_n385_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n735_), .A2(new_n257_), .A3(new_n527_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND2_X1  g545(.A1(new_n740_), .A2(new_n704_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(G106gat), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT115), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT52), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n748_), .A2(new_n749_), .A3(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n735_), .A2(new_n258_), .A3(new_n704_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(KEYINPUT115), .A2(KEYINPUT52), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n749_), .A2(new_n750_), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n747_), .A2(G106gat), .A3(new_n753_), .A4(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n751_), .A2(new_n752_), .A3(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT53), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT53), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n751_), .A2(new_n758_), .A3(new_n752_), .A4(new_n755_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(G1339gat));
  NAND2_X1  g559(.A1(new_n275_), .A2(KEYINPUT118), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(KEYINPUT55), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n271_), .B(new_n272_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n269_), .B1(new_n763_), .B2(new_n268_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT55), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n275_), .A2(KEYINPUT118), .A3(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n762_), .A2(new_n765_), .A3(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(new_n289_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT56), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n331_), .A2(new_n329_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n328_), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n338_), .B(new_n771_), .C1(new_n772_), .C2(new_n329_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(new_n341_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT56), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n768_), .A2(new_n776_), .A3(new_n289_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n770_), .A2(new_n291_), .A3(new_n775_), .A4(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT58), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n774_), .B1(new_n769_), .B2(KEYINPUT56), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n781_), .A2(KEYINPUT58), .A3(new_n291_), .A4(new_n777_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n780_), .A2(new_n586_), .A3(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT57), .ZN(new_n784_));
  NOR2_X1   g583(.A1(KEYINPUT119), .A2(KEYINPUT56), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n275_), .A2(KEYINPUT118), .A3(new_n766_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n766_), .B1(new_n275_), .B2(KEYINPUT118), .ZN(new_n788_));
  NOR3_X1   g587(.A1(new_n787_), .A2(new_n788_), .A3(new_n764_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n786_), .B1(new_n789_), .B2(new_n288_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n768_), .A2(new_n289_), .A3(new_n785_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n790_), .A2(new_n710_), .A3(new_n291_), .A4(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n290_), .A2(new_n291_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(new_n775_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n626_), .A2(new_n570_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n784_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  AOI211_X1 g596(.A(KEYINPUT57), .B(new_n627_), .C1(new_n792_), .C2(new_n794_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n783_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n624_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n342_), .B1(new_n615_), .B2(new_n618_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT116), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  OAI211_X1 g602(.A(KEYINPUT116), .B(new_n342_), .C1(new_n615_), .C2(new_n618_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n585_), .A2(new_n709_), .A3(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(KEYINPUT117), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT117), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n585_), .A2(new_n709_), .A3(new_n805_), .A4(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n807_), .A2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT54), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n807_), .A2(KEYINPUT54), .A3(new_n809_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n800_), .A2(new_n814_), .ZN(new_n815_));
  NOR3_X1   g614(.A1(new_n633_), .A2(new_n531_), .A3(new_n529_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(G113gat), .B1(new_n818_), .B2(new_n710_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n817_), .A2(KEYINPUT59), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n799_), .A2(new_n619_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n814_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT59), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n822_), .A2(new_n823_), .A3(new_n816_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n820_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n710_), .A2(G113gat), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n819_), .B1(new_n826_), .B2(new_n827_), .ZN(G1340gat));
  INV_X1    g627(.A(KEYINPUT120), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n829_), .B1(new_n825_), .B2(new_n709_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n820_), .A2(KEYINPUT120), .A3(new_n294_), .A4(new_n824_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n830_), .A2(G120gat), .A3(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(G120gat), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n833_), .B1(new_n709_), .B2(KEYINPUT60), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n818_), .B(new_n834_), .C1(KEYINPUT60), .C2(new_n833_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n832_), .A2(new_n835_), .ZN(G1341gat));
  INV_X1    g635(.A(G127gat), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n837_), .B1(new_n817_), .B2(new_n619_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n625_), .A2(G127gat), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n838_), .B1(new_n825_), .B2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT121), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  OAI211_X1 g641(.A(KEYINPUT121), .B(new_n838_), .C1(new_n825_), .C2(new_n839_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(G1342gat));
  INV_X1    g643(.A(new_n628_), .ZN(new_n845_));
  AOI21_X1  g644(.A(G134gat), .B1(new_n818_), .B2(new_n845_), .ZN(new_n846_));
  XOR2_X1   g645(.A(KEYINPUT122), .B(G134gat), .Z(new_n847_));
  NOR2_X1   g646(.A1(new_n585_), .A2(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n846_), .B1(new_n826_), .B2(new_n848_), .ZN(G1343gat));
  NAND2_X1  g648(.A1(new_n812_), .A2(new_n813_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n850_), .B1(new_n624_), .B2(new_n799_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n851_), .A2(new_n522_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n633_), .A2(new_n531_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n854_), .A2(new_n342_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(new_n392_), .ZN(G1344gat));
  NOR2_X1   g655(.A1(new_n854_), .A2(new_n709_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(new_n393_), .ZN(G1345gat));
  NOR2_X1   g657(.A1(new_n854_), .A2(new_n619_), .ZN(new_n859_));
  XOR2_X1   g658(.A(KEYINPUT61), .B(G155gat), .Z(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(KEYINPUT123), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n859_), .B(new_n861_), .ZN(G1346gat));
  NOR3_X1   g661(.A1(new_n854_), .A2(new_n562_), .A3(new_n675_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n854_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n845_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n863_), .B1(new_n562_), .B2(new_n865_), .ZN(G1347gat));
  INV_X1    g665(.A(KEYINPUT124), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n634_), .A2(new_n468_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n527_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n869_), .A2(new_n649_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n822_), .A2(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n867_), .B1(new_n871_), .B2(new_n342_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n822_), .A2(KEYINPUT124), .A3(new_n710_), .A4(new_n870_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n872_), .A2(G169gat), .A3(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(KEYINPUT62), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT62), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n872_), .A2(new_n876_), .A3(G169gat), .A4(new_n873_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n875_), .A2(new_n877_), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n822_), .A2(new_n870_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(KEYINPUT22), .B(G169gat), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n879_), .A2(new_n710_), .A3(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n878_), .A2(new_n881_), .ZN(G1348gat));
  INV_X1    g681(.A(KEYINPUT126), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n869_), .A2(new_n709_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT125), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n885_), .B1(new_n815_), .B2(new_n441_), .ZN(new_n886_));
  AOI211_X1 g685(.A(KEYINPUT125), .B(new_n704_), .C1(new_n800_), .C2(new_n814_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n884_), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(G176gat), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n879_), .A2(new_n360_), .A3(new_n294_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n883_), .B1(new_n889_), .B2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n884_), .ZN(new_n892_));
  OAI21_X1  g691(.A(KEYINPUT125), .B1(new_n851_), .B2(new_n704_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n795_), .A2(new_n796_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(KEYINPUT57), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n795_), .A2(new_n784_), .A3(new_n796_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n625_), .B1(new_n897_), .B2(new_n783_), .ZN(new_n898_));
  OAI211_X1 g697(.A(new_n885_), .B(new_n441_), .C1(new_n898_), .C2(new_n850_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n892_), .B1(new_n893_), .B2(new_n899_), .ZN(new_n900_));
  OAI211_X1 g699(.A(new_n883_), .B(new_n890_), .C1(new_n900_), .C2(new_n360_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n891_), .A2(new_n902_), .ZN(G1349gat));
  NOR3_X1   g702(.A1(new_n871_), .A2(new_n624_), .A3(new_n356_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n869_), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n715_), .B(new_n905_), .C1(new_n886_), .C2(new_n887_), .ZN(new_n906_));
  INV_X1    g705(.A(G183gat), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n904_), .B1(new_n906_), .B2(new_n907_), .ZN(G1350gat));
  NAND3_X1  g707(.A1(new_n879_), .A2(new_n357_), .A3(new_n845_), .ZN(new_n909_));
  OAI21_X1  g708(.A(G190gat), .B1(new_n871_), .B2(new_n585_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(G1351gat));
  NAND3_X1  g710(.A1(new_n852_), .A2(new_n710_), .A3(new_n868_), .ZN(new_n912_));
  OR3_X1    g711(.A1(new_n912_), .A2(KEYINPUT127), .A3(new_n337_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n337_), .ZN(new_n914_));
  OAI21_X1  g713(.A(KEYINPUT127), .B1(new_n912_), .B2(new_n337_), .ZN(new_n915_));
  AND3_X1   g714(.A1(new_n913_), .A2(new_n914_), .A3(new_n915_), .ZN(G1352gat));
  AND2_X1   g715(.A1(new_n852_), .A2(new_n868_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(new_n294_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(G204gat), .ZN(G1353gat));
  AND3_X1   g718(.A1(new_n852_), .A2(new_n625_), .A3(new_n868_), .ZN(new_n920_));
  NOR3_X1   g719(.A1(new_n920_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n921_));
  XOR2_X1   g720(.A(KEYINPUT63), .B(G211gat), .Z(new_n922_));
  AOI21_X1  g721(.A(new_n921_), .B1(new_n920_), .B2(new_n922_), .ZN(G1354gat));
  AOI21_X1  g722(.A(G218gat), .B1(new_n917_), .B2(new_n845_), .ZN(new_n924_));
  AND2_X1   g723(.A1(new_n586_), .A2(G218gat), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n924_), .B1(new_n917_), .B2(new_n925_), .ZN(G1355gat));
endmodule


