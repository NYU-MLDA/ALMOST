//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 0 0 0 1 1 1 1 1 0 0 1 1 1 1 1 1 1 0 1 0 0 0 0 1 0 1 1 1 0 1 1 0 0 0 0 0 1 1 1 0 1 1 1 0 1 1 0 1 0 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n663_, new_n664_, new_n665_, new_n667_,
    new_n668_, new_n669_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n787_, new_n788_, new_n789_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n803_, new_n805_,
    new_n806_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n843_, new_n844_, new_n846_, new_n847_,
    new_n848_, new_n850_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n861_, new_n862_,
    new_n863_, new_n864_;
  XOR2_X1   g000(.A(G113gat), .B(G120gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G127gat), .B(G134gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  NOR2_X1   g003(.A1(G141gat), .A2(G148gat), .ZN(new_n205_));
  NOR2_X1   g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206_));
  AND2_X1   g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT1), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n206_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(G155gat), .ZN(new_n210_));
  INV_X1    g009(.A(G162gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT1), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n205_), .B1(new_n209_), .B2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G141gat), .A2(G148gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT86), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT85), .B(KEYINPUT3), .ZN(new_n216_));
  OR2_X1    g015(.A1(G141gat), .A2(G148gat), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n215_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT3), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n219_), .A2(KEYINPUT85), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n219_), .A2(KEYINPUT85), .ZN(new_n221_));
  OAI211_X1 g020(.A(KEYINPUT86), .B(new_n205_), .C1(new_n220_), .C2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n214_), .A2(KEYINPUT2), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT2), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n224_), .A2(G141gat), .A3(G148gat), .ZN(new_n225_));
  AOI22_X1  g024(.A1(new_n223_), .A2(new_n225_), .B1(new_n217_), .B2(KEYINPUT3), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n218_), .A2(new_n222_), .A3(new_n226_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n207_), .A2(new_n206_), .ZN(new_n228_));
  AOI221_X4 g027(.A(KEYINPUT87), .B1(new_n213_), .B2(new_n214_), .C1(new_n227_), .C2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT87), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n227_), .A2(new_n228_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n213_), .A2(new_n214_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n230_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n204_), .B1(new_n229_), .B2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n231_), .A2(new_n232_), .ZN(new_n235_));
  OR2_X1    g034(.A1(new_n235_), .A2(new_n204_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n234_), .A2(KEYINPUT4), .A3(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT92), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n234_), .A2(KEYINPUT4), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT92), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n234_), .A2(new_n240_), .A3(KEYINPUT4), .A4(new_n236_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n238_), .A2(new_n239_), .A3(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G225gat), .A2(G233gat), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n244_), .B1(new_n234_), .B2(new_n236_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G1gat), .B(G29gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(G85gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT0), .B(G57gat), .ZN(new_n251_));
  XOR2_X1   g050(.A(new_n250_), .B(new_n251_), .Z(new_n252_));
  NAND2_X1  g051(.A1(new_n248_), .A2(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n246_), .B1(new_n242_), .B2(new_n244_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n252_), .ZN(new_n255_));
  AOI21_X1  g054(.A(KEYINPUT95), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n253_), .A2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n248_), .A2(KEYINPUT95), .A3(new_n252_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n257_), .A2(KEYINPUT96), .A3(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n258_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT96), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n229_), .A2(new_n233_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT29), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G22gat), .B(G50gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT28), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n265_), .B(new_n267_), .ZN(new_n268_));
  XOR2_X1   g067(.A(G78gat), .B(G106gat), .Z(new_n269_));
  NAND2_X1  g068(.A1(G228gat), .A2(G233gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G211gat), .B(G218gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT21), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G197gat), .B(G204gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n272_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n271_), .A2(KEYINPUT21), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n274_), .B1(new_n277_), .B2(new_n273_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  OAI211_X1 g078(.A(new_n270_), .B(new_n279_), .C1(new_n263_), .C2(new_n264_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n264_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n281_));
  OAI211_X1 g080(.A(G228gat), .B(G233gat), .C1(new_n281_), .C2(new_n278_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n269_), .B1(new_n280_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT88), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n268_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(KEYINPUT89), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT89), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n268_), .B(new_n287_), .C1(new_n283_), .C2(new_n284_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  AND3_X1   g088(.A1(new_n280_), .A2(new_n269_), .A3(new_n282_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n290_), .A2(new_n283_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n289_), .A2(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n291_), .B1(new_n286_), .B2(new_n288_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT27), .ZN(new_n295_));
  INV_X1    g094(.A(G183gat), .ZN(new_n296_));
  INV_X1    g095(.A(G190gat), .ZN(new_n297_));
  OR3_X1    g096(.A1(new_n296_), .A2(new_n297_), .A3(KEYINPUT23), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT23), .B1(new_n296_), .B2(new_n297_), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n299_), .A2(KEYINPUT82), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n299_), .A2(KEYINPUT82), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n298_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  XOR2_X1   g101(.A(KEYINPUT79), .B(G190gat), .Z(new_n303_));
  OAI21_X1  g102(.A(new_n302_), .B1(G183gat), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G169gat), .A2(G176gat), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(KEYINPUT22), .B(G169gat), .ZN(new_n307_));
  INV_X1    g106(.A(G176gat), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n306_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n304_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT80), .ZN(new_n311_));
  INV_X1    g110(.A(G169gat), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n311_), .A2(new_n312_), .A3(new_n308_), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT80), .B1(G169gat), .B2(G176gat), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n313_), .A2(KEYINPUT24), .A3(new_n305_), .A4(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT81), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n298_), .A2(new_n299_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(KEYINPUT25), .B(G183gat), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT26), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(G190gat), .ZN(new_n320_));
  OAI211_X1 g119(.A(new_n318_), .B(new_n320_), .C1(new_n303_), .C2(new_n319_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n313_), .A2(new_n314_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT24), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n316_), .A2(new_n317_), .A3(new_n321_), .A4(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n310_), .A2(new_n325_), .A3(new_n278_), .ZN(new_n326_));
  AND2_X1   g125(.A1(new_n324_), .A2(new_n315_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT26), .B(G190gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(new_n318_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n327_), .A2(new_n302_), .A3(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT90), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n327_), .A2(new_n302_), .A3(KEYINPUT90), .A4(new_n329_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n317_), .B1(G183gat), .B2(G190gat), .ZN(new_n334_));
  AOI22_X1  g133(.A1(new_n332_), .A2(new_n333_), .B1(new_n309_), .B2(new_n334_), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n326_), .B(KEYINPUT20), .C1(new_n335_), .C2(new_n278_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G226gat), .A2(G233gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT19), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n335_), .A2(new_n278_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n338_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT20), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n310_), .A2(new_n325_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n342_), .B1(new_n343_), .B2(new_n279_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n340_), .A2(new_n341_), .A3(new_n344_), .ZN(new_n345_));
  XOR2_X1   g144(.A(KEYINPUT91), .B(KEYINPUT18), .Z(new_n346_));
  XNOR2_X1  g145(.A(G8gat), .B(G36gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G64gat), .B(G92gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n339_), .A2(new_n345_), .A3(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n351_), .B1(new_n339_), .B2(new_n345_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n295_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n334_), .A2(new_n309_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n278_), .A2(new_n330_), .A3(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n341_), .B1(new_n344_), .B2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n336_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n358_), .B1(new_n359_), .B2(new_n341_), .ZN(new_n360_));
  OAI211_X1 g159(.A(KEYINPUT27), .B(new_n352_), .C1(new_n360_), .C2(new_n351_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n355_), .A2(new_n361_), .ZN(new_n362_));
  NOR3_X1   g161(.A1(new_n293_), .A2(new_n294_), .A3(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G227gat), .A2(G233gat), .ZN(new_n364_));
  INV_X1    g163(.A(G71gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n343_), .B(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G15gat), .B(G43gat), .ZN(new_n368_));
  INV_X1    g167(.A(G99gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(KEYINPUT83), .B(KEYINPUT30), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  OR2_X1    g172(.A1(new_n367_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n367_), .A2(new_n373_), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n374_), .A2(new_n375_), .A3(KEYINPUT84), .ZN(new_n376_));
  AOI21_X1  g175(.A(KEYINPUT84), .B1(new_n374_), .B2(new_n375_), .ZN(new_n377_));
  XOR2_X1   g176(.A(new_n204_), .B(KEYINPUT31), .Z(new_n378_));
  OR3_X1    g177(.A1(new_n376_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n376_), .A2(new_n378_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  AND4_X1   g181(.A1(new_n259_), .A2(new_n262_), .A3(new_n363_), .A4(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT33), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n253_), .A2(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n353_), .A2(new_n354_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n234_), .A2(new_n244_), .A3(new_n236_), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n255_), .B(new_n387_), .C1(new_n242_), .C2(new_n244_), .ZN(new_n388_));
  AND2_X1   g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n255_), .B1(new_n245_), .B2(new_n247_), .ZN(new_n390_));
  AOI21_X1  g189(.A(KEYINPUT93), .B1(new_n390_), .B2(KEYINPUT33), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT93), .ZN(new_n392_));
  NOR4_X1   g191(.A1(new_n254_), .A2(new_n392_), .A3(new_n384_), .A4(new_n255_), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n385_), .B(new_n389_), .C1(new_n391_), .C2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n351_), .A2(KEYINPUT32), .ZN(new_n395_));
  OR2_X1    g194(.A1(new_n360_), .A2(new_n395_), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n339_), .A2(new_n345_), .ZN(new_n397_));
  AOI21_X1  g196(.A(KEYINPUT94), .B1(new_n397_), .B2(new_n395_), .ZN(new_n398_));
  AND4_X1   g197(.A1(KEYINPUT94), .A2(new_n339_), .A3(new_n345_), .A4(new_n395_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n257_), .A2(new_n258_), .A3(new_n396_), .A4(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n394_), .A2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n289_), .B(new_n292_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n362_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n262_), .A2(new_n403_), .A3(new_n259_), .A4(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n405_), .A2(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n383_), .B1(new_n408_), .B2(new_n381_), .ZN(new_n409_));
  XOR2_X1   g208(.A(G1gat), .B(G8gat), .Z(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(KEYINPUT76), .ZN(new_n411_));
  OR2_X1    g210(.A1(G15gat), .A2(G22gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G15gat), .A2(G22gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G1gat), .A2(G8gat), .ZN(new_n414_));
  AOI22_X1  g213(.A1(new_n412_), .A2(new_n413_), .B1(KEYINPUT14), .B2(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n411_), .B(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G29gat), .B(G36gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(G50gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT73), .B(G43gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n416_), .A2(new_n420_), .ZN(new_n421_));
  XOR2_X1   g220(.A(new_n420_), .B(KEYINPUT15), .Z(new_n422_));
  AOI21_X1  g221(.A(new_n421_), .B1(new_n422_), .B2(new_n416_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G229gat), .A2(G233gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(KEYINPUT78), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n423_), .A2(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n416_), .B(new_n420_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n427_), .A2(G229gat), .A3(G233gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n426_), .A2(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G113gat), .B(G141gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G169gat), .B(G197gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n430_), .B(new_n431_), .ZN(new_n432_));
  OR2_X1    g231(.A1(new_n429_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n429_), .A2(new_n432_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G230gat), .A2(G233gat), .ZN(new_n437_));
  XOR2_X1   g236(.A(new_n437_), .B(KEYINPUT64), .Z(new_n438_));
  AND2_X1   g237(.A1(G85gat), .A2(G92gat), .ZN(new_n439_));
  NOR2_X1   g238(.A1(G85gat), .A2(G92gat), .ZN(new_n440_));
  OR2_X1    g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n441_), .A2(KEYINPUT8), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G99gat), .A2(G106gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(KEYINPUT6), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT6), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n445_), .A2(G99gat), .A3(G106gat), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n444_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT7), .ZN(new_n448_));
  INV_X1    g247(.A(G106gat), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n448_), .A2(new_n369_), .A3(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n442_), .B1(new_n447_), .B2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n444_), .A2(new_n446_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT67), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n452_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n447_), .A2(KEYINPUT67), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n441_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT8), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n453_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(KEYINPUT9), .B1(new_n439_), .B2(new_n440_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT65), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT9), .ZN(new_n463_));
  INV_X1    g262(.A(G85gat), .ZN(new_n464_));
  INV_X1    g263(.A(G92gat), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n463_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n461_), .A2(new_n462_), .A3(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n439_), .A2(KEYINPUT65), .A3(KEYINPUT9), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT66), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  XOR2_X1   g270(.A(KEYINPUT10), .B(G99gat), .Z(new_n472_));
  AOI21_X1  g271(.A(new_n447_), .B1(new_n449_), .B2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n467_), .A2(KEYINPUT66), .A3(new_n468_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n471_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT68), .B(G71gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(G78gat), .ZN(new_n477_));
  XOR2_X1   g276(.A(G57gat), .B(G64gat), .Z(new_n478_));
  INV_X1    g277(.A(KEYINPUT11), .ZN(new_n479_));
  OR2_X1    g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n479_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n477_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(G78gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n476_), .B(new_n483_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n478_), .A2(new_n479_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n482_), .A2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n460_), .A2(new_n475_), .A3(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(KEYINPUT69), .A2(KEYINPUT12), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n460_), .A2(new_n475_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n487_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT69), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT12), .ZN(new_n494_));
  AOI22_X1  g293(.A1(new_n491_), .A2(new_n492_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n493_), .A2(new_n494_), .ZN(new_n496_));
  AOI211_X1 g295(.A(new_n496_), .B(new_n487_), .C1(new_n460_), .C2(new_n475_), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n438_), .B(new_n490_), .C1(new_n495_), .C2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n491_), .A2(new_n492_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(new_n488_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n438_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(KEYINPUT5), .B(G176gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(G204gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G120gat), .B(G148gat), .ZN(new_n505_));
  XOR2_X1   g304(.A(new_n504_), .B(new_n505_), .Z(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n498_), .A2(new_n502_), .A3(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT70), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n507_), .B1(new_n498_), .B2(new_n502_), .ZN(new_n511_));
  AND2_X1   g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n510_), .A2(new_n511_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n514_), .A2(KEYINPUT13), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT13), .ZN(new_n516_));
  NOR3_X1   g315(.A1(new_n512_), .A2(new_n513_), .A3(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT71), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  NOR3_X1   g319(.A1(new_n409_), .A2(new_n436_), .A3(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G232gat), .A2(G233gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT35), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n422_), .A2(new_n491_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT74), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n491_), .A2(new_n420_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT75), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n531_), .B1(new_n525_), .B2(new_n524_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n527_), .B1(new_n529_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT36), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G190gat), .B(G218gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G134gat), .B(G162gat), .ZN(new_n537_));
  XOR2_X1   g336(.A(new_n536_), .B(new_n537_), .Z(new_n538_));
  NAND3_X1  g337(.A1(new_n529_), .A2(new_n532_), .A3(new_n527_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n534_), .A2(new_n535_), .A3(new_n538_), .A4(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT37), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n538_), .B(KEYINPUT36), .ZN(new_n542_));
  INV_X1    g341(.A(new_n539_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n542_), .B1(new_n543_), .B2(new_n533_), .ZN(new_n544_));
  AND3_X1   g343(.A1(new_n540_), .A2(new_n541_), .A3(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n541_), .B1(new_n540_), .B2(new_n544_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G231gat), .A2(G233gat), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n487_), .B(new_n548_), .Z(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(new_n416_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G127gat), .B(G155gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(G211gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(KEYINPUT16), .B(G183gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n555_), .A2(KEYINPUT77), .A3(KEYINPUT17), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n556_), .B1(KEYINPUT17), .B2(new_n555_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n551_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n550_), .A2(new_n556_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n547_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n521_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n262_), .A2(new_n259_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NOR3_X1   g364(.A1(new_n563_), .A2(G1gat), .A3(new_n565_), .ZN(new_n566_));
  XOR2_X1   g365(.A(new_n566_), .B(KEYINPUT38), .Z(new_n567_));
  INV_X1    g366(.A(new_n409_), .ZN(new_n568_));
  OR2_X1    g367(.A1(new_n518_), .A2(KEYINPUT71), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n518_), .A2(KEYINPUT71), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n436_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n540_), .A2(new_n544_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n573_), .A2(new_n561_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n568_), .A2(new_n571_), .A3(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(G1gat), .B1(new_n575_), .B2(new_n565_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT97), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n567_), .A2(new_n577_), .ZN(G1324gat));
  OAI21_X1  g377(.A(G8gat), .B1(new_n575_), .B2(new_n406_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(KEYINPUT98), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT98), .ZN(new_n581_));
  OAI211_X1 g380(.A(new_n581_), .B(G8gat), .C1(new_n575_), .C2(new_n406_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n580_), .A2(KEYINPUT39), .A3(new_n582_), .ZN(new_n583_));
  OR3_X1    g382(.A1(new_n563_), .A2(G8gat), .A3(new_n406_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT39), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n579_), .A2(KEYINPUT98), .A3(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n583_), .A2(new_n584_), .A3(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(G1325gat));
  OAI21_X1  g388(.A(G15gat), .B1(new_n575_), .B2(new_n381_), .ZN(new_n590_));
  XOR2_X1   g389(.A(KEYINPUT100), .B(KEYINPUT41), .Z(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n381_), .A2(G15gat), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n592_), .B1(new_n563_), .B2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT101), .ZN(G1326gat));
  OAI21_X1  g394(.A(G22gat), .B1(new_n575_), .B2(new_n404_), .ZN(new_n596_));
  XOR2_X1   g395(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n404_), .A2(G22gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT103), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n598_), .B1(new_n563_), .B2(new_n600_), .ZN(G1327gat));
  INV_X1    g400(.A(new_n547_), .ZN(new_n602_));
  OAI21_X1  g401(.A(KEYINPUT43), .B1(new_n409_), .B2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT43), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n382_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n605_));
  OAI211_X1 g404(.A(new_n604_), .B(new_n547_), .C1(new_n605_), .C2(new_n383_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n603_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n571_), .A2(new_n561_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(KEYINPUT44), .B1(new_n607_), .B2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT44), .ZN(new_n611_));
  AOI211_X1 g410(.A(new_n611_), .B(new_n608_), .C1(new_n603_), .C2(new_n606_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(new_n564_), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n614_), .A2(KEYINPUT104), .A3(G29gat), .ZN(new_n615_));
  AOI21_X1  g414(.A(KEYINPUT104), .B1(new_n614_), .B2(G29gat), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n572_), .A2(new_n560_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n521_), .A2(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n565_), .A2(G29gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT105), .ZN(new_n620_));
  OAI22_X1  g419(.A1(new_n615_), .A2(new_n616_), .B1(new_n618_), .B2(new_n620_), .ZN(G1328gat));
  INV_X1    g420(.A(KEYINPUT46), .ZN(new_n622_));
  NOR3_X1   g421(.A1(new_n610_), .A2(new_n612_), .A3(new_n406_), .ZN(new_n623_));
  INV_X1    g422(.A(G36gat), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NOR3_X1   g424(.A1(new_n618_), .A2(G36gat), .A3(new_n406_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT45), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n622_), .B1(new_n625_), .B2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT45), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n626_), .B(new_n629_), .ZN(new_n630_));
  OAI211_X1 g429(.A(new_n630_), .B(KEYINPUT46), .C1(new_n624_), .C2(new_n623_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n628_), .A2(new_n631_), .ZN(G1329gat));
  INV_X1    g431(.A(G43gat), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n633_), .B1(new_n618_), .B2(new_n381_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT107), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n381_), .A2(new_n633_), .ZN(new_n636_));
  AOI21_X1  g435(.A(KEYINPUT106), .B1(new_n613_), .B2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT106), .ZN(new_n638_));
  INV_X1    g437(.A(new_n636_), .ZN(new_n639_));
  NOR4_X1   g438(.A1(new_n610_), .A2(new_n612_), .A3(new_n638_), .A4(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n635_), .B1(new_n637_), .B2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(KEYINPUT47), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT47), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n643_), .B(new_n635_), .C1(new_n637_), .C2(new_n640_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n644_), .ZN(G1330gat));
  OR3_X1    g444(.A1(new_n618_), .A2(G50gat), .A3(new_n404_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n613_), .A2(new_n403_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT108), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n647_), .A2(new_n648_), .A3(G50gat), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n648_), .B1(new_n647_), .B2(G50gat), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n646_), .B1(new_n649_), .B2(new_n650_), .ZN(G1331gat));
  NAND4_X1  g450(.A1(new_n568_), .A2(new_n436_), .A3(new_n520_), .A4(new_n574_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  OAI21_X1  g452(.A(G57gat), .B1(new_n565_), .B2(KEYINPUT110), .ZN(new_n654_));
  OAI211_X1 g453(.A(new_n653_), .B(new_n654_), .C1(KEYINPUT110), .C2(G57gat), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n562_), .A2(new_n520_), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n656_), .A2(KEYINPUT109), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(KEYINPUT109), .ZN(new_n658_));
  NAND4_X1  g457(.A1(new_n657_), .A2(new_n436_), .A3(new_n568_), .A4(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n659_), .A2(new_n565_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n655_), .B1(new_n660_), .B2(G57gat), .ZN(new_n661_));
  XOR2_X1   g460(.A(new_n661_), .B(KEYINPUT111), .Z(G1332gat));
  OAI21_X1  g461(.A(G64gat), .B1(new_n652_), .B2(new_n406_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT48), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n406_), .A2(G64gat), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n664_), .B1(new_n659_), .B2(new_n665_), .ZN(G1333gat));
  OAI21_X1  g465(.A(G71gat), .B1(new_n652_), .B2(new_n381_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT49), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n659_), .A2(G71gat), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n668_), .B1(new_n381_), .B2(new_n669_), .ZN(G1334gat));
  OR3_X1    g469(.A1(new_n659_), .A2(G78gat), .A3(new_n404_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT50), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n653_), .A2(new_n403_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n672_), .B1(new_n673_), .B2(G78gat), .ZN(new_n674_));
  AOI211_X1 g473(.A(KEYINPUT50), .B(new_n483_), .C1(new_n653_), .C2(new_n403_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n671_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT112), .ZN(G1335gat));
  AND4_X1   g476(.A1(new_n436_), .A2(new_n568_), .A3(new_n520_), .A4(new_n617_), .ZN(new_n678_));
  AOI21_X1  g477(.A(G85gat), .B1(new_n678_), .B2(new_n564_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT113), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n520_), .A2(new_n436_), .A3(new_n561_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(KEYINPUT114), .B1(new_n607_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT114), .ZN(new_n684_));
  AOI211_X1 g483(.A(new_n684_), .B(new_n681_), .C1(new_n603_), .C2(new_n606_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n683_), .A2(new_n685_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n565_), .A2(new_n464_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n680_), .B1(new_n686_), .B2(new_n687_), .ZN(G1336gat));
  AOI21_X1  g487(.A(G92gat), .B1(new_n678_), .B2(new_n362_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n406_), .A2(new_n465_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n689_), .B1(new_n686_), .B2(new_n690_), .ZN(G1337gat));
  OR2_X1    g490(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n692_));
  NAND2_X1  g491(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n369_), .B1(new_n686_), .B2(new_n382_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n678_), .A2(new_n472_), .A3(new_n382_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n692_), .B(new_n693_), .C1(new_n694_), .C2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n683_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n685_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n698_), .A2(new_n699_), .A3(new_n382_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(G99gat), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n701_), .A2(KEYINPUT115), .A3(KEYINPUT51), .A4(new_n695_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n697_), .A2(new_n702_), .ZN(G1338gat));
  NAND3_X1  g502(.A1(new_n678_), .A2(new_n449_), .A3(new_n403_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT116), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n607_), .A2(new_n403_), .A3(new_n682_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n706_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(G106gat), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT52), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n705_), .A2(new_n707_), .A3(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT53), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT53), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n705_), .A2(new_n713_), .A3(new_n707_), .A4(new_n710_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n714_), .ZN(G1339gat));
  INV_X1    g514(.A(KEYINPUT54), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n515_), .A2(new_n517_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT117), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n717_), .A2(new_n718_), .A3(new_n436_), .A4(new_n560_), .ZN(new_n719_));
  OAI211_X1 g518(.A(new_n436_), .B(new_n560_), .C1(new_n515_), .C2(new_n517_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(KEYINPUT117), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n716_), .B1(new_n722_), .B2(new_n602_), .ZN(new_n723_));
  AOI211_X1 g522(.A(KEYINPUT54), .B(new_n547_), .C1(new_n719_), .C2(new_n721_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n435_), .A2(new_n508_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n498_), .A2(KEYINPUT118), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(KEYINPUT55), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n490_), .B1(new_n495_), .B2(new_n497_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(new_n501_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT55), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n498_), .A2(KEYINPUT118), .A3(new_n731_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n728_), .A2(new_n730_), .A3(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT119), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NAND4_X1  g534(.A1(new_n728_), .A2(new_n730_), .A3(KEYINPUT119), .A4(new_n732_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(KEYINPUT56), .B1(new_n737_), .B2(new_n506_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT56), .ZN(new_n739_));
  AOI211_X1 g538(.A(new_n739_), .B(new_n507_), .C1(new_n735_), .C2(new_n736_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n726_), .B1(new_n738_), .B2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT120), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n427_), .A2(new_n425_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n423_), .ZN(new_n745_));
  OAI211_X1 g544(.A(new_n432_), .B(new_n744_), .C1(new_n745_), .C2(new_n425_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n433_), .A2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(new_n514_), .ZN(new_n748_));
  OAI211_X1 g547(.A(KEYINPUT120), .B(new_n726_), .C1(new_n738_), .C2(new_n740_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n743_), .A2(new_n748_), .A3(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(new_n572_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT57), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n750_), .A2(KEYINPUT57), .A3(new_n572_), .ZN(new_n754_));
  OR2_X1    g553(.A1(new_n738_), .A2(new_n740_), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n755_), .A2(KEYINPUT58), .A3(new_n508_), .A4(new_n747_), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n508_), .B(new_n747_), .C1(new_n738_), .C2(new_n740_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT58), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n756_), .A2(new_n547_), .A3(new_n759_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n753_), .A2(new_n754_), .A3(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n725_), .B1(new_n761_), .B2(new_n561_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n564_), .A2(new_n382_), .A3(new_n363_), .ZN(new_n763_));
  XOR2_X1   g562(.A(new_n763_), .B(KEYINPUT121), .Z(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n762_), .A2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT59), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(KEYINPUT59), .B1(new_n762_), .B2(new_n765_), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n768_), .A2(new_n769_), .A3(G113gat), .A4(new_n435_), .ZN(new_n770_));
  INV_X1    g569(.A(G113gat), .ZN(new_n771_));
  AND3_X1   g570(.A1(new_n750_), .A2(KEYINPUT57), .A3(new_n572_), .ZN(new_n772_));
  AOI21_X1  g571(.A(KEYINPUT57), .B1(new_n750_), .B2(new_n572_), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n756_), .A2(new_n547_), .A3(new_n759_), .ZN(new_n774_));
  NOR3_X1   g573(.A1(new_n772_), .A2(new_n773_), .A3(new_n774_), .ZN(new_n775_));
  OAI22_X1  g574(.A1(new_n775_), .A2(new_n560_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n764_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n771_), .B1(new_n777_), .B2(new_n436_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n770_), .A2(new_n778_), .ZN(G1340gat));
  NAND3_X1  g578(.A1(new_n768_), .A2(new_n769_), .A3(new_n520_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(G120gat), .ZN(new_n781_));
  INV_X1    g580(.A(G120gat), .ZN(new_n782_));
  INV_X1    g581(.A(new_n520_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n782_), .B1(new_n783_), .B2(KEYINPUT60), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n766_), .B(new_n784_), .C1(KEYINPUT60), .C2(new_n782_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n781_), .A2(new_n785_), .ZN(G1341gat));
  AOI21_X1  g585(.A(G127gat), .B1(new_n766_), .B2(new_n560_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n768_), .A2(new_n769_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n560_), .A2(G127gat), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n787_), .B1(new_n788_), .B2(new_n789_), .ZN(G1342gat));
  INV_X1    g589(.A(G134gat), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n791_), .B1(new_n777_), .B2(new_n572_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT122), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n768_), .A2(new_n769_), .A3(G134gat), .A4(new_n547_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT122), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n795_), .B(new_n791_), .C1(new_n777_), .C2(new_n572_), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n793_), .A2(new_n794_), .A3(new_n796_), .ZN(G1343gat));
  NOR3_X1   g596(.A1(new_n565_), .A2(new_n404_), .A3(new_n362_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  NOR3_X1   g598(.A1(new_n762_), .A2(new_n382_), .A3(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n435_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n801_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n520_), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n803_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g603(.A1(new_n800_), .A2(new_n560_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(KEYINPUT61), .B(G155gat), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n805_), .B(new_n806_), .ZN(G1346gat));
  AOI21_X1  g606(.A(G162gat), .B1(new_n800_), .B2(new_n573_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n776_), .A2(G162gat), .A3(new_n381_), .A4(new_n798_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n809_), .A2(new_n602_), .ZN(new_n810_));
  OAI21_X1  g609(.A(KEYINPUT123), .B1(new_n808_), .B2(new_n810_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n776_), .A2(new_n381_), .A3(new_n573_), .A4(new_n798_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n211_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT123), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n813_), .B(new_n814_), .C1(new_n602_), .C2(new_n809_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n811_), .A2(new_n815_), .ZN(G1347gat));
  NOR2_X1   g615(.A1(new_n564_), .A2(new_n381_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n362_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n776_), .A2(new_n435_), .A3(new_n404_), .A4(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT62), .ZN(new_n821_));
  AND3_X1   g620(.A1(new_n820_), .A2(new_n821_), .A3(G169gat), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n821_), .B1(new_n820_), .B2(G169gat), .ZN(new_n823_));
  NOR3_X1   g622(.A1(new_n762_), .A2(new_n403_), .A3(new_n818_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n435_), .A2(new_n307_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n826_), .B(KEYINPUT124), .ZN(new_n827_));
  OAI22_X1  g626(.A1(new_n822_), .A2(new_n823_), .B1(new_n825_), .B2(new_n827_), .ZN(G1348gat));
  XOR2_X1   g627(.A(KEYINPUT125), .B(G176gat), .Z(new_n829_));
  OAI21_X1  g628(.A(new_n829_), .B1(new_n825_), .B2(new_n783_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n308_), .A2(KEYINPUT125), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n824_), .A2(new_n520_), .A3(new_n831_), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n830_), .A2(new_n832_), .ZN(G1349gat));
  AOI21_X1  g632(.A(new_n296_), .B1(new_n824_), .B2(new_n560_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n776_), .A2(new_n404_), .A3(new_n560_), .A4(new_n819_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n318_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(KEYINPUT126), .B1(new_n834_), .B2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n835_), .A2(G183gat), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT126), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n839_), .B(new_n840_), .C1(new_n836_), .C2(new_n835_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n838_), .A2(new_n841_), .ZN(G1350gat));
  OAI21_X1  g641(.A(G190gat), .B1(new_n825_), .B2(new_n602_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n824_), .A2(new_n328_), .A3(new_n573_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(G1351gat));
  NOR2_X1   g644(.A1(new_n762_), .A2(new_n382_), .ZN(new_n846_));
  NOR3_X1   g645(.A1(new_n564_), .A2(new_n404_), .A3(new_n406_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n846_), .A2(new_n435_), .A3(new_n847_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n848_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g648(.A1(new_n846_), .A2(new_n520_), .A3(new_n847_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g650(.A(KEYINPUT127), .ZN(new_n852_));
  AND4_X1   g651(.A1(new_n381_), .A2(new_n776_), .A3(new_n560_), .A4(new_n847_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n852_), .B1(new_n853_), .B2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n846_), .A2(new_n847_), .ZN(new_n857_));
  OAI211_X1 g656(.A(KEYINPUT127), .B(new_n854_), .C1(new_n857_), .C2(new_n561_), .ZN(new_n858_));
  XOR2_X1   g657(.A(KEYINPUT63), .B(G211gat), .Z(new_n859_));
  AOI22_X1  g658(.A1(new_n856_), .A2(new_n858_), .B1(new_n853_), .B2(new_n859_), .ZN(G1354gat));
  INV_X1    g659(.A(G218gat), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n857_), .A2(new_n861_), .A3(new_n602_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n857_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n573_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n862_), .B1(new_n861_), .B2(new_n864_), .ZN(G1355gat));
endmodule


