//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 0 1 0 0 0 1 1 1 1 1 1 1 1 0 1 0 1 1 1 1 0 1 1 1 0 1 1 1 1 0 1 1 1 0 1 0 0 0 1 0 0 0 0 1 0 0 0 1 1 1 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n659_, new_n660_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n824_, new_n825_, new_n827_, new_n828_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n873_, new_n874_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n897_;
  NOR3_X1   g000(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT66), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G99gat), .A2(G106gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT6), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G99gat), .ZN(new_n209_));
  INV_X1    g008(.A(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT7), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n204_), .A2(new_n208_), .A3(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G85gat), .ZN(new_n214_));
  INV_X1    g013(.A(G92gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G85gat), .A2(G92gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n213_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT67), .ZN(new_n221_));
  AOI21_X1  g020(.A(KEYINPUT8), .B1(new_n219_), .B2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT9), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT65), .ZN(new_n224_));
  AND3_X1   g023(.A1(new_n217_), .A2(new_n224_), .A3(new_n223_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n224_), .B1(new_n217_), .B2(new_n223_), .ZN(new_n226_));
  OAI221_X1 g025(.A(new_n216_), .B1(new_n223_), .B2(new_n217_), .C1(new_n225_), .C2(new_n226_), .ZN(new_n227_));
  XOR2_X1   g026(.A(KEYINPUT10), .B(G99gat), .Z(new_n228_));
  AOI21_X1  g027(.A(new_n207_), .B1(new_n210_), .B2(new_n228_), .ZN(new_n229_));
  AOI22_X1  g028(.A1(new_n220_), .A2(new_n222_), .B1(new_n227_), .B2(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n207_), .B1(KEYINPUT7), .B2(new_n211_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n218_), .B1(new_n231_), .B2(new_n204_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n222_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n230_), .A2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G57gat), .B(G64gat), .ZN(new_n236_));
  OR2_X1    g035(.A1(new_n236_), .A2(KEYINPUT11), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(KEYINPUT11), .ZN(new_n238_));
  XOR2_X1   g037(.A(G71gat), .B(G78gat), .Z(new_n239_));
  NAND3_X1  g038(.A1(new_n237_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  OR2_X1    g039(.A1(new_n238_), .A2(new_n239_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n235_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT69), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT12), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n244_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n242_), .B1(new_n230_), .B2(new_n234_), .ZN(new_n248_));
  OAI21_X1  g047(.A(KEYINPUT69), .B1(new_n248_), .B2(KEYINPUT12), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n235_), .A2(new_n243_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n229_), .A2(new_n227_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n252_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n220_), .A2(new_n222_), .ZN(new_n254_));
  OAI211_X1 g053(.A(KEYINPUT12), .B(new_n243_), .C1(new_n253_), .C2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT68), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n235_), .A2(new_n257_), .A3(KEYINPUT12), .A4(new_n243_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n251_), .B1(new_n256_), .B2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G230gat), .A2(G233gat), .ZN(new_n260_));
  XOR2_X1   g059(.A(new_n260_), .B(KEYINPUT64), .Z(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n250_), .A2(new_n259_), .A3(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n261_), .B1(new_n251_), .B2(new_n248_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  XOR2_X1   g064(.A(G120gat), .B(G148gat), .Z(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G176gat), .B(G204gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n265_), .A2(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n263_), .A2(new_n264_), .A3(new_n270_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n274_), .A2(KEYINPUT13), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(KEYINPUT13), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  XOR2_X1   g076(.A(new_n277_), .B(KEYINPUT71), .Z(new_n278_));
  XOR2_X1   g077(.A(G127gat), .B(G155gat), .Z(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G183gat), .B(G211gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G231gat), .A2(G233gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n242_), .B(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G1gat), .B(G8gat), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT72), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(G15gat), .ZN(new_n290_));
  INV_X1    g089(.A(G22gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G15gat), .A2(G22gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G1gat), .A2(G8gat), .ZN(new_n294_));
  AOI22_X1  g093(.A1(new_n292_), .A2(new_n293_), .B1(KEYINPUT14), .B2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n289_), .B(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n286_), .B(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT74), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n284_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n299_), .A2(KEYINPUT17), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT17), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n301_), .B1(new_n297_), .B2(new_n284_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n299_), .A2(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n300_), .A2(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G29gat), .B(G36gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G43gat), .B(G50gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT15), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n235_), .A2(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n230_), .A2(new_n307_), .A3(new_n234_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G232gat), .A2(G233gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT34), .ZN(new_n312_));
  OAI211_X1 g111(.A(new_n309_), .B(new_n310_), .C1(KEYINPUT35), .C2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(KEYINPUT35), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G190gat), .B(G218gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G134gat), .B(G162gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT36), .ZN(new_n319_));
  OR2_X1    g118(.A1(new_n315_), .A2(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n318_), .A2(KEYINPUT36), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n315_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT37), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT37), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n320_), .A2(new_n325_), .A3(new_n322_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n324_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NOR3_X1   g127(.A1(new_n278_), .A2(new_n304_), .A3(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n296_), .B(new_n307_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G229gat), .A2(G233gat), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n296_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(new_n308_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n296_), .A2(new_n307_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  OAI211_X1 g136(.A(new_n333_), .B(KEYINPUT75), .C1(new_n332_), .C2(new_n337_), .ZN(new_n338_));
  OR3_X1    g137(.A1(new_n337_), .A2(KEYINPUT75), .A3(new_n332_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G113gat), .B(G141gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G169gat), .B(G197gat), .ZN(new_n342_));
  XOR2_X1   g141(.A(new_n341_), .B(new_n342_), .Z(new_n343_));
  NAND2_X1  g142(.A1(new_n340_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n343_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n338_), .A2(new_n339_), .A3(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G183gat), .A2(G190gat), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT78), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(KEYINPUT78), .A2(G183gat), .A3(G190gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n349_), .B1(new_n354_), .B2(KEYINPUT23), .ZN(new_n355_));
  INV_X1    g154(.A(G183gat), .ZN(new_n356_));
  INV_X1    g155(.A(G190gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n355_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G169gat), .A2(G176gat), .ZN(new_n360_));
  INV_X1    g159(.A(G169gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT22), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT22), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(G169gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT79), .B(G176gat), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n360_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT80), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT80), .ZN(new_n369_));
  OAI211_X1 g168(.A(new_n369_), .B(new_n360_), .C1(new_n365_), .C2(new_n366_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n359_), .A2(new_n368_), .A3(new_n370_), .ZN(new_n371_));
  NOR3_X1   g170(.A1(KEYINPUT77), .A2(G169gat), .A3(G176gat), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT77), .B1(G169gat), .B2(G176gat), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n373_), .A2(KEYINPUT24), .A3(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n360_), .A2(KEYINPUT24), .ZN(new_n376_));
  INV_X1    g175(.A(new_n374_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n376_), .B1(new_n377_), .B2(new_n372_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n375_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT76), .ZN(new_n380_));
  OR3_X1    g179(.A1(new_n380_), .A2(new_n357_), .A3(KEYINPUT26), .ZN(new_n381_));
  XNOR2_X1  g180(.A(KEYINPUT25), .B(G183gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n357_), .A2(KEYINPUT26), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n380_), .B1(new_n357_), .B2(KEYINPUT26), .ZN(new_n384_));
  NAND4_X1  g183(.A1(new_n381_), .A2(new_n382_), .A3(new_n383_), .A4(new_n384_), .ZN(new_n385_));
  AND2_X1   g184(.A1(new_n350_), .A2(KEYINPUT23), .ZN(new_n386_));
  AOI21_X1  g185(.A(KEYINPUT23), .B1(new_n352_), .B2(new_n353_), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n379_), .B(new_n385_), .C1(new_n386_), .C2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n371_), .A2(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT30), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(KEYINPUT82), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT83), .ZN(new_n392_));
  XOR2_X1   g191(.A(G127gat), .B(G134gat), .Z(new_n393_));
  XOR2_X1   g192(.A(G113gat), .B(G120gat), .Z(new_n394_));
  XOR2_X1   g193(.A(new_n393_), .B(new_n394_), .Z(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT31), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n392_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n398_), .B1(new_n397_), .B2(new_n396_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n391_), .B(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G227gat), .A2(G233gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(G15gat), .ZN(new_n402_));
  XOR2_X1   g201(.A(KEYINPUT81), .B(G43gat), .Z(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G71gat), .B(G99gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n406_), .B1(new_n390_), .B2(KEYINPUT82), .ZN(new_n407_));
  XOR2_X1   g206(.A(new_n400_), .B(new_n407_), .Z(new_n408_));
  NOR2_X1   g207(.A1(G155gat), .A2(G162gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G155gat), .A2(G162gat), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n409_), .B1(KEYINPUT1), .B2(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n411_), .B1(KEYINPUT1), .B2(new_n410_), .ZN(new_n412_));
  XOR2_X1   g211(.A(G141gat), .B(G148gat), .Z(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT3), .ZN(new_n415_));
  INV_X1    g214(.A(G141gat), .ZN(new_n416_));
  INV_X1    g215(.A(G148gat), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n415_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G141gat), .A2(G148gat), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT2), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n418_), .A2(new_n421_), .A3(new_n422_), .A4(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT84), .ZN(new_n425_));
  XOR2_X1   g224(.A(G155gat), .B(G162gat), .Z(new_n426_));
  AND3_X1   g225(.A1(new_n424_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n425_), .B1(new_n424_), .B2(new_n426_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n414_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT85), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT85), .ZN(new_n431_));
  OAI211_X1 g230(.A(new_n431_), .B(new_n414_), .C1(new_n427_), .C2(new_n428_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n430_), .A2(new_n432_), .A3(new_n395_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT89), .ZN(new_n434_));
  INV_X1    g233(.A(new_n428_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n424_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n436_));
  AOI22_X1  g235(.A1(new_n435_), .A2(new_n436_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n434_), .B1(new_n437_), .B2(new_n396_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n433_), .A2(new_n438_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n430_), .A2(new_n434_), .A3(new_n432_), .A4(new_n395_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n439_), .A2(KEYINPUT4), .A3(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT4), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n433_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n441_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(G225gat), .A2(G233gat), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n444_), .A2(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G1gat), .B(G29gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(KEYINPUT91), .ZN(new_n449_));
  XOR2_X1   g248(.A(G57gat), .B(G85gat), .Z(new_n450_));
  XNOR2_X1  g249(.A(new_n449_), .B(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(KEYINPUT90), .B(KEYINPUT0), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n451_), .B(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n446_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n447_), .A2(new_n454_), .A3(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n445_), .B1(new_n441_), .B2(new_n443_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n453_), .B1(new_n458_), .B2(new_n455_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n457_), .A2(KEYINPUT92), .A3(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT92), .ZN(new_n461_));
  OAI211_X1 g260(.A(new_n461_), .B(new_n453_), .C1(new_n458_), .C2(new_n455_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G226gat), .A2(G233gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n358_), .B1(new_n387_), .B2(new_n386_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n365_), .A2(KEYINPUT88), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT88), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n362_), .A2(new_n364_), .A3(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n470_), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n467_), .B(new_n360_), .C1(new_n471_), .C2(new_n366_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(G197gat), .A2(G204gat), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G197gat), .A2(G204gat), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n474_), .A2(KEYINPUT21), .A3(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G211gat), .B(G218gat), .ZN(new_n477_));
  OR2_X1    g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT21), .ZN(new_n479_));
  INV_X1    g278(.A(new_n475_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n479_), .B1(new_n480_), .B2(new_n473_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n476_), .A2(new_n481_), .A3(new_n477_), .ZN(new_n482_));
  AND2_X1   g281(.A1(new_n478_), .A2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT26), .B(G190gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n382_), .A2(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n379_), .A2(new_n355_), .A3(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n472_), .A2(new_n483_), .A3(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT20), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n483_), .B1(new_n371_), .B2(new_n388_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n466_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n472_), .A2(new_n486_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n483_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n371_), .A2(new_n388_), .A3(new_n483_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n493_), .A2(new_n494_), .A3(KEYINPUT20), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n490_), .B1(new_n466_), .B2(new_n495_), .ZN(new_n496_));
  XOR2_X1   g295(.A(G8gat), .B(G36gat), .Z(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT18), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G64gat), .B(G92gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n496_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n495_), .A2(new_n466_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n489_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n466_), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n504_), .A2(KEYINPUT20), .A3(new_n505_), .A4(new_n487_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n503_), .A2(new_n506_), .A3(new_n500_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n502_), .A2(KEYINPUT27), .A3(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NOR3_X1   g308(.A1(new_n488_), .A2(new_n489_), .A3(new_n466_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT20), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n511_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n505_), .B1(new_n512_), .B2(new_n494_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n501_), .B1(new_n510_), .B2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(new_n507_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT27), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(KEYINPUT93), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT93), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n515_), .A2(new_n519_), .A3(new_n516_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n509_), .B1(new_n518_), .B2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G22gat), .B(G50gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n430_), .A2(new_n432_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT28), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT29), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n523_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n524_), .B1(new_n523_), .B2(new_n525_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n522_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n528_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n522_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n530_), .A2(new_n526_), .A3(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n529_), .A2(new_n532_), .ZN(new_n533_));
  XOR2_X1   g332(.A(G78gat), .B(G106gat), .Z(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n430_), .A2(KEYINPUT29), .A3(new_n432_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(KEYINPUT86), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT86), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n430_), .A2(new_n538_), .A3(KEYINPUT29), .A4(new_n432_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n537_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(G228gat), .ZN(new_n541_));
  INV_X1    g340(.A(G233gat), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n492_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n540_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n429_), .A2(KEYINPUT29), .ZN(new_n546_));
  AOI211_X1 g345(.A(new_n541_), .B(new_n542_), .C1(new_n546_), .C2(new_n492_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n535_), .B1(new_n545_), .B2(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n543_), .B1(new_n537_), .B2(new_n539_), .ZN(new_n550_));
  NOR3_X1   g349(.A1(new_n550_), .A2(new_n534_), .A3(new_n547_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n533_), .B1(new_n549_), .B2(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n545_), .A2(new_n535_), .A3(new_n548_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n534_), .B1(new_n550_), .B2(new_n547_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n553_), .A2(new_n554_), .A3(new_n532_), .A4(new_n529_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n552_), .A2(new_n555_), .ZN(new_n556_));
  AND3_X1   g355(.A1(new_n463_), .A2(new_n521_), .A3(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n500_), .A2(KEYINPUT32), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n558_), .B1(new_n510_), .B2(new_n513_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n559_), .B1(new_n558_), .B2(new_n496_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n460_), .A2(new_n462_), .A3(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT33), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n457_), .A2(new_n562_), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n447_), .A2(KEYINPUT33), .A3(new_n454_), .A4(new_n456_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n444_), .A2(new_n445_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n439_), .A2(new_n440_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n454_), .B1(new_n566_), .B2(new_n446_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n515_), .B1(new_n565_), .B2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n563_), .A2(new_n564_), .A3(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n556_), .B1(new_n561_), .B2(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n408_), .B1(new_n557_), .B2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n556_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT94), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n572_), .A2(new_n521_), .A3(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n519_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n575_));
  AOI211_X1 g374(.A(KEYINPUT93), .B(KEYINPUT27), .C1(new_n514_), .C2(new_n507_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n508_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  OAI21_X1  g376(.A(KEYINPUT94), .B1(new_n577_), .B2(new_n556_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n574_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n463_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n580_), .A2(new_n408_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n348_), .B1(new_n571_), .B2(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n583_), .A2(KEYINPUT95), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n583_), .A2(KEYINPUT95), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n329_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n586_), .A2(KEYINPUT96), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(KEYINPUT96), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n463_), .A2(G1gat), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n587_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT38), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n323_), .B(KEYINPUT97), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n594_), .B1(new_n571_), .B2(new_n582_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n277_), .A2(new_n347_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n596_), .A2(new_n304_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  OAI21_X1  g397(.A(G1gat), .B1(new_n598_), .B2(new_n463_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n590_), .A2(new_n591_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n592_), .A2(new_n599_), .A3(new_n600_), .ZN(G1324gat));
  NOR2_X1   g400(.A1(new_n521_), .A2(G8gat), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n587_), .A2(new_n588_), .A3(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(G8gat), .B1(new_n598_), .B2(new_n521_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT39), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n603_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT40), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n603_), .A2(KEYINPUT40), .A3(new_n605_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(G1325gat));
  OAI21_X1  g409(.A(G15gat), .B1(new_n598_), .B2(new_n408_), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT41), .Z(new_n612_));
  INV_X1    g411(.A(new_n586_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n408_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n613_), .A2(new_n290_), .A3(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n612_), .A2(new_n615_), .ZN(G1326gat));
  NAND3_X1  g415(.A1(new_n613_), .A2(new_n291_), .A3(new_n556_), .ZN(new_n617_));
  OAI21_X1  g416(.A(G22gat), .B1(new_n598_), .B2(new_n572_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT42), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT98), .ZN(G1327gat));
  OR2_X1    g420(.A1(new_n585_), .A2(new_n584_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n277_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n304_), .ZN(new_n624_));
  NOR3_X1   g423(.A1(new_n623_), .A2(new_n624_), .A3(new_n323_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n622_), .A2(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(G29gat), .B1(new_n626_), .B2(new_n580_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n596_), .A2(new_n624_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT43), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n571_), .A2(new_n582_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n629_), .B1(new_n630_), .B2(new_n328_), .ZN(new_n631_));
  AOI211_X1 g430(.A(KEYINPUT43), .B(new_n327_), .C1(new_n571_), .C2(new_n582_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n628_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT44), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  OAI211_X1 g434(.A(KEYINPUT44), .B(new_n628_), .C1(new_n631_), .C2(new_n632_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n580_), .A2(G29gat), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n627_), .B1(new_n637_), .B2(new_n638_), .ZN(G1328gat));
  NOR2_X1   g438(.A1(new_n521_), .A2(G36gat), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n625_), .B(new_n640_), .C1(new_n585_), .C2(new_n584_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT45), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n635_), .A2(new_n577_), .A3(new_n636_), .ZN(new_n643_));
  AND3_X1   g442(.A1(new_n643_), .A2(KEYINPUT99), .A3(G36gat), .ZN(new_n644_));
  AOI21_X1  g443(.A(KEYINPUT99), .B1(new_n643_), .B2(G36gat), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n642_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT46), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  OAI211_X1 g447(.A(KEYINPUT46), .B(new_n642_), .C1(new_n644_), .C2(new_n645_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(G1329gat));
  NAND2_X1  g449(.A1(new_n626_), .A2(new_n614_), .ZN(new_n651_));
  INV_X1    g450(.A(G43gat), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n637_), .A2(G43gat), .A3(new_n614_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(KEYINPUT100), .B(KEYINPUT47), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n653_), .A2(new_n654_), .A3(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n655_), .B1(new_n653_), .B2(new_n654_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n656_), .A2(new_n657_), .ZN(G1330gat));
  AOI21_X1  g457(.A(G50gat), .B1(new_n626_), .B2(new_n556_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n556_), .A2(G50gat), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n659_), .B1(new_n637_), .B2(new_n660_), .ZN(G1331gat));
  INV_X1    g460(.A(G57gat), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n304_), .A2(new_n347_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n278_), .A2(new_n595_), .A3(new_n663_), .ZN(new_n664_));
  XOR2_X1   g463(.A(new_n664_), .B(KEYINPUT101), .Z(new_n665_));
  AOI21_X1  g464(.A(new_n662_), .B1(new_n665_), .B2(new_n580_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n347_), .B1(new_n571_), .B2(new_n582_), .ZN(new_n667_));
  AND4_X1   g466(.A1(new_n623_), .A2(new_n667_), .A3(new_n624_), .A4(new_n327_), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n668_), .A2(new_n662_), .A3(new_n580_), .ZN(new_n669_));
  OR2_X1    g468(.A1(new_n666_), .A2(new_n669_), .ZN(G1332gat));
  NOR2_X1   g469(.A1(new_n521_), .A2(G64gat), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n671_), .B(KEYINPUT103), .Z(new_n672_));
  NAND2_X1  g471(.A1(new_n668_), .A2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n665_), .A2(new_n577_), .ZN(new_n674_));
  XOR2_X1   g473(.A(KEYINPUT102), .B(KEYINPUT48), .Z(new_n675_));
  AND3_X1   g474(.A1(new_n674_), .A2(G64gat), .A3(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n674_), .B2(G64gat), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n673_), .B1(new_n676_), .B2(new_n677_), .ZN(G1333gat));
  INV_X1    g477(.A(G71gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n668_), .A2(new_n679_), .A3(new_n614_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n665_), .A2(new_n614_), .ZN(new_n681_));
  XOR2_X1   g480(.A(KEYINPUT104), .B(KEYINPUT49), .Z(new_n682_));
  AND3_X1   g481(.A1(new_n681_), .A2(G71gat), .A3(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n682_), .B1(new_n681_), .B2(G71gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n680_), .B1(new_n683_), .B2(new_n684_), .ZN(G1334gat));
  INV_X1    g484(.A(G78gat), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n668_), .A2(new_n686_), .A3(new_n556_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT50), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n665_), .A2(new_n556_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n689_), .B2(G78gat), .ZN(new_n690_));
  AOI211_X1 g489(.A(KEYINPUT50), .B(new_n686_), .C1(new_n665_), .C2(new_n556_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n687_), .B1(new_n690_), .B2(new_n691_), .ZN(G1335gat));
  NOR3_X1   g491(.A1(new_n277_), .A2(new_n347_), .A3(new_n624_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n693_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n694_), .A2(KEYINPUT105), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n694_), .A2(KEYINPUT105), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(G85gat), .B1(new_n697_), .B2(new_n463_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n323_), .ZN(new_n699_));
  AND4_X1   g498(.A1(new_n278_), .A2(new_n304_), .A3(new_n699_), .A4(new_n667_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n700_), .A2(new_n214_), .A3(new_n580_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n698_), .A2(new_n701_), .ZN(G1336gat));
  OAI21_X1  g501(.A(G92gat), .B1(new_n697_), .B2(new_n521_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n700_), .A2(new_n215_), .A3(new_n577_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(G1337gat));
  INV_X1    g504(.A(KEYINPUT106), .ZN(new_n706_));
  OR2_X1    g505(.A1(new_n706_), .A2(KEYINPUT51), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(KEYINPUT51), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n694_), .B(KEYINPUT105), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n209_), .B1(new_n709_), .B2(new_n614_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n700_), .A2(new_n614_), .A3(new_n228_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  OAI211_X1 g511(.A(new_n707_), .B(new_n708_), .C1(new_n710_), .C2(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(G99gat), .B1(new_n697_), .B2(new_n408_), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n714_), .A2(new_n706_), .A3(KEYINPUT51), .A4(new_n711_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n713_), .A2(new_n715_), .ZN(G1338gat));
  OAI21_X1  g515(.A(G106gat), .B1(new_n694_), .B2(new_n572_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT107), .ZN(new_n718_));
  OR2_X1    g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n718_), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n719_), .A2(KEYINPUT52), .A3(new_n720_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n700_), .A2(new_n210_), .A3(new_n556_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n722_), .B1(new_n720_), .B2(KEYINPUT52), .ZN(new_n723_));
  OAI21_X1  g522(.A(KEYINPUT53), .B1(new_n721_), .B2(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n719_), .A2(KEYINPUT52), .A3(new_n720_), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n720_), .A2(KEYINPUT52), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT53), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n725_), .A2(new_n726_), .A3(new_n727_), .A4(new_n722_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n724_), .A2(new_n728_), .ZN(G1339gat));
  XOR2_X1   g528(.A(KEYINPUT115), .B(KEYINPUT59), .Z(new_n730_));
  INV_X1    g529(.A(KEYINPUT111), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n331_), .B1(new_n337_), .B2(new_n731_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n732_), .B1(new_n731_), .B2(new_n337_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n343_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  OR2_X1    g534(.A1(new_n735_), .A2(KEYINPUT112), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(KEYINPUT112), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n736_), .A2(new_n344_), .A3(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(new_n273_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT110), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n263_), .A2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT55), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n250_), .A2(new_n259_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(new_n261_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT55), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n263_), .A2(new_n740_), .A3(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n742_), .A2(new_n744_), .A3(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(new_n271_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT56), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n747_), .A2(KEYINPUT56), .A3(new_n271_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n739_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n328_), .B1(new_n752_), .B2(KEYINPUT58), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(KEYINPUT113), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n752_), .A2(KEYINPUT58), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT113), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n756_), .B(new_n328_), .C1(new_n752_), .C2(KEYINPUT58), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n754_), .A2(new_n755_), .A3(new_n757_), .ZN(new_n758_));
  AND3_X1   g557(.A1(new_n347_), .A2(KEYINPUT109), .A3(new_n273_), .ZN(new_n759_));
  AOI21_X1  g558(.A(KEYINPUT109), .B1(new_n347_), .B2(new_n273_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n747_), .A2(KEYINPUT56), .A3(new_n271_), .ZN(new_n762_));
  AOI21_X1  g561(.A(KEYINPUT56), .B1(new_n747_), .B2(new_n271_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n761_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n738_), .A2(new_n274_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(KEYINPUT57), .B1(new_n766_), .B2(new_n323_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT57), .ZN(new_n768_));
  AOI211_X1 g567(.A(new_n768_), .B(new_n699_), .C1(new_n764_), .C2(new_n765_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n767_), .A2(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n624_), .B1(new_n758_), .B2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT54), .ZN(new_n772_));
  XOR2_X1   g571(.A(new_n663_), .B(KEYINPUT108), .Z(new_n773_));
  NOR2_X1   g572(.A1(new_n773_), .A2(new_n328_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n772_), .B1(new_n774_), .B2(new_n277_), .ZN(new_n775_));
  NOR4_X1   g574(.A1(new_n773_), .A2(new_n623_), .A3(new_n328_), .A4(KEYINPUT54), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n771_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n579_), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n779_), .A2(new_n463_), .A3(new_n408_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n730_), .B1(new_n778_), .B2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT59), .ZN(new_n783_));
  OAI221_X1 g582(.A(new_n780_), .B1(KEYINPUT115), .B2(new_n783_), .C1(new_n771_), .C2(new_n777_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n782_), .A2(G113gat), .A3(new_n347_), .A4(new_n784_), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n347_), .B(new_n780_), .C1(new_n771_), .C2(new_n777_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT114), .ZN(new_n787_));
  INV_X1    g586(.A(G113gat), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n786_), .A2(new_n787_), .A3(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n786_), .A2(new_n788_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT114), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n785_), .A2(new_n789_), .A3(new_n791_), .ZN(G1340gat));
  NAND3_X1  g591(.A1(new_n782_), .A2(new_n278_), .A3(new_n784_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(G120gat), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n758_), .A2(new_n770_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n304_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n777_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT60), .ZN(new_n799_));
  AOI21_X1  g598(.A(G120gat), .B1(new_n623_), .B2(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n800_), .B1(new_n799_), .B2(G120gat), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n798_), .A2(new_n780_), .A3(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n794_), .A2(new_n802_), .ZN(G1341gat));
  AND2_X1   g602(.A1(new_n782_), .A2(new_n784_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n304_), .A2(KEYINPUT116), .ZN(new_n805_));
  MUX2_X1   g604(.A(KEYINPUT116), .B(new_n805_), .S(G127gat), .Z(new_n806_));
  INV_X1    g605(.A(G127gat), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n798_), .A2(new_n624_), .A3(new_n780_), .ZN(new_n808_));
  AOI22_X1  g607(.A1(new_n804_), .A2(new_n806_), .B1(new_n807_), .B2(new_n808_), .ZN(G1342gat));
  NAND4_X1  g608(.A1(new_n782_), .A2(G134gat), .A3(new_n328_), .A4(new_n784_), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n594_), .B(new_n780_), .C1(new_n771_), .C2(new_n777_), .ZN(new_n811_));
  INV_X1    g610(.A(G134gat), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n811_), .A2(KEYINPUT117), .A3(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n811_), .A2(new_n812_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT117), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  AND3_X1   g615(.A1(new_n810_), .A2(new_n813_), .A3(new_n816_), .ZN(G1343gat));
  NOR2_X1   g616(.A1(new_n614_), .A2(new_n572_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n818_), .A2(new_n580_), .A3(new_n521_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n778_), .A2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n347_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(KEYINPUT118), .B(G141gat), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n821_), .B(new_n822_), .ZN(G1344gat));
  NAND2_X1  g622(.A1(new_n820_), .A2(new_n278_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(KEYINPUT119), .B(G148gat), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n824_), .B(new_n825_), .ZN(G1345gat));
  NAND2_X1  g625(.A1(new_n820_), .A2(new_n624_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(KEYINPUT61), .B(G155gat), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n827_), .B(new_n828_), .ZN(G1346gat));
  INV_X1    g628(.A(new_n819_), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n594_), .B(new_n830_), .C1(new_n771_), .C2(new_n777_), .ZN(new_n831_));
  INV_X1    g630(.A(G162gat), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(KEYINPUT120), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT120), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n831_), .A2(new_n835_), .A3(new_n832_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n327_), .A2(new_n832_), .ZN(new_n837_));
  AOI22_X1  g636(.A1(new_n834_), .A2(new_n836_), .B1(new_n820_), .B2(new_n837_), .ZN(G1347gat));
  NAND3_X1  g637(.A1(new_n581_), .A2(new_n572_), .A3(new_n577_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n798_), .A2(new_n347_), .A3(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(G169gat), .ZN(new_n842_));
  XNOR2_X1  g641(.A(KEYINPUT121), .B(KEYINPUT62), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n843_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n841_), .A2(G169gat), .A3(new_n845_), .ZN(new_n846_));
  OR2_X1    g645(.A1(new_n841_), .A2(new_n471_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n844_), .A2(new_n846_), .A3(new_n847_), .ZN(G1348gat));
  AOI21_X1  g647(.A(new_n839_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n366_), .B1(new_n849_), .B2(new_n623_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n278_), .A2(G176gat), .ZN(new_n851_));
  NOR3_X1   g650(.A1(new_n778_), .A2(new_n839_), .A3(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(KEYINPUT122), .B1(new_n850_), .B2(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n849_), .A2(G176gat), .A3(new_n278_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT122), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n778_), .A2(new_n277_), .A3(new_n839_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n854_), .B(new_n855_), .C1(new_n856_), .C2(new_n366_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n853_), .A2(new_n857_), .ZN(G1349gat));
  INV_X1    g657(.A(new_n382_), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n798_), .A2(new_n859_), .A3(new_n624_), .A4(new_n840_), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n624_), .B(new_n840_), .C1(new_n771_), .C2(new_n777_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n356_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT123), .ZN(new_n863_));
  AND3_X1   g662(.A1(new_n860_), .A2(new_n862_), .A3(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n863_), .B1(new_n860_), .B2(new_n862_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n864_), .A2(new_n865_), .ZN(G1350gat));
  INV_X1    g665(.A(KEYINPUT124), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n357_), .B1(new_n849_), .B2(new_n328_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n594_), .A2(new_n484_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n778_), .A2(new_n839_), .A3(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n867_), .B1(new_n868_), .B2(new_n870_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n849_), .A2(new_n484_), .A3(new_n594_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n778_), .A2(new_n327_), .A3(new_n839_), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n872_), .B(KEYINPUT124), .C1(new_n873_), .C2(new_n357_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n871_), .A2(new_n874_), .ZN(G1351gat));
  AND3_X1   g674(.A1(new_n818_), .A2(KEYINPUT125), .A3(new_n463_), .ZN(new_n876_));
  AOI21_X1  g675(.A(KEYINPUT125), .B1(new_n818_), .B2(new_n463_), .ZN(new_n877_));
  OR3_X1    g676(.A1(new_n876_), .A2(new_n877_), .A3(new_n521_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n778_), .A2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(KEYINPUT126), .A2(G197gat), .ZN(new_n880_));
  OR2_X1    g679(.A1(KEYINPUT126), .A2(G197gat), .ZN(new_n881_));
  AOI22_X1  g680(.A1(new_n879_), .A2(new_n347_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n778_), .A2(new_n348_), .A3(new_n878_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n882_), .B1(new_n883_), .B2(new_n881_), .ZN(G1352gat));
  NAND2_X1  g683(.A1(new_n879_), .A2(new_n278_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n885_), .B1(KEYINPUT127), .B2(G204gat), .ZN(new_n886_));
  XNOR2_X1  g685(.A(KEYINPUT127), .B(G204gat), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n879_), .A2(new_n278_), .A3(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n888_), .ZN(G1353gat));
  NOR3_X1   g688(.A1(new_n778_), .A2(new_n304_), .A3(new_n878_), .ZN(new_n890_));
  OR2_X1    g689(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  XOR2_X1   g691(.A(KEYINPUT63), .B(G211gat), .Z(new_n893_));
  AOI21_X1  g692(.A(new_n892_), .B1(new_n890_), .B2(new_n893_), .ZN(G1354gat));
  INV_X1    g693(.A(G218gat), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n879_), .A2(new_n895_), .A3(new_n594_), .ZN(new_n896_));
  NOR3_X1   g695(.A1(new_n778_), .A2(new_n327_), .A3(new_n878_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n895_), .B2(new_n897_), .ZN(G1355gat));
endmodule


