//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 1 0 0 0 0 1 1 0 1 0 0 1 0 1 0 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 1 1 1 1 1 1 0 1 1 0 0 1 1 0 1 1 0 1 0 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n587_,
    new_n588_, new_n589_, new_n591_, new_n592_, new_n593_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n669_, new_n670_, new_n671_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n829_, new_n831_, new_n832_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n852_, new_n853_, new_n854_, new_n856_, new_n857_, new_n859_,
    new_n860_, new_n861_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n874_,
    new_n875_, new_n876_, new_n877_;
  NAND2_X1  g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(new_n202_), .B(KEYINPUT94), .Z(new_n203_));
  INV_X1    g002(.A(G155gat), .ZN(new_n204_));
  INV_X1    g003(.A(G162gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT93), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n208_), .A2(KEYINPUT2), .ZN(new_n209_));
  OR3_X1    g008(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT2), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n210_), .B(new_n211_), .C1(new_n212_), .C2(new_n207_), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n203_), .B(new_n206_), .C1(new_n209_), .C2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT95), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n214_), .B(new_n215_), .ZN(new_n216_));
  AOI22_X1  g015(.A1(new_n203_), .A2(KEYINPUT1), .B1(new_n204_), .B2(new_n205_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n217_), .B1(KEYINPUT1), .B2(new_n203_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n208_), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n218_), .B(new_n219_), .C1(G141gat), .C2(G148gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n216_), .A2(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(G127gat), .B(G134gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G113gat), .B(G120gat), .ZN(new_n223_));
  XOR2_X1   g022(.A(new_n222_), .B(new_n223_), .Z(new_n224_));
  OR2_X1    g023(.A1(new_n221_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n221_), .A2(new_n224_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(KEYINPUT4), .A3(new_n226_), .ZN(new_n227_));
  OR2_X1    g026(.A1(new_n226_), .A2(KEYINPUT4), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G225gat), .A2(G233gat), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G1gat), .B(G29gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(G85gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT0), .B(G57gat), .ZN(new_n235_));
  XOR2_X1   g034(.A(new_n234_), .B(new_n235_), .Z(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n225_), .A2(new_n226_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(new_n230_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n232_), .A2(new_n237_), .A3(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n239_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n230_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n236_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n240_), .A2(new_n243_), .A3(KEYINPUT105), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT105), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n232_), .A2(new_n245_), .A3(new_n237_), .A4(new_n239_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT20), .ZN(new_n247_));
  INV_X1    g046(.A(G204gat), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n248_), .A2(G197gat), .ZN(new_n249_));
  INV_X1    g048(.A(G197gat), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n250_), .A2(G204gat), .ZN(new_n251_));
  OAI21_X1  g050(.A(KEYINPUT21), .B1(new_n249_), .B2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G211gat), .B(G218gat), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT99), .B1(new_n248_), .B2(G197gat), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT99), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n255_), .A2(new_n250_), .A3(G204gat), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n254_), .B(new_n256_), .C1(new_n250_), .C2(G204gat), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n252_), .B(new_n253_), .C1(new_n257_), .C2(KEYINPUT21), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT100), .ZN(new_n259_));
  INV_X1    g058(.A(new_n253_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n257_), .A2(KEYINPUT21), .A3(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G183gat), .A2(G190gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT23), .ZN(new_n264_));
  OR2_X1    g063(.A1(G169gat), .A2(G176gat), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n264_), .B1(KEYINPUT24), .B2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT25), .B(G183gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT26), .B(G190gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G169gat), .A2(G176gat), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n265_), .A2(KEYINPUT24), .A3(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n266_), .B1(KEYINPUT104), .B2(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n273_), .B1(KEYINPUT104), .B2(new_n272_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n264_), .B1(G183gat), .B2(G190gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT22), .B(G169gat), .ZN(new_n276_));
  INV_X1    g075(.A(G176gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n275_), .A2(new_n270_), .A3(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n274_), .A2(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n247_), .B1(new_n262_), .B2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n278_), .B(KEYINPUT87), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n282_), .A2(new_n270_), .A3(new_n275_), .ZN(new_n283_));
  OAI211_X1 g082(.A(new_n269_), .B(new_n264_), .C1(KEYINPUT24), .C2(new_n265_), .ZN(new_n284_));
  XOR2_X1   g083(.A(new_n271_), .B(KEYINPUT86), .Z(new_n285_));
  OAI21_X1  g084(.A(new_n283_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n281_), .B1(new_n262_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G226gat), .A2(G233gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT19), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n287_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n289_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n262_), .A2(new_n280_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n292_), .A2(new_n247_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n262_), .A2(new_n286_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n291_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n290_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n287_), .A2(new_n289_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n293_), .A2(new_n291_), .A3(new_n294_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G8gat), .B(G36gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT18), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G64gat), .B(G92gat), .ZN(new_n302_));
  XOR2_X1   g101(.A(new_n301_), .B(new_n302_), .Z(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT32), .ZN(new_n304_));
  MUX2_X1   g103(.A(new_n296_), .B(new_n299_), .S(new_n304_), .Z(new_n305_));
  NAND3_X1  g104(.A1(new_n244_), .A2(new_n246_), .A3(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT33), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n243_), .A2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n299_), .B(new_n303_), .ZN(new_n309_));
  OAI211_X1 g108(.A(KEYINPUT33), .B(new_n236_), .C1(new_n241_), .C2(new_n242_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n227_), .A2(new_n230_), .A3(new_n228_), .ZN(new_n311_));
  OAI211_X1 g110(.A(new_n311_), .B(new_n237_), .C1(new_n230_), .C2(new_n238_), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n308_), .A2(new_n309_), .A3(new_n310_), .A4(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n306_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G228gat), .A2(G233gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n262_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n221_), .A2(KEYINPUT29), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT98), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n221_), .A2(KEYINPUT98), .A3(KEYINPUT29), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n316_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT101), .B(KEYINPUT29), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n221_), .A2(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n315_), .B1(new_n323_), .B2(new_n262_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G78gat), .B(G106gat), .ZN(new_n325_));
  NOR3_X1   g124(.A1(new_n321_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  OR2_X1    g125(.A1(new_n326_), .A2(KEYINPUT102), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(KEYINPUT102), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n325_), .B1(new_n321_), .B2(new_n324_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n327_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  XOR2_X1   g129(.A(KEYINPUT96), .B(KEYINPUT28), .Z(new_n331_));
  OAI21_X1  g130(.A(new_n331_), .B1(new_n221_), .B2(KEYINPUT29), .ZN(new_n332_));
  XOR2_X1   g131(.A(G22gat), .B(G50gat), .Z(new_n333_));
  INV_X1    g132(.A(KEYINPUT29), .ZN(new_n334_));
  INV_X1    g133(.A(new_n331_), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n216_), .A2(new_n334_), .A3(new_n220_), .A4(new_n335_), .ZN(new_n336_));
  AND3_X1   g135(.A1(new_n332_), .A2(new_n333_), .A3(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n333_), .B1(new_n332_), .B2(new_n336_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT97), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n329_), .A2(new_n339_), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT103), .B1(new_n341_), .B2(new_n326_), .ZN(new_n342_));
  OR3_X1    g141(.A1(new_n321_), .A2(new_n325_), .A3(new_n324_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT103), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n343_), .A2(new_n339_), .A3(new_n344_), .A4(new_n329_), .ZN(new_n345_));
  AOI22_X1  g144(.A1(new_n330_), .A2(new_n340_), .B1(new_n342_), .B2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n314_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n342_), .A2(new_n345_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n328_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n329_), .B1(new_n326_), .B2(KEYINPUT102), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n340_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n348_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n244_), .A2(new_n246_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n309_), .A2(KEYINPUT27), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n296_), .A2(new_n303_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n303_), .ZN(new_n356_));
  OAI21_X1  g155(.A(KEYINPUT27), .B1(new_n299_), .B2(new_n356_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n354_), .A2(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n352_), .A2(new_n353_), .A3(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n347_), .A2(new_n360_), .ZN(new_n361_));
  XOR2_X1   g160(.A(new_n286_), .B(KEYINPUT30), .Z(new_n362_));
  OR2_X1    g161(.A1(new_n362_), .A2(KEYINPUT90), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(KEYINPUT90), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G227gat), .A2(G233gat), .ZN(new_n365_));
  XOR2_X1   g164(.A(new_n365_), .B(G15gat), .Z(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(G71gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(G99gat), .ZN(new_n368_));
  XOR2_X1   g167(.A(KEYINPUT88), .B(G43gat), .Z(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT89), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n368_), .B(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n363_), .A2(new_n364_), .A3(new_n371_), .ZN(new_n372_));
  OR2_X1    g171(.A1(new_n364_), .A2(new_n371_), .ZN(new_n373_));
  XOR2_X1   g172(.A(new_n224_), .B(KEYINPUT31), .Z(new_n374_));
  XOR2_X1   g173(.A(new_n374_), .B(KEYINPUT91), .Z(new_n375_));
  NAND3_X1  g174(.A1(new_n372_), .A2(new_n373_), .A3(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT92), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n374_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n376_), .A2(new_n377_), .ZN(new_n381_));
  OR2_X1    g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n359_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n383_), .A2(new_n352_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n353_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n382_), .A2(new_n385_), .ZN(new_n386_));
  AOI22_X1  g185(.A1(new_n361_), .A2(new_n382_), .B1(new_n384_), .B2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G230gat), .A2(G233gat), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  XOR2_X1   g188(.A(KEYINPUT10), .B(G99gat), .Z(new_n390_));
  INV_X1    g189(.A(G106gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  XOR2_X1   g191(.A(G85gat), .B(G92gat), .Z(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(KEYINPUT9), .ZN(new_n394_));
  INV_X1    g193(.A(G85gat), .ZN(new_n395_));
  INV_X1    g194(.A(G92gat), .ZN(new_n396_));
  OR3_X1    g195(.A1(new_n395_), .A2(new_n396_), .A3(KEYINPUT9), .ZN(new_n397_));
  AND3_X1   g196(.A1(new_n392_), .A2(new_n394_), .A3(new_n397_), .ZN(new_n398_));
  AND2_X1   g197(.A1(G99gat), .A2(G106gat), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT64), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n401_), .A2(KEYINPUT6), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT6), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n403_), .A2(KEYINPUT64), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n400_), .B1(new_n402_), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(KEYINPUT64), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n401_), .A2(KEYINPUT6), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n406_), .A2(new_n407_), .A3(new_n399_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n405_), .A2(KEYINPUT65), .A3(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT65), .ZN(new_n410_));
  AND3_X1   g209(.A1(new_n406_), .A2(new_n407_), .A3(new_n399_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n399_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n410_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n398_), .A2(new_n409_), .A3(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(G99gat), .A2(G106gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT7), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n413_), .A2(new_n409_), .A3(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT66), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT66), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n413_), .A2(new_n409_), .A3(new_n420_), .A4(new_n417_), .ZN(new_n421_));
  XOR2_X1   g220(.A(KEYINPUT67), .B(KEYINPUT8), .Z(new_n422_));
  AND2_X1   g221(.A1(new_n422_), .A2(new_n393_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n419_), .A2(new_n421_), .A3(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT68), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n425_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n405_), .A2(KEYINPUT68), .A3(new_n408_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n426_), .A2(new_n427_), .A3(new_n417_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(new_n393_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT8), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n415_), .B1(new_n424_), .B2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G57gat), .B(G64gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(KEYINPUT11), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G71gat), .B(G78gat), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n433_), .A2(new_n435_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n432_), .A2(KEYINPUT11), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n437_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n389_), .B1(new_n431_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(KEYINPUT70), .A2(KEYINPUT12), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n424_), .A2(new_n430_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(new_n414_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n440_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n442_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n442_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(KEYINPUT70), .A2(KEYINPUT12), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NOR3_X1   g249(.A1(new_n431_), .A2(new_n440_), .A3(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n441_), .B1(new_n446_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT71), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n431_), .A2(new_n440_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT69), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n444_), .A2(new_n445_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n431_), .A2(KEYINPUT69), .A3(new_n440_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n456_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(new_n389_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT71), .ZN(new_n461_));
  OAI211_X1 g260(.A(new_n461_), .B(new_n441_), .C1(new_n446_), .C2(new_n451_), .ZN(new_n462_));
  XOR2_X1   g261(.A(G120gat), .B(G148gat), .Z(new_n463_));
  XNOR2_X1  g262(.A(G176gat), .B(G204gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n465_), .B(new_n466_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n453_), .A2(new_n460_), .A3(new_n462_), .A4(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT73), .ZN(new_n469_));
  AND2_X1   g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n468_), .A2(new_n469_), .ZN(new_n471_));
  AND3_X1   g270(.A1(new_n453_), .A2(new_n460_), .A3(new_n462_), .ZN(new_n472_));
  OAI22_X1  g271(.A1(new_n470_), .A2(new_n471_), .B1(new_n472_), .B2(new_n467_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT13), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n473_), .A2(new_n474_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(KEYINPUT79), .B(G15gat), .ZN(new_n478_));
  INV_X1    g277(.A(G22gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(G1gat), .ZN(new_n481_));
  INV_X1    g280(.A(G8gat), .ZN(new_n482_));
  OAI21_X1  g281(.A(KEYINPUT14), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n480_), .A2(new_n483_), .ZN(new_n484_));
  XOR2_X1   g283(.A(G1gat), .B(G8gat), .Z(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G29gat), .B(G36gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G43gat), .B(G50gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT82), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n486_), .B(new_n490_), .Z(new_n491_));
  NAND3_X1  g290(.A1(new_n491_), .A2(G229gat), .A3(G233gat), .ZN(new_n492_));
  INV_X1    g291(.A(new_n486_), .ZN(new_n493_));
  OR2_X1    g292(.A1(new_n493_), .A2(new_n490_), .ZN(new_n494_));
  XOR2_X1   g293(.A(KEYINPUT74), .B(KEYINPUT15), .Z(new_n495_));
  XNOR2_X1  g294(.A(new_n489_), .B(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n493_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G229gat), .A2(G233gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT83), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n494_), .A2(new_n497_), .A3(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n492_), .A2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G113gat), .B(G141gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT85), .ZN(new_n503_));
  XOR2_X1   g302(.A(G169gat), .B(G197gat), .Z(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n506_), .A2(KEYINPUT84), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n501_), .B(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n477_), .A2(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n387_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G190gat), .B(G218gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G134gat), .B(G162gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  XOR2_X1   g312(.A(new_n513_), .B(KEYINPUT36), .Z(new_n514_));
  INV_X1    g313(.A(KEYINPUT35), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G232gat), .A2(G233gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT34), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  AOI22_X1  g317(.A1(new_n444_), .A2(new_n496_), .B1(new_n515_), .B2(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n518_), .A2(new_n515_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT75), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n431_), .A2(new_n522_), .A3(new_n489_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n522_), .B1(new_n431_), .B2(new_n489_), .ZN(new_n525_));
  OAI211_X1 g324(.A(new_n519_), .B(new_n521_), .C1(new_n524_), .C2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n443_), .A2(new_n414_), .A3(new_n489_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT75), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(new_n523_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n521_), .B1(new_n530_), .B2(new_n519_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n514_), .B1(new_n527_), .B2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(KEYINPUT77), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n519_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(new_n520_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(new_n526_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT77), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n536_), .A2(new_n537_), .A3(new_n514_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n513_), .A2(KEYINPUT36), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n535_), .A2(new_n539_), .A3(new_n526_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT76), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n535_), .A2(KEYINPUT76), .A3(new_n539_), .A4(new_n526_), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n533_), .A2(new_n538_), .A3(new_n542_), .A4(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(KEYINPUT37), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT78), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n536_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n535_), .A2(KEYINPUT78), .A3(new_n526_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n547_), .A2(new_n548_), .A3(new_n514_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT37), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n549_), .A2(new_n550_), .A3(new_n540_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n545_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  XOR2_X1   g352(.A(G127gat), .B(G155gat), .Z(new_n554_));
  XNOR2_X1  g353(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  XOR2_X1   g355(.A(G183gat), .B(G211gat), .Z(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G231gat), .A2(G233gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n486_), .B(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(new_n440_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n558_), .B1(new_n561_), .B2(KEYINPUT81), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n558_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n562_), .B1(KEYINPUT17), .B2(new_n563_), .ZN(new_n564_));
  AND2_X1   g363(.A1(new_n562_), .A2(KEYINPUT17), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n553_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n510_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n570_), .A2(new_n481_), .A3(new_n385_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT38), .ZN(new_n572_));
  OR2_X1    g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n549_), .A2(new_n540_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NOR4_X1   g374(.A1(new_n387_), .A2(new_n509_), .A3(new_n567_), .A4(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  OAI21_X1  g376(.A(G1gat), .B1(new_n577_), .B2(new_n353_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n571_), .A2(new_n572_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n573_), .A2(new_n578_), .A3(new_n579_), .ZN(G1324gat));
  AOI21_X1  g379(.A(new_n482_), .B1(new_n576_), .B2(new_n383_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT39), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n570_), .A2(new_n482_), .A3(new_n383_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  XOR2_X1   g384(.A(new_n585_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g385(.A(G15gat), .B1(new_n577_), .B2(new_n382_), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n587_), .B(KEYINPUT41), .Z(new_n588_));
  OR2_X1    g387(.A1(new_n382_), .A2(G15gat), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n588_), .B1(new_n569_), .B2(new_n589_), .ZN(G1326gat));
  AOI21_X1  g389(.A(new_n479_), .B1(new_n576_), .B2(new_n352_), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n591_), .B(KEYINPUT42), .Z(new_n592_));
  NAND3_X1  g391(.A1(new_n570_), .A2(new_n479_), .A3(new_n352_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(G1327gat));
  NOR2_X1   g393(.A1(new_n566_), .A2(new_n574_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NOR3_X1   g395(.A1(new_n387_), .A2(new_n509_), .A3(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(G29gat), .B1(new_n597_), .B2(new_n385_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT43), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n599_), .B1(new_n553_), .B2(KEYINPUT106), .ZN(new_n600_));
  OR3_X1    g399(.A1(new_n387_), .A2(new_n552_), .A3(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n600_), .B1(new_n387_), .B2(new_n552_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n509_), .A2(new_n566_), .ZN(new_n604_));
  AOI21_X1  g403(.A(KEYINPUT44), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT44), .ZN(new_n606_));
  INV_X1    g405(.A(new_n604_), .ZN(new_n607_));
  AOI211_X1 g406(.A(new_n606_), .B(new_n607_), .C1(new_n601_), .C2(new_n602_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n605_), .A2(new_n608_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n385_), .A2(G29gat), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n598_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT107), .ZN(G1328gat));
  INV_X1    g411(.A(KEYINPUT108), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n359_), .A2(G36gat), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n613_), .B1(new_n597_), .B2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n597_), .A2(new_n613_), .A3(new_n614_), .ZN(new_n617_));
  AND3_X1   g416(.A1(new_n616_), .A2(KEYINPUT45), .A3(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(KEYINPUT45), .B1(new_n616_), .B2(new_n617_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NOR3_X1   g419(.A1(new_n605_), .A2(new_n608_), .A3(new_n359_), .ZN(new_n621_));
  INV_X1    g420(.A(G36gat), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n620_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT46), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  OAI211_X1 g424(.A(new_n620_), .B(KEYINPUT46), .C1(new_n621_), .C2(new_n622_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(G1329gat));
  INV_X1    g426(.A(new_n382_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(G43gat), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n605_), .A2(new_n608_), .A3(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(G43gat), .B1(new_n597_), .B2(new_n628_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT109), .Z(new_n632_));
  OR3_X1    g431(.A1(new_n630_), .A2(new_n632_), .A3(KEYINPUT47), .ZN(new_n633_));
  OAI21_X1  g432(.A(KEYINPUT47), .B1(new_n630_), .B2(new_n632_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(G1330gat));
  INV_X1    g434(.A(KEYINPUT110), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n603_), .A2(new_n604_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(new_n606_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n603_), .A2(KEYINPUT44), .A3(new_n604_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n638_), .A2(new_n352_), .A3(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(G50gat), .ZN(new_n641_));
  INV_X1    g440(.A(new_n597_), .ZN(new_n642_));
  NOR3_X1   g441(.A1(new_n642_), .A2(G50gat), .A3(new_n346_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n636_), .B1(new_n641_), .B2(new_n644_), .ZN(new_n645_));
  AOI211_X1 g444(.A(KEYINPUT110), .B(new_n643_), .C1(new_n640_), .C2(G50gat), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n645_), .A2(new_n646_), .ZN(G1331gat));
  NOR2_X1   g446(.A1(new_n387_), .A2(new_n575_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n477_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n508_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n566_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n648_), .A2(new_n649_), .A3(new_n652_), .ZN(new_n653_));
  OR2_X1    g452(.A1(new_n653_), .A2(KEYINPUT111), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(KEYINPUT111), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(G57gat), .B1(new_n656_), .B2(new_n353_), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n387_), .A2(new_n508_), .A3(new_n477_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(new_n568_), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n353_), .A2(G57gat), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n657_), .B1(new_n659_), .B2(new_n660_), .ZN(G1332gat));
  OR3_X1    g460(.A1(new_n659_), .A2(G64gat), .A3(new_n359_), .ZN(new_n662_));
  OAI21_X1  g461(.A(G64gat), .B1(new_n656_), .B2(new_n359_), .ZN(new_n663_));
  XOR2_X1   g462(.A(KEYINPUT112), .B(KEYINPUT48), .Z(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n663_), .A2(new_n665_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n663_), .A2(new_n665_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n662_), .B1(new_n666_), .B2(new_n667_), .ZN(G1333gat));
  OAI21_X1  g467(.A(G71gat), .B1(new_n656_), .B2(new_n382_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT49), .ZN(new_n670_));
  OR3_X1    g469(.A1(new_n659_), .A2(G71gat), .A3(new_n382_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(G1334gat));
  OR3_X1    g471(.A1(new_n659_), .A2(G78gat), .A3(new_n346_), .ZN(new_n673_));
  OAI21_X1  g472(.A(G78gat), .B1(new_n656_), .B2(new_n346_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n674_), .A2(KEYINPUT50), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n674_), .A2(KEYINPUT50), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n673_), .B1(new_n675_), .B2(new_n676_), .ZN(G1335gat));
  NOR3_X1   g476(.A1(new_n477_), .A2(new_n566_), .A3(new_n508_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT113), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n603_), .A2(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n601_), .A2(KEYINPUT113), .A3(new_n602_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n679_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(G85gat), .B1(new_n684_), .B2(new_n353_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n658_), .A2(new_n595_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n687_), .A2(new_n395_), .A3(new_n385_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n685_), .A2(new_n688_), .ZN(G1336gat));
  OAI21_X1  g488(.A(G92gat), .B1(new_n684_), .B2(new_n359_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n687_), .A2(new_n396_), .A3(new_n383_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1337gat));
  INV_X1    g491(.A(G99gat), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n693_), .B1(new_n683_), .B2(new_n628_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n687_), .A2(new_n390_), .A3(new_n628_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n695_), .A2(new_n696_), .A3(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n697_), .ZN(new_n699_));
  OAI211_X1 g498(.A(KEYINPUT114), .B(KEYINPUT51), .C1(new_n694_), .C2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n698_), .A2(new_n700_), .ZN(G1338gat));
  NAND2_X1  g500(.A1(new_n678_), .A2(new_n352_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n391_), .B1(new_n603_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT52), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n704_), .B(new_n705_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n687_), .A2(new_n391_), .A3(new_n352_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(KEYINPUT53), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT53), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n706_), .A2(new_n710_), .A3(new_n707_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n709_), .A2(new_n711_), .ZN(G1339gat));
  NOR2_X1   g511(.A1(new_n553_), .A2(new_n651_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT54), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n713_), .A2(new_n714_), .A3(new_n477_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n713_), .B2(new_n477_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n505_), .B1(new_n492_), .B2(new_n500_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n491_), .A2(new_n499_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n499_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n494_), .A2(new_n497_), .A3(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n506_), .B1(new_n719_), .B2(new_n721_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n718_), .A2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n473_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT115), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n726_), .B(new_n508_), .C1(new_n470_), .C2(new_n471_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT56), .ZN(new_n728_));
  INV_X1    g527(.A(new_n441_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n457_), .A2(new_n447_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n451_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n729_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  OAI211_X1 g531(.A(new_n456_), .B(new_n458_), .C1(new_n446_), .C2(new_n451_), .ZN(new_n733_));
  AOI22_X1  g532(.A1(new_n732_), .A2(KEYINPUT55), .B1(new_n733_), .B2(new_n389_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT55), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n453_), .A2(new_n735_), .A3(new_n462_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n467_), .B1(new_n734_), .B2(new_n736_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n728_), .B1(new_n737_), .B2(KEYINPUT116), .ZN(new_n738_));
  INV_X1    g537(.A(new_n467_), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n453_), .A2(new_n735_), .A3(new_n462_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n732_), .A2(KEYINPUT55), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n733_), .A2(new_n389_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n739_), .B1(new_n740_), .B2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT116), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n744_), .A2(new_n745_), .A3(KEYINPUT56), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n727_), .A2(new_n738_), .A3(new_n746_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n468_), .B(new_n469_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n726_), .B1(new_n748_), .B2(new_n508_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n725_), .B1(new_n747_), .B2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT57), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n575_), .A2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n748_), .A2(new_n724_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT58), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(KEYINPUT117), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n737_), .A2(new_n728_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n744_), .A2(KEYINPUT56), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n754_), .A2(new_n756_), .A3(new_n757_), .A4(new_n758_), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n758_), .A2(new_n748_), .A3(new_n724_), .A4(new_n757_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n756_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n759_), .A2(new_n762_), .A3(new_n553_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n508_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(KEYINPUT115), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n765_), .A2(new_n727_), .A3(new_n738_), .A4(new_n746_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n575_), .B1(new_n766_), .B2(new_n725_), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n753_), .B(new_n763_), .C1(new_n767_), .C2(KEYINPUT57), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n566_), .B1(new_n768_), .B2(KEYINPUT118), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n552_), .B1(new_n761_), .B2(new_n760_), .ZN(new_n770_));
  AOI22_X1  g569(.A1(new_n759_), .A2(new_n770_), .B1(new_n750_), .B2(new_n752_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n750_), .A2(new_n574_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(new_n751_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT118), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n771_), .A2(new_n773_), .A3(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n717_), .B1(new_n769_), .B2(new_n775_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n382_), .A2(new_n353_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(new_n384_), .ZN(new_n778_));
  OAI21_X1  g577(.A(KEYINPUT59), .B1(new_n776_), .B2(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n566_), .B1(new_n771_), .B2(new_n773_), .ZN(new_n780_));
  OR2_X1    g579(.A1(new_n780_), .A2(new_n717_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT59), .ZN(new_n782_));
  INV_X1    g581(.A(new_n778_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n781_), .A2(new_n782_), .A3(new_n783_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n779_), .A2(G113gat), .A3(new_n508_), .A4(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(KEYINPUT119), .B1(new_n776_), .B2(new_n778_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n753_), .A2(new_n763_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT57), .B1(new_n750_), .B2(new_n574_), .ZN(new_n789_));
  OAI21_X1  g588(.A(KEYINPUT118), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n790_), .A2(new_n775_), .A3(new_n567_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n717_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT119), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n793_), .A2(new_n794_), .A3(new_n783_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n787_), .A2(new_n795_), .A3(new_n508_), .ZN(new_n796_));
  INV_X1    g595(.A(G113gat), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT120), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n796_), .A2(KEYINPUT120), .A3(new_n797_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n786_), .B1(new_n800_), .B2(new_n801_), .ZN(G1340gat));
  INV_X1    g601(.A(KEYINPUT60), .ZN(new_n803_));
  AOI21_X1  g602(.A(G120gat), .B1(new_n649_), .B2(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(new_n803_), .B2(G120gat), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n787_), .A2(new_n795_), .A3(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n779_), .A2(new_n649_), .A3(new_n784_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT121), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(G120gat), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n807_), .A2(new_n808_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n806_), .B1(new_n810_), .B2(new_n811_), .ZN(G1341gat));
  AND2_X1   g611(.A1(new_n779_), .A2(new_n784_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n567_), .A2(KEYINPUT122), .ZN(new_n814_));
  MUX2_X1   g613(.A(KEYINPUT122), .B(new_n814_), .S(G127gat), .Z(new_n815_));
  NAND3_X1  g614(.A1(new_n787_), .A2(new_n795_), .A3(new_n566_), .ZN(new_n816_));
  INV_X1    g615(.A(G127gat), .ZN(new_n817_));
  AOI22_X1  g616(.A1(new_n813_), .A2(new_n815_), .B1(new_n816_), .B2(new_n817_), .ZN(G1342gat));
  NAND2_X1  g617(.A1(new_n553_), .A2(G134gat), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n819_), .B(KEYINPUT123), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n787_), .A2(new_n795_), .A3(new_n575_), .ZN(new_n821_));
  INV_X1    g620(.A(G134gat), .ZN(new_n822_));
  AOI22_X1  g621(.A1(new_n813_), .A2(new_n820_), .B1(new_n821_), .B2(new_n822_), .ZN(G1343gat));
  NOR4_X1   g622(.A1(new_n628_), .A2(new_n353_), .A3(new_n346_), .A4(new_n383_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n793_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n508_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n649_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n829_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g629(.A1(new_n825_), .A2(new_n567_), .ZN(new_n831_));
  XOR2_X1   g630(.A(KEYINPUT61), .B(G155gat), .Z(new_n832_));
  XNOR2_X1  g631(.A(new_n831_), .B(new_n832_), .ZN(G1346gat));
  OAI21_X1  g632(.A(G162gat), .B1(new_n825_), .B2(new_n552_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n575_), .A2(new_n205_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n834_), .B1(new_n825_), .B2(new_n835_), .ZN(G1347gat));
  NAND2_X1  g635(.A1(new_n386_), .A2(new_n383_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n837_), .A2(new_n352_), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n508_), .B(new_n838_), .C1(new_n780_), .C2(new_n717_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n839_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n840_));
  INV_X1    g639(.A(new_n276_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n840_), .B1(new_n841_), .B2(new_n839_), .ZN(new_n842_));
  AOI21_X1  g641(.A(KEYINPUT62), .B1(new_n839_), .B2(G169gat), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(KEYINPUT124), .ZN(G1348gat));
  NAND2_X1  g644(.A1(new_n781_), .A2(new_n838_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(G176gat), .B1(new_n847_), .B2(new_n649_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n776_), .A2(new_n352_), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n837_), .A2(new_n477_), .A3(new_n277_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n848_), .B1(new_n849_), .B2(new_n850_), .ZN(G1349gat));
  NOR3_X1   g650(.A1(new_n846_), .A2(new_n567_), .A3(new_n267_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n849_), .A2(new_n566_), .A3(new_n383_), .A4(new_n386_), .ZN(new_n853_));
  INV_X1    g652(.A(G183gat), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n852_), .B1(new_n853_), .B2(new_n854_), .ZN(G1350gat));
  OAI21_X1  g654(.A(G190gat), .B1(new_n846_), .B2(new_n552_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n575_), .A2(new_n268_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n856_), .B1(new_n846_), .B2(new_n857_), .ZN(G1351gat));
  NOR4_X1   g657(.A1(new_n628_), .A2(new_n385_), .A3(new_n346_), .A4(new_n359_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n793_), .A2(new_n859_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n860_), .A2(new_n650_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(new_n250_), .ZN(G1352gat));
  INV_X1    g661(.A(new_n860_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n649_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT125), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n865_), .B2(G204gat), .ZN(new_n866_));
  XNOR2_X1  g665(.A(KEYINPUT125), .B(G204gat), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n866_), .B1(new_n864_), .B2(new_n867_), .ZN(G1353gat));
  NOR2_X1   g667(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n869_));
  AND2_X1   g668(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n870_));
  NOR4_X1   g669(.A1(new_n860_), .A2(new_n567_), .A3(new_n869_), .A4(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n863_), .A2(new_n566_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n871_), .B1(new_n872_), .B2(new_n869_), .ZN(G1354gat));
  AND3_X1   g672(.A1(new_n863_), .A2(G218gat), .A3(new_n553_), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n860_), .A2(KEYINPUT126), .A3(new_n574_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n875_), .A2(G218gat), .ZN(new_n876_));
  OAI21_X1  g675(.A(KEYINPUT126), .B1(new_n860_), .B2(new_n574_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n874_), .B1(new_n876_), .B2(new_n877_), .ZN(G1355gat));
endmodule


