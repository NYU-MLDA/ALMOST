//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 1 0 0 0 0 1 0 1 0 0 1 0 1 1 0 1 0 1 0 1 0 0 0 0 0 0 1 1 1 0 1 0 0 0 0 1 1 0 1 0 0 1 0 0 1 0 1 0 0 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n654_, new_n655_, new_n656_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n708_, new_n709_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n754_,
    new_n755_, new_n757_, new_n758_, new_n759_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n839_, new_n840_, new_n841_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n854_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n893_, new_n894_,
    new_n895_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_;
  INV_X1    g000(.A(KEYINPUT68), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT6), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT65), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT65), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT6), .ZN(new_n206_));
  AND2_X1   g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  AND3_X1   g006(.A1(new_n204_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n207_), .B1(new_n204_), .B2(new_n206_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  OAI22_X1  g009(.A1(KEYINPUT66), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT66), .B1(KEYINPUT67), .B2(KEYINPUT7), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  OAI221_X1 g012(.A(KEYINPUT66), .B1(KEYINPUT67), .B2(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n202_), .B1(new_n210_), .B2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n204_), .A2(new_n206_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n207_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n204_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  AND2_X1   g020(.A1(new_n213_), .A2(new_n214_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n221_), .A2(new_n222_), .A3(KEYINPUT68), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT8), .ZN(new_n224_));
  XOR2_X1   g023(.A(G85gat), .B(G92gat), .Z(new_n225_));
  NAND4_X1  g024(.A1(new_n216_), .A2(new_n223_), .A3(new_n224_), .A4(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT69), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  XOR2_X1   g027(.A(KEYINPUT70), .B(KEYINPUT6), .Z(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(new_n207_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n222_), .A2(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n229_), .A2(new_n207_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n225_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT8), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n214_), .B(new_n213_), .C1(new_n208_), .C2(new_n209_), .ZN(new_n235_));
  AOI21_X1  g034(.A(KEYINPUT8), .B1(new_n235_), .B2(new_n202_), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n236_), .A2(KEYINPUT69), .A3(new_n225_), .A4(new_n223_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n228_), .A2(new_n234_), .A3(new_n237_), .ZN(new_n238_));
  XOR2_X1   g037(.A(KEYINPUT10), .B(G99gat), .Z(new_n239_));
  XNOR2_X1  g038(.A(KEYINPUT64), .B(G106gat), .ZN(new_n240_));
  AOI22_X1  g039(.A1(KEYINPUT9), .A2(new_n225_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G85gat), .A2(G92gat), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n241_), .B(new_n221_), .C1(KEYINPUT9), .C2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n238_), .A2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G57gat), .B(G64gat), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT71), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT11), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G71gat), .B(G78gat), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT11), .ZN(new_n252_));
  OR3_X1    g051(.A1(new_n247_), .A2(new_n252_), .A3(new_n250_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n244_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT72), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT12), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n256_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n254_), .B1(new_n238_), .B2(new_n243_), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT12), .B1(new_n260_), .B2(KEYINPUT72), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G230gat), .A2(G233gat), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n238_), .A2(new_n254_), .A3(new_n243_), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n259_), .A2(new_n261_), .A3(new_n262_), .A4(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n256_), .A2(new_n263_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n262_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G120gat), .B(G148gat), .ZN(new_n268_));
  INV_X1    g067(.A(G204gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT5), .ZN(new_n271_));
  INV_X1    g070(.A(G176gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n264_), .A2(new_n267_), .A3(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT73), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n264_), .A2(KEYINPUT73), .A3(new_n267_), .A4(new_n273_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n264_), .A2(new_n267_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n273_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n278_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT13), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT13), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n278_), .A2(new_n284_), .A3(new_n281_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT15), .ZN(new_n288_));
  INV_X1    g087(.A(G29gat), .ZN(new_n289_));
  INV_X1    g088(.A(G36gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G29gat), .A2(G36gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(G43gat), .ZN(new_n294_));
  INV_X1    g093(.A(G43gat), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n291_), .A2(new_n295_), .A3(new_n292_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n294_), .A2(G50gat), .A3(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(G50gat), .B1(new_n294_), .B2(new_n296_), .ZN(new_n299_));
  NOR3_X1   g098(.A1(new_n298_), .A2(new_n299_), .A3(KEYINPUT74), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT74), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n294_), .A2(new_n296_), .ZN(new_n302_));
  INV_X1    g101(.A(G50gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n301_), .B1(new_n304_), .B2(new_n297_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n288_), .B1(new_n300_), .B2(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(KEYINPUT74), .B1(new_n298_), .B2(new_n299_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n304_), .A2(new_n301_), .A3(new_n297_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n307_), .A2(KEYINPUT15), .A3(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n306_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G15gat), .B(G22gat), .ZN(new_n312_));
  INV_X1    g111(.A(G1gat), .ZN(new_n313_));
  INV_X1    g112(.A(G8gat), .ZN(new_n314_));
  OAI21_X1  g113(.A(KEYINPUT14), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n312_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G1gat), .B(G8gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n311_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n318_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n298_), .A2(new_n299_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n319_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G229gat), .A2(G233gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n320_), .B(new_n321_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n326_), .A2(G229gat), .A3(G233gat), .ZN(new_n327_));
  OR2_X1    g126(.A1(new_n327_), .A2(KEYINPUT80), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(KEYINPUT80), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n325_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G113gat), .B(G141gat), .ZN(new_n331_));
  INV_X1    g130(.A(G169gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(G197gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n330_), .B(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n287_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G231gat), .A2(G233gat), .ZN(new_n339_));
  XOR2_X1   g138(.A(new_n318_), .B(new_n339_), .Z(new_n340_));
  XNOR2_X1  g139(.A(new_n254_), .B(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT16), .B(G183gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(G211gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G127gat), .B(G155gat), .ZN(new_n344_));
  XOR2_X1   g143(.A(new_n343_), .B(new_n344_), .Z(new_n345_));
  INV_X1    g144(.A(KEYINPUT17), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n341_), .A2(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT78), .ZN(new_n349_));
  AND2_X1   g148(.A1(new_n345_), .A2(new_n346_), .ZN(new_n350_));
  OR3_X1    g149(.A1(new_n341_), .A2(new_n347_), .A3(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n349_), .A2(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT0), .B(G57gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(G85gat), .ZN(new_n354_));
  XOR2_X1   g153(.A(G1gat), .B(G29gat), .Z(new_n355_));
  XOR2_X1   g154(.A(new_n354_), .B(new_n355_), .Z(new_n356_));
  NAND2_X1  g155(.A1(G225gat), .A2(G233gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT103), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT91), .ZN(new_n360_));
  INV_X1    g159(.A(G155gat), .ZN(new_n361_));
  INV_X1    g160(.A(G162gat), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n360_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G155gat), .A2(G162gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(KEYINPUT1), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT1), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n366_), .A2(G155gat), .A3(G162gat), .ZN(new_n367_));
  OAI21_X1  g166(.A(KEYINPUT91), .B1(G155gat), .B2(G162gat), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n363_), .A2(new_n365_), .A3(new_n367_), .A4(new_n368_), .ZN(new_n369_));
  XOR2_X1   g168(.A(G141gat), .B(G148gat), .Z(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT92), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n369_), .A2(KEYINPUT92), .A3(new_n370_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT3), .ZN(new_n378_));
  INV_X1    g177(.A(G141gat), .ZN(new_n379_));
  INV_X1    g178(.A(G148gat), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n378_), .A2(new_n379_), .A3(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n382_));
  NAND3_X1  g181(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n377_), .A2(new_n381_), .A3(new_n382_), .A4(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(KEYINPUT93), .ZN(new_n385_));
  INV_X1    g184(.A(new_n383_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n386_), .A2(new_n376_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT93), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n387_), .A2(new_n388_), .A3(new_n382_), .A4(new_n381_), .ZN(new_n389_));
  AND2_X1   g188(.A1(new_n363_), .A2(new_n368_), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n385_), .A2(new_n389_), .A3(new_n390_), .A4(new_n364_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n375_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT94), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n375_), .A2(new_n391_), .A3(KEYINPUT94), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  XOR2_X1   g195(.A(G127gat), .B(G134gat), .Z(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(G113gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(G120gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n396_), .A2(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n399_), .A2(new_n392_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT4), .ZN(new_n404_));
  INV_X1    g203(.A(new_n399_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n405_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n406_));
  OR2_X1    g205(.A1(new_n406_), .A2(KEYINPUT4), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n359_), .B1(new_n404_), .B2(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n403_), .A2(new_n358_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n356_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n409_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n356_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n406_), .A2(KEYINPUT4), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n413_), .B1(new_n403_), .B2(KEYINPUT4), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n411_), .B(new_n412_), .C1(new_n414_), .C2(new_n359_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT104), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n410_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n408_), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n418_), .A2(KEYINPUT104), .A3(new_n411_), .A4(new_n412_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(new_n419_), .ZN(new_n420_));
  XOR2_X1   g219(.A(G211gat), .B(G218gat), .Z(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT96), .B(G204gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT95), .B(G197gat), .ZN(new_n423_));
  AOI22_X1  g222(.A1(G197gat), .A2(new_n422_), .B1(new_n423_), .B2(G204gat), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT21), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n421_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  OAI22_X1  g225(.A1(G197gat), .A2(new_n422_), .B1(new_n423_), .B2(G204gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT21), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n426_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n424_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n430_), .A2(KEYINPUT21), .A3(new_n421_), .ZN(new_n431_));
  AND2_X1   g230(.A1(new_n429_), .A2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(KEYINPUT98), .B(KEYINPUT24), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n332_), .A2(new_n272_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G169gat), .A2(G176gat), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n433_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(KEYINPUT25), .B(G183gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT26), .B(G190gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT99), .ZN(new_n440_));
  AND3_X1   g239(.A1(new_n436_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n440_), .B1(new_n436_), .B2(new_n439_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G183gat), .A2(G190gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(KEYINPUT23), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT23), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n445_), .A2(G183gat), .A3(G190gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n444_), .A2(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n447_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n448_));
  NOR3_X1   g247(.A1(new_n441_), .A2(new_n442_), .A3(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT84), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n443_), .A2(new_n450_), .A3(KEYINPUT23), .ZN(new_n451_));
  OAI221_X1 g250(.A(new_n451_), .B1(G183gat), .B2(G190gat), .C1(new_n447_), .C2(new_n450_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n435_), .B(KEYINPUT83), .ZN(new_n453_));
  XOR2_X1   g252(.A(KEYINPUT86), .B(G176gat), .Z(new_n454_));
  XNOR2_X1  g253(.A(KEYINPUT22), .B(G169gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  AND3_X1   g255(.A1(new_n452_), .A2(new_n453_), .A3(new_n456_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n449_), .A2(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(KEYINPUT100), .B1(new_n432_), .B2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n429_), .A2(new_n431_), .ZN(new_n460_));
  XOR2_X1   g259(.A(KEYINPUT82), .B(G190gat), .Z(new_n461_));
  XNOR2_X1  g260(.A(KEYINPUT81), .B(G183gat), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n447_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT22), .ZN(new_n464_));
  OAI21_X1  g263(.A(G169gat), .B1(new_n464_), .B2(KEYINPUT85), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n332_), .A2(KEYINPUT22), .ZN(new_n466_));
  OAI211_X1 g265(.A(new_n454_), .B(new_n465_), .C1(KEYINPUT85), .C2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n463_), .A2(new_n453_), .A3(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n453_), .A2(KEYINPUT24), .A3(new_n434_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n447_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT84), .ZN(new_n471_));
  OR2_X1    g270(.A1(new_n434_), .A2(KEYINPUT24), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n469_), .A2(new_n471_), .A3(new_n451_), .A4(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT26), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(G190gat), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n475_), .B1(new_n461_), .B2(new_n474_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n477_), .B1(new_n462_), .B2(KEYINPUT25), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n476_), .A2(new_n478_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n468_), .B1(new_n473_), .B2(new_n479_), .ZN(new_n480_));
  OR2_X1    g279(.A1(new_n460_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT100), .ZN(new_n482_));
  OAI211_X1 g281(.A(new_n460_), .B(new_n482_), .C1(new_n457_), .C2(new_n449_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n459_), .A2(KEYINPUT20), .A3(new_n481_), .A4(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G226gat), .A2(G233gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT19), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n484_), .A2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n460_), .A2(KEYINPUT101), .A3(new_n480_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(KEYINPUT101), .B1(new_n460_), .B2(new_n480_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT102), .ZN(new_n492_));
  INV_X1    g291(.A(new_n486_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT20), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n494_), .B1(new_n432_), .B2(new_n458_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n491_), .A2(new_n492_), .A3(new_n493_), .A4(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n460_), .A2(new_n480_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT101), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n495_), .A2(new_n499_), .A3(new_n493_), .A4(new_n488_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT102), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n487_), .A2(new_n496_), .A3(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(KEYINPUT18), .B(G64gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(G92gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G8gat), .B(G36gat), .ZN(new_n505_));
  XOR2_X1   g304(.A(new_n504_), .B(new_n505_), .Z(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n502_), .B(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT27), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n491_), .A2(new_n495_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(new_n486_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n512_), .B1(new_n486_), .B2(new_n484_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(new_n507_), .ZN(new_n514_));
  OAI211_X1 g313(.A(new_n514_), .B(KEYINPUT27), .C1(new_n507_), .C2(new_n502_), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n510_), .A2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G22gat), .B(G50gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT28), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  AND3_X1   g318(.A1(new_n375_), .A2(new_n391_), .A3(KEYINPUT94), .ZN(new_n520_));
  AOI21_X1  g319(.A(KEYINPUT94), .B1(new_n375_), .B2(new_n391_), .ZN(new_n521_));
  OAI21_X1  g320(.A(KEYINPUT29), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G228gat), .A2(G233gat), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n522_), .A2(new_n523_), .A3(new_n460_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT97), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n392_), .A2(KEYINPUT29), .ZN(new_n527_));
  OAI211_X1 g326(.A(G228gat), .B(G233gat), .C1(new_n527_), .C2(new_n432_), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n522_), .A2(KEYINPUT97), .A3(new_n523_), .A4(new_n460_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n526_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n396_), .A2(KEYINPUT29), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G78gat), .B(G106gat), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n531_), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n526_), .A2(new_n535_), .A3(new_n528_), .A4(new_n529_), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n532_), .A2(new_n534_), .A3(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n534_), .B1(new_n532_), .B2(new_n536_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n519_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n532_), .A2(new_n536_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(new_n533_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n532_), .A2(new_n534_), .A3(new_n536_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n541_), .A2(new_n518_), .A3(new_n542_), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n480_), .A2(KEYINPUT30), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT88), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT30), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n468_), .B(new_n546_), .C1(new_n473_), .C2(new_n479_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  OR3_X1    g347(.A1(new_n544_), .A2(new_n545_), .A3(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n545_), .B1(new_n544_), .B2(new_n548_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G227gat), .A2(G233gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT87), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G71gat), .B(G99gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(G15gat), .B(G43gat), .Z(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n549_), .A2(new_n550_), .A3(new_n556_), .ZN(new_n557_));
  OR4_X1    g356(.A1(new_n545_), .A2(new_n544_), .A3(new_n548_), .A4(new_n556_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n399_), .B(KEYINPUT31), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT89), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT90), .ZN(new_n563_));
  NOR3_X1   g362(.A1(new_n559_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n559_), .A2(new_n560_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(KEYINPUT90), .ZN(new_n566_));
  OR2_X1    g365(.A1(new_n559_), .A2(new_n562_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n564_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  AND3_X1   g367(.A1(new_n539_), .A2(new_n543_), .A3(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n568_), .B1(new_n539_), .B2(new_n543_), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n420_), .B(new_n516_), .C1(new_n569_), .C2(new_n570_), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n506_), .A2(KEYINPUT32), .ZN(new_n572_));
  OR2_X1    g371(.A1(new_n502_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n513_), .A2(new_n572_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n417_), .A2(new_n419_), .A3(new_n573_), .A4(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n502_), .B(new_n506_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n400_), .A2(new_n358_), .A3(new_n402_), .ZN(new_n577_));
  OAI211_X1 g376(.A(new_n356_), .B(new_n577_), .C1(new_n414_), .C2(new_n358_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT33), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n415_), .A2(new_n579_), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n418_), .A2(KEYINPUT33), .A3(new_n411_), .A4(new_n412_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n576_), .A2(new_n578_), .A3(new_n580_), .A4(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n575_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n543_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n539_), .ZN(new_n585_));
  OAI211_X1 g384(.A(new_n583_), .B(new_n568_), .C1(new_n584_), .C2(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n352_), .B1(new_n571_), .B2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(G232gat), .A2(G233gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT34), .ZN(new_n589_));
  AND3_X1   g388(.A1(new_n238_), .A2(new_n243_), .A3(new_n321_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n310_), .B1(new_n238_), .B2(new_n243_), .ZN(new_n591_));
  OAI211_X1 g390(.A(KEYINPUT35), .B(new_n589_), .C1(new_n590_), .C2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n244_), .A2(new_n311_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n589_), .A2(KEYINPUT35), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n589_), .A2(KEYINPUT35), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n238_), .A2(new_n243_), .A3(new_n321_), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n593_), .A2(new_n594_), .A3(new_n595_), .A4(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT75), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n592_), .A2(new_n597_), .A3(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G190gat), .B(G218gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(G134gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(G162gat), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n602_), .A2(KEYINPUT36), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n599_), .A2(new_n604_), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n592_), .A2(new_n597_), .A3(new_n598_), .A4(new_n603_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT36), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n607_), .B1(new_n592_), .B2(new_n597_), .ZN(new_n608_));
  AOI22_X1  g407(.A1(new_n605_), .A2(new_n606_), .B1(new_n602_), .B2(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n338_), .A2(new_n587_), .A3(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(G1gat), .B1(new_n610_), .B2(new_n420_), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT105), .Z(new_n612_));
  NAND2_X1  g411(.A1(new_n571_), .A2(new_n586_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n352_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT37), .ZN(new_n615_));
  OAI21_X1  g414(.A(KEYINPUT76), .B1(new_n609_), .B2(KEYINPUT77), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n605_), .A2(new_n606_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n608_), .A2(new_n602_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT76), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n615_), .B1(new_n616_), .B2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT77), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n619_), .A2(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(KEYINPUT37), .B1(new_n624_), .B2(KEYINPUT76), .ZN(new_n625_));
  OAI211_X1 g424(.A(new_n286_), .B(new_n614_), .C1(new_n622_), .C2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT79), .ZN(new_n627_));
  OAI211_X1 g426(.A(new_n336_), .B(new_n613_), .C1(new_n626_), .C2(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n620_), .B1(new_n619_), .B2(new_n623_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n609_), .A2(KEYINPUT76), .ZN(new_n630_));
  OAI21_X1  g429(.A(KEYINPUT37), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n616_), .A2(new_n615_), .ZN(new_n632_));
  AOI22_X1  g431(.A1(new_n631_), .A2(new_n632_), .B1(new_n283_), .B2(new_n285_), .ZN(new_n633_));
  AOI21_X1  g432(.A(KEYINPUT79), .B1(new_n633_), .B2(new_n614_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n628_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n420_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n635_), .A2(new_n313_), .A3(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT38), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n638_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n612_), .A2(new_n639_), .A3(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT106), .ZN(G1324gat));
  INV_X1    g441(.A(new_n635_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n516_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(new_n314_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n643_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT107), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n646_), .B(new_n647_), .ZN(new_n648_));
  OAI21_X1  g447(.A(G8gat), .B1(new_n610_), .B2(new_n516_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT39), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n648_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT40), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n651_), .B(new_n652_), .ZN(G1325gat));
  OAI21_X1  g452(.A(G15gat), .B1(new_n610_), .B2(new_n568_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT41), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n643_), .A2(G15gat), .A3(new_n568_), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n655_), .A2(new_n656_), .ZN(G1326gat));
  NOR2_X1   g456(.A1(new_n585_), .A2(new_n584_), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n658_), .B(KEYINPUT108), .Z(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  OAI21_X1  g459(.A(G22gat), .B1(new_n610_), .B2(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT42), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n660_), .A2(G22gat), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n662_), .B1(new_n643_), .B2(new_n663_), .ZN(G1327gat));
  INV_X1    g463(.A(KEYINPUT109), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n631_), .A2(new_n665_), .A3(new_n632_), .ZN(new_n666_));
  OAI21_X1  g465(.A(KEYINPUT109), .B1(new_n622_), .B2(new_n625_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n613_), .A2(new_n666_), .A3(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(KEYINPUT43), .ZN(new_n669_));
  AOI21_X1  g468(.A(KEYINPUT43), .B1(new_n571_), .B2(new_n586_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n622_), .A2(new_n625_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n669_), .A2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n338_), .A2(new_n352_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT110), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(KEYINPUT44), .ZN(new_n677_));
  OR2_X1    g476(.A1(new_n676_), .A2(KEYINPUT44), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n673_), .A2(new_n675_), .A3(new_n677_), .A4(new_n678_), .ZN(new_n679_));
  AOI22_X1  g478(.A1(new_n668_), .A2(KEYINPUT43), .B1(new_n671_), .B2(new_n670_), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n676_), .B(KEYINPUT44), .C1(new_n680_), .C2(new_n674_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n682_), .A2(G29gat), .A3(new_n636_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n609_), .B1(new_n571_), .B2(new_n586_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n675_), .A2(new_n684_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n685_), .A2(new_n636_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n683_), .B1(G29gat), .B2(new_n686_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT111), .ZN(G1328gat));
  INV_X1    g487(.A(KEYINPUT46), .ZN(new_n689_));
  AOI21_X1  g488(.A(KEYINPUT112), .B1(new_n682_), .B2(new_n644_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT112), .ZN(new_n691_));
  AOI211_X1 g490(.A(new_n691_), .B(new_n516_), .C1(new_n679_), .C2(new_n681_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n690_), .A2(new_n692_), .A3(new_n290_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n685_), .A2(new_n290_), .A3(new_n644_), .ZN(new_n694_));
  XOR2_X1   g493(.A(new_n694_), .B(KEYINPUT45), .Z(new_n695_));
  OAI21_X1  g494(.A(new_n689_), .B1(new_n693_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n690_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n682_), .A2(KEYINPUT112), .A3(new_n644_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n697_), .A2(G36gat), .A3(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n695_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n699_), .A2(new_n700_), .A3(KEYINPUT46), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n696_), .A2(new_n701_), .ZN(G1329gat));
  INV_X1    g501(.A(new_n568_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n295_), .B1(new_n682_), .B2(new_n703_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n568_), .A2(G43gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n685_), .B2(new_n705_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g506(.A1(new_n685_), .A2(new_n303_), .A3(new_n659_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n682_), .A2(new_n658_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n708_), .B1(new_n709_), .B2(new_n303_), .ZN(G1331gat));
  NAND3_X1  g509(.A1(new_n587_), .A2(new_n287_), .A3(new_n337_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n711_), .A2(new_n671_), .ZN(new_n712_));
  AOI21_X1  g511(.A(G57gat), .B1(new_n712_), .B2(new_n636_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT113), .ZN(new_n714_));
  OR3_X1    g513(.A1(new_n711_), .A2(new_n714_), .A3(new_n619_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n714_), .B1(new_n711_), .B2(new_n619_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  OR2_X1    g516(.A1(new_n420_), .A2(KEYINPUT114), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(G57gat), .B2(new_n718_), .ZN(new_n719_));
  OR2_X1    g518(.A1(KEYINPUT114), .A2(G57gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n713_), .B1(new_n719_), .B2(new_n720_), .ZN(G1332gat));
  INV_X1    g520(.A(G64gat), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n712_), .A2(new_n722_), .A3(new_n644_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT48), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n715_), .A2(new_n716_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(new_n644_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n724_), .B1(new_n726_), .B2(G64gat), .ZN(new_n727_));
  AOI211_X1 g526(.A(KEYINPUT48), .B(new_n722_), .C1(new_n725_), .C2(new_n644_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n723_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(KEYINPUT115), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT115), .ZN(new_n731_));
  OAI211_X1 g530(.A(new_n731_), .B(new_n723_), .C1(new_n727_), .C2(new_n728_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n730_), .A2(new_n732_), .ZN(G1333gat));
  INV_X1    g532(.A(G71gat), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n712_), .A2(new_n734_), .A3(new_n703_), .ZN(new_n735_));
  OAI21_X1  g534(.A(G71gat), .B1(new_n717_), .B2(new_n568_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n736_), .A2(KEYINPUT49), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n736_), .A2(KEYINPUT49), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n735_), .B1(new_n737_), .B2(new_n738_), .ZN(G1334gat));
  INV_X1    g538(.A(G78gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n712_), .A2(new_n740_), .A3(new_n659_), .ZN(new_n741_));
  OAI21_X1  g540(.A(G78gat), .B1(new_n717_), .B2(new_n660_), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n742_), .A2(KEYINPUT116), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(KEYINPUT116), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n743_), .A2(KEYINPUT50), .A3(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(KEYINPUT50), .B1(new_n743_), .B2(new_n744_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n741_), .B1(new_n745_), .B2(new_n746_), .ZN(G1335gat));
  NOR3_X1   g546(.A1(new_n286_), .A2(new_n614_), .A3(new_n336_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n684_), .A2(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(G85gat), .B1(new_n749_), .B2(new_n636_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n673_), .A2(new_n748_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n636_), .A2(G85gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n750_), .B1(new_n751_), .B2(new_n752_), .ZN(G1336gat));
  AOI21_X1  g552(.A(G92gat), .B1(new_n749_), .B2(new_n644_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n644_), .A2(G92gat), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n751_), .B2(new_n755_), .ZN(G1337gat));
  NAND2_X1  g555(.A1(new_n751_), .A2(new_n703_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n703_), .A2(new_n239_), .ZN(new_n758_));
  AOI22_X1  g557(.A1(new_n757_), .A2(G99gat), .B1(new_n749_), .B2(new_n758_), .ZN(new_n759_));
  XOR2_X1   g558(.A(new_n759_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g559(.A1(new_n749_), .A2(new_n240_), .A3(new_n658_), .ZN(new_n761_));
  INV_X1    g560(.A(G106gat), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n762_), .B1(new_n751_), .B2(new_n658_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT52), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n763_), .A2(new_n764_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n761_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT53), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT53), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n769_), .B(new_n761_), .C1(new_n765_), .C2(new_n766_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(G1339gat));
  OAI21_X1  g570(.A(KEYINPUT117), .B1(new_n626_), .B2(new_n336_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT117), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n633_), .A2(new_n773_), .A3(new_n614_), .A4(new_n337_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n772_), .A2(new_n774_), .A3(KEYINPUT54), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n772_), .A2(new_n774_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT54), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  AND3_X1   g577(.A1(new_n259_), .A2(new_n263_), .A3(new_n261_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT118), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n779_), .A2(new_n780_), .A3(KEYINPUT55), .A4(new_n262_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT55), .ZN(new_n782_));
  OAI21_X1  g581(.A(KEYINPUT118), .B1(new_n264_), .B2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n264_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n259_), .A2(new_n261_), .A3(new_n263_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n782_), .B1(new_n785_), .B2(new_n266_), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n781_), .B(new_n783_), .C1(new_n784_), .C2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT56), .ZN(new_n788_));
  AND3_X1   g587(.A1(new_n787_), .A2(new_n788_), .A3(new_n280_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n788_), .B1(new_n787_), .B2(new_n280_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  MUX2_X1   g590(.A(new_n323_), .B(new_n326_), .S(new_n324_), .Z(new_n792_));
  MUX2_X1   g591(.A(new_n330_), .B(new_n792_), .S(new_n335_), .Z(new_n793_));
  NAND4_X1  g592(.A1(new_n791_), .A2(KEYINPUT58), .A3(new_n278_), .A4(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n781_), .A2(new_n783_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n786_), .A2(new_n784_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n280_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT56), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n787_), .A2(new_n788_), .A3(new_n280_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n798_), .A2(new_n278_), .A3(new_n793_), .A4(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT58), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  AND3_X1   g601(.A1(new_n794_), .A2(new_n671_), .A3(new_n802_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n798_), .A2(new_n278_), .A3(new_n336_), .A4(new_n799_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n282_), .A2(new_n793_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT57), .B1(new_n806_), .B2(new_n609_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT57), .ZN(new_n808_));
  AOI211_X1 g607(.A(new_n808_), .B(new_n619_), .C1(new_n804_), .C2(new_n805_), .ZN(new_n809_));
  NOR3_X1   g608(.A1(new_n803_), .A2(new_n807_), .A3(new_n809_), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n775_), .B(new_n778_), .C1(new_n810_), .C2(new_n614_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n644_), .A2(new_n420_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n811_), .A2(new_n570_), .A3(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(G113gat), .B1(new_n814_), .B2(new_n336_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT59), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n813_), .A2(new_n816_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n811_), .A2(KEYINPUT59), .A3(new_n570_), .A4(new_n812_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n337_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n815_), .B1(new_n819_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g619(.A(G120gat), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n821_), .A2(KEYINPUT60), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT60), .ZN(new_n823_));
  AOI21_X1  g622(.A(G120gat), .B1(new_n287_), .B2(new_n823_), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n813_), .A2(new_n822_), .A3(new_n824_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n825_), .A2(KEYINPUT119), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT119), .ZN(new_n827_));
  NOR4_X1   g626(.A1(new_n813_), .A2(new_n827_), .A3(new_n822_), .A4(new_n824_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n286_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n829_));
  OAI22_X1  g628(.A1(new_n826_), .A2(new_n828_), .B1(new_n829_), .B2(new_n821_), .ZN(G1341gat));
  INV_X1    g629(.A(G127gat), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n831_), .B1(new_n813_), .B2(new_n352_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT120), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  OAI211_X1 g633(.A(KEYINPUT120), .B(new_n831_), .C1(new_n813_), .C2(new_n352_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  AOI211_X1 g635(.A(new_n831_), .B(new_n352_), .C1(new_n817_), .C2(new_n818_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n836_), .A2(new_n837_), .ZN(G1342gat));
  AOI21_X1  g637(.A(G134gat), .B1(new_n814_), .B2(new_n619_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n671_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n840_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n839_), .B1(new_n841_), .B2(G134gat), .ZN(G1343gat));
  NAND2_X1  g641(.A1(new_n806_), .A2(new_n609_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n808_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n806_), .A2(KEYINPUT57), .A3(new_n609_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n794_), .A2(new_n802_), .A3(new_n671_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n844_), .A2(new_n845_), .A3(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n352_), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n848_), .A2(new_n775_), .A3(new_n778_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n812_), .A2(new_n569_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n336_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n287_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g654(.A1(new_n851_), .A2(new_n614_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(KEYINPUT61), .B(G155gat), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n856_), .B(new_n857_), .ZN(G1346gat));
  AND3_X1   g657(.A1(new_n666_), .A2(new_n667_), .A3(G162gat), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n851_), .A2(new_n859_), .ZN(new_n860_));
  NOR3_X1   g659(.A1(new_n849_), .A2(new_n609_), .A3(new_n850_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(G162gat), .B2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT121), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT121), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n860_), .B(new_n864_), .C1(G162gat), .C2(new_n861_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n863_), .A2(new_n865_), .ZN(G1347gat));
  NOR2_X1   g665(.A1(new_n516_), .A2(new_n636_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n868_), .A2(new_n568_), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n811_), .A2(new_n336_), .A3(new_n660_), .A4(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(G169gat), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(KEYINPUT122), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT122), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n870_), .A2(new_n873_), .A3(G169gat), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n872_), .A2(KEYINPUT62), .A3(new_n874_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n811_), .A2(new_n660_), .A3(new_n869_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n877_), .A2(new_n336_), .A3(new_n455_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT62), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n871_), .A2(KEYINPUT122), .A3(new_n879_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n875_), .A2(new_n878_), .A3(new_n880_), .ZN(G1348gat));
  OAI21_X1  g680(.A(new_n454_), .B1(new_n876_), .B2(new_n286_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT123), .ZN(new_n883_));
  OR2_X1    g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n882_), .A2(new_n883_), .ZN(new_n885_));
  AND3_X1   g684(.A1(new_n811_), .A2(new_n570_), .A3(new_n867_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n286_), .A2(new_n272_), .ZN(new_n887_));
  AOI22_X1  g686(.A1(new_n884_), .A2(new_n885_), .B1(new_n886_), .B2(new_n887_), .ZN(G1349gat));
  AOI21_X1  g687(.A(new_n462_), .B1(new_n886_), .B2(new_n614_), .ZN(new_n889_));
  OR2_X1    g688(.A1(new_n352_), .A2(new_n437_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n889_), .B1(new_n877_), .B2(new_n891_), .ZN(G1350gat));
  OAI21_X1  g691(.A(G190gat), .B1(new_n876_), .B2(new_n840_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n619_), .A2(new_n438_), .ZN(new_n894_));
  XOR2_X1   g693(.A(new_n894_), .B(KEYINPUT124), .Z(new_n895_));
  OAI21_X1  g694(.A(new_n893_), .B1(new_n876_), .B2(new_n895_), .ZN(G1351gat));
  INV_X1    g695(.A(new_n569_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n868_), .A2(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n849_), .A2(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n336_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g701(.A1(new_n900_), .A2(new_n287_), .ZN(new_n903_));
  MUX2_X1   g702(.A(new_n422_), .B(G204gat), .S(new_n903_), .Z(G1353gat));
  AND3_X1   g703(.A1(new_n772_), .A2(new_n774_), .A3(KEYINPUT54), .ZN(new_n905_));
  AOI21_X1  g704(.A(KEYINPUT54), .B1(new_n772_), .B2(new_n774_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  AOI211_X1 g706(.A(new_n352_), .B(new_n899_), .C1(new_n907_), .C2(new_n848_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT125), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT126), .ZN(new_n910_));
  NAND2_X1  g709(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n911_));
  NAND4_X1  g710(.A1(new_n908_), .A2(new_n909_), .A3(new_n910_), .A4(new_n911_), .ZN(new_n912_));
  NAND4_X1  g711(.A1(new_n811_), .A2(new_n614_), .A3(new_n898_), .A4(new_n911_), .ZN(new_n913_));
  OAI21_X1  g712(.A(KEYINPUT126), .B1(new_n913_), .B2(KEYINPUT125), .ZN(new_n914_));
  NOR2_X1   g713(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n915_), .B1(new_n913_), .B2(KEYINPUT125), .ZN(new_n916_));
  AND3_X1   g715(.A1(new_n912_), .A2(new_n914_), .A3(new_n916_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n916_), .B1(new_n912_), .B2(new_n914_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n917_), .A2(new_n918_), .ZN(G1354gat));
  NAND3_X1  g718(.A1(new_n811_), .A2(new_n619_), .A3(new_n898_), .ZN(new_n920_));
  OR2_X1    g719(.A1(new_n920_), .A2(KEYINPUT127), .ZN(new_n921_));
  INV_X1    g720(.A(G218gat), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n920_), .A2(KEYINPUT127), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n921_), .A2(new_n922_), .A3(new_n923_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n900_), .A2(G218gat), .A3(new_n671_), .ZN(new_n925_));
  AND2_X1   g724(.A1(new_n924_), .A2(new_n925_), .ZN(G1355gat));
endmodule


