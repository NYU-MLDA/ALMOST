//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 1 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0 0 0 1 1 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 0 0 0 0 1 0 1 0 1 1 1 1 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n706_,
    new_n707_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n744_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n833_, new_n834_, new_n836_, new_n837_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n853_, new_n854_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n902_, new_n904_, new_n905_, new_n906_,
    new_n908_, new_n909_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_, new_n920_;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G85gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT0), .B(G57gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n207_), .B1(new_n208_), .B2(KEYINPUT1), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT1), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n210_), .A2(KEYINPUT89), .A3(G155gat), .A4(G162gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT89), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n212_), .B1(new_n207_), .B2(KEYINPUT1), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n209_), .A2(new_n211_), .A3(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(G141gat), .ZN(new_n215_));
  INV_X1    g014(.A(G148gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n215_), .A2(new_n216_), .A3(KEYINPUT88), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT88), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n218_), .B1(G141gat), .B2(G148gat), .ZN(new_n219_));
  AOI22_X1  g018(.A1(new_n217_), .A2(new_n219_), .B1(G141gat), .B2(G148gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n214_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(G134gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(G127gat), .ZN(new_n223_));
  INV_X1    g022(.A(G127gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(G134gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n223_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(G120gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(G113gat), .ZN(new_n228_));
  INV_X1    g027(.A(G113gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(G120gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n226_), .A2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G127gat), .B(G134gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G113gat), .B(G120gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n232_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT2), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n237_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n239_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n241_));
  OAI21_X1  g040(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n238_), .A2(new_n240_), .A3(new_n241_), .A4(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n208_), .ZN(new_n244_));
  AND2_X1   g043(.A1(new_n244_), .A2(new_n207_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n221_), .A2(new_n236_), .A3(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT86), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n226_), .A2(new_n231_), .ZN(new_n249_));
  AOI22_X1  g048(.A1(new_n223_), .A2(new_n225_), .B1(new_n228_), .B2(new_n230_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n248_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n248_), .B1(new_n226_), .B2(new_n231_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  AOI22_X1  g053(.A1(new_n214_), .A2(new_n220_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n255_));
  OAI211_X1 g054(.A(KEYINPUT99), .B(new_n247_), .C1(new_n254_), .C2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n255_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT99), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n252_), .B1(new_n236_), .B2(new_n248_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n257_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n256_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G225gat), .A2(G233gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT100), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n261_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n267_), .B1(new_n256_), .B2(new_n260_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n257_), .A2(new_n259_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n263_), .B1(new_n269_), .B2(KEYINPUT4), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n268_), .A2(new_n270_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n206_), .B1(new_n266_), .B2(new_n271_), .ZN(new_n272_));
  OAI211_X1 g071(.A(new_n265_), .B(new_n205_), .C1(new_n268_), .C2(new_n270_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G169gat), .A2(G176gat), .ZN(new_n275_));
  AND3_X1   g074(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n276_));
  AOI21_X1  g075(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT80), .ZN(new_n279_));
  INV_X1    g078(.A(G183gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(KEYINPUT80), .A2(G183gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n278_), .B1(new_n283_), .B2(G190gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(KEYINPUT22), .B(G169gat), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT84), .ZN(new_n286_));
  INV_X1    g085(.A(G176gat), .ZN(new_n287_));
  AND3_X1   g086(.A1(new_n285_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n286_), .B1(new_n285_), .B2(new_n287_), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n275_), .B(new_n284_), .C1(new_n288_), .C2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT81), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n291_), .B1(new_n280_), .B2(KEYINPUT25), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT25), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n293_), .A2(KEYINPUT81), .A3(G183gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n281_), .A2(KEYINPUT25), .A3(new_n282_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT26), .B(G190gat), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n295_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT82), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n295_), .A2(new_n296_), .A3(KEYINPUT82), .A4(new_n297_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(G169gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(new_n287_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n304_), .A2(KEYINPUT24), .A3(new_n275_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT83), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT24), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n307_), .A2(new_n303_), .A3(new_n287_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n306_), .B1(new_n278_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G183gat), .A2(G190gat), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT23), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n313_));
  AND4_X1   g112(.A1(new_n306_), .A2(new_n308_), .A3(new_n312_), .A4(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n305_), .B1(new_n309_), .B2(new_n314_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n290_), .B1(new_n302_), .B2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT30), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT87), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n259_), .B(KEYINPUT31), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(G99gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G227gat), .A2(G233gat), .ZN(new_n322_));
  INV_X1    g121(.A(G15gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(G71gat), .ZN(new_n325_));
  OR2_X1    g124(.A1(new_n321_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n321_), .A2(new_n325_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT85), .B(G43gat), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n326_), .A2(new_n327_), .A3(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n329_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n319_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n332_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n334_), .A2(new_n318_), .A3(new_n330_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n274_), .B1(new_n333_), .B2(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n278_), .B1(G183gat), .B2(G190gat), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT94), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT22), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n339_), .A2(G169gat), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n303_), .A2(KEYINPUT22), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n338_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n303_), .A2(KEYINPUT22), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n339_), .A2(G169gat), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n343_), .A2(new_n344_), .A3(KEYINPUT94), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n342_), .A2(new_n287_), .A3(new_n345_), .ZN(new_n346_));
  AND3_X1   g145(.A1(new_n346_), .A2(KEYINPUT95), .A3(new_n275_), .ZN(new_n347_));
  AOI21_X1  g146(.A(KEYINPUT95), .B1(new_n346_), .B2(new_n275_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n337_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  OR2_X1    g148(.A1(G197gat), .A2(G204gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G197gat), .A2(G204gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT21), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n350_), .A2(KEYINPUT21), .A3(new_n351_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G211gat), .B(G218gat), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n354_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  OR2_X1    g156(.A1(new_n355_), .A2(new_n356_), .ZN(new_n358_));
  AND2_X1   g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT25), .B(G183gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT93), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(new_n297_), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n362_), .A2(new_n278_), .A3(new_n305_), .A4(new_n308_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n349_), .A2(new_n359_), .A3(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G226gat), .A2(G233gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT20), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT96), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n308_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(KEYINPUT83), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n278_), .A2(new_n306_), .A3(new_n308_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n374_), .A2(new_n300_), .A3(new_n305_), .A4(new_n301_), .ZN(new_n375_));
  AOI211_X1 g174(.A(new_n370_), .B(new_n359_), .C1(new_n375_), .C2(new_n290_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n357_), .A2(new_n358_), .ZN(new_n377_));
  AOI21_X1  g176(.A(KEYINPUT96), .B1(new_n316_), .B2(new_n377_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n364_), .B(new_n369_), .C1(new_n376_), .C2(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n359_), .B1(new_n349_), .B2(new_n363_), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT20), .B1(new_n316_), .B2(new_n377_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n367_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  XOR2_X1   g181(.A(G8gat), .B(G36gat), .Z(new_n383_));
  XNOR2_X1  g182(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G64gat), .B(G92gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n379_), .A2(new_n382_), .A3(new_n387_), .ZN(new_n388_));
  NOR3_X1   g187(.A1(new_n380_), .A2(new_n381_), .A3(new_n367_), .ZN(new_n389_));
  OAI211_X1 g188(.A(KEYINPUT20), .B(new_n364_), .C1(new_n376_), .C2(new_n378_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n389_), .B1(new_n367_), .B2(new_n390_), .ZN(new_n391_));
  OAI211_X1 g190(.A(KEYINPUT27), .B(new_n388_), .C1(new_n391_), .C2(new_n387_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT27), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n379_), .A2(new_n382_), .A3(new_n387_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n387_), .B1(new_n379_), .B2(new_n382_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n393_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n392_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT29), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n377_), .B1(new_n255_), .B2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n399_), .A2(G228gat), .A3(G233gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G228gat), .A2(G233gat), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n377_), .B(new_n401_), .C1(new_n255_), .C2(new_n398_), .ZN(new_n402_));
  XOR2_X1   g201(.A(G78gat), .B(G106gat), .Z(new_n403_));
  AND3_X1   g202(.A1(new_n400_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n403_), .B1(new_n400_), .B2(new_n402_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n255_), .A2(new_n398_), .ZN(new_n407_));
  XOR2_X1   g206(.A(G22gat), .B(G50gat), .Z(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT28), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n407_), .B(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n410_), .B1(new_n405_), .B2(KEYINPUT90), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT91), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT91), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n413_), .B(new_n410_), .C1(new_n405_), .C2(KEYINPUT90), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n406_), .B1(new_n412_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n412_), .A2(new_n406_), .A3(new_n414_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n397_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n336_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n274_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n417_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n422_), .B1(new_n423_), .B2(new_n415_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n424_), .A2(new_n397_), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT98), .B1(new_n394_), .B2(new_n395_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n379_), .A2(new_n382_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n387_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT98), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n429_), .A2(new_n430_), .A3(new_n388_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n264_), .B1(new_n269_), .B2(KEYINPUT4), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n268_), .A2(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n264_), .B1(new_n256_), .B2(new_n260_), .ZN(new_n434_));
  NOR3_X1   g233(.A1(new_n433_), .A2(new_n205_), .A3(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n273_), .A2(KEYINPUT33), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n261_), .A2(KEYINPUT4), .ZN(new_n437_));
  INV_X1    g236(.A(new_n270_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT33), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n439_), .A2(new_n440_), .A3(new_n265_), .A4(new_n205_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n435_), .B1(new_n436_), .B2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n426_), .A2(new_n431_), .A3(new_n442_), .ZN(new_n443_));
  AND2_X1   g242(.A1(new_n387_), .A2(KEYINPUT32), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n379_), .A2(new_n382_), .A3(new_n445_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n274_), .B(new_n446_), .C1(new_n391_), .C2(new_n445_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n443_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n418_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT101), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n425_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n418_), .B1(new_n443_), .B2(new_n447_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT101), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n333_), .A2(new_n335_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n421_), .B1(new_n455_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT79), .ZN(new_n459_));
  XOR2_X1   g258(.A(G15gat), .B(G22gat), .Z(new_n460_));
  XNOR2_X1  g259(.A(KEYINPUT75), .B(G1gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(KEYINPUT76), .B(G8gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n460_), .B1(new_n463_), .B2(KEYINPUT14), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G1gat), .B(G8gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G29gat), .B(G36gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(KEYINPUT73), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G43gat), .B(G50gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n459_), .B1(new_n467_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n470_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n469_), .B(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n466_), .A2(new_n474_), .A3(KEYINPUT79), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n472_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G229gat), .A2(G233gat), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n467_), .A2(new_n471_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n476_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n474_), .A2(KEYINPUT15), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT15), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n471_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n481_), .A2(new_n483_), .ZN(new_n484_));
  AOI22_X1  g283(.A1(new_n475_), .A2(new_n472_), .B1(new_n484_), .B2(new_n467_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n480_), .B1(new_n485_), .B2(new_n478_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G113gat), .B(G141gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G169gat), .B(G197gat), .ZN(new_n488_));
  XOR2_X1   g287(.A(new_n487_), .B(new_n488_), .Z(new_n489_));
  NAND2_X1  g288(.A1(new_n486_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n489_), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n480_), .B(new_n491_), .C1(new_n485_), .C2(new_n478_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n458_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT13), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G99gat), .A2(G106gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(KEYINPUT6), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT6), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n499_), .A2(G99gat), .A3(G106gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n498_), .A2(new_n500_), .ZN(new_n501_));
  XOR2_X1   g300(.A(KEYINPUT10), .B(G99gat), .Z(new_n502_));
  INV_X1    g301(.A(G106gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  XOR2_X1   g303(.A(KEYINPUT64), .B(G85gat), .Z(new_n505_));
  OR2_X1    g304(.A1(G85gat), .A2(G92gat), .ZN(new_n506_));
  AOI22_X1  g305(.A1(new_n505_), .A2(G92gat), .B1(KEYINPUT9), .B2(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT65), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n501_), .B(new_n504_), .C1(new_n507_), .C2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT8), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT67), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n501_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n498_), .A2(new_n500_), .A3(KEYINPUT67), .ZN(new_n514_));
  INV_X1    g313(.A(G99gat), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n515_), .A2(new_n503_), .A3(KEYINPUT66), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT7), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT7), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n518_), .A2(new_n515_), .A3(new_n503_), .A4(KEYINPUT66), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n513_), .A2(new_n514_), .A3(new_n517_), .A4(new_n519_), .ZN(new_n520_));
  XOR2_X1   g319(.A(G85gat), .B(G92gat), .Z(new_n521_));
  AOI21_X1  g320(.A(new_n511_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n511_), .ZN(new_n523_));
  AND2_X1   g322(.A1(new_n517_), .A2(new_n519_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n523_), .B1(new_n524_), .B2(new_n501_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n510_), .B1(new_n522_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT68), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT68), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n528_), .B(new_n510_), .C1(new_n522_), .C2(new_n525_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G57gat), .B(G64gat), .ZN(new_n531_));
  OR2_X1    g330(.A1(new_n531_), .A2(KEYINPUT11), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(KEYINPUT11), .ZN(new_n533_));
  XOR2_X1   g332(.A(G71gat), .B(G78gat), .Z(new_n534_));
  NAND3_X1  g333(.A1(new_n532_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n535_));
  OR2_X1    g334(.A1(new_n533_), .A2(new_n534_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n530_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n537_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n527_), .A2(new_n529_), .A3(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G230gat), .A2(G233gat), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n541_), .A2(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n543_), .B1(new_n530_), .B2(new_n537_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT12), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n540_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT69), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n510_), .B(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n522_), .A2(new_n525_), .ZN(new_n550_));
  OAI211_X1 g349(.A(KEYINPUT12), .B(new_n539_), .C1(new_n549_), .C2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n545_), .A2(new_n547_), .A3(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n544_), .A2(new_n552_), .ZN(new_n553_));
  XOR2_X1   g352(.A(G176gat), .B(G204gat), .Z(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT71), .ZN(new_n555_));
  XOR2_X1   g354(.A(G120gat), .B(G148gat), .Z(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n553_), .A2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n544_), .A2(new_n552_), .A3(new_n559_), .ZN(new_n562_));
  AND3_X1   g361(.A1(new_n561_), .A2(KEYINPUT72), .A3(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(KEYINPUT72), .B1(new_n561_), .B2(new_n562_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n496_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n561_), .A2(new_n562_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT72), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n561_), .A2(KEYINPUT72), .A3(new_n562_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n568_), .A2(new_n569_), .A3(KEYINPUT13), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n565_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G231gat), .A2(G233gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n537_), .B(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(new_n467_), .ZN(new_n574_));
  XOR2_X1   g373(.A(G127gat), .B(G155gat), .Z(new_n575_));
  XNOR2_X1  g374(.A(G183gat), .B(G211gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n579_), .A2(KEYINPUT77), .A3(KEYINPUT17), .ZN(new_n580_));
  OAI211_X1 g379(.A(new_n574_), .B(new_n580_), .C1(KEYINPUT17), .C2(new_n579_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n581_), .B1(new_n574_), .B2(new_n580_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G190gat), .B(G218gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G134gat), .B(G162gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  XOR2_X1   g384(.A(new_n585_), .B(KEYINPUT36), .Z(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(G232gat), .A2(G233gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT34), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n549_), .A2(new_n550_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n590_), .B1(new_n481_), .B2(new_n483_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n471_), .B1(new_n527_), .B2(new_n529_), .ZN(new_n592_));
  OAI211_X1 g391(.A(KEYINPUT35), .B(new_n589_), .C1(new_n591_), .C2(new_n592_), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n549_), .A2(new_n550_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT35), .ZN(new_n595_));
  INV_X1    g394(.A(new_n589_), .ZN(new_n596_));
  AOI22_X1  g395(.A1(new_n594_), .A2(new_n484_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(new_n595_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n592_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n597_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n587_), .B1(new_n593_), .B2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n585_), .A2(KEYINPUT36), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n593_), .A2(new_n601_), .A3(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(KEYINPUT74), .B(KEYINPUT37), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n603_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n606_), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n593_), .A2(new_n601_), .A3(new_n604_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n608_), .B1(new_n609_), .B2(new_n602_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n582_), .B1(new_n607_), .B2(new_n610_), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n495_), .A2(new_n571_), .A3(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n422_), .A2(new_n461_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  XOR2_X1   g413(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n571_), .A2(new_n493_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n617_), .A2(new_n582_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n454_), .ZN(new_n619_));
  OAI22_X1  g418(.A1(new_n453_), .A2(KEYINPUT101), .B1(new_n424_), .B2(new_n397_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n457_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(new_n420_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n603_), .A2(new_n605_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n618_), .A2(new_n622_), .A3(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT103), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n623_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n458_), .A2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n628_), .A2(KEYINPUT103), .A3(new_n618_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n626_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(G1gat), .B1(new_n631_), .B2(new_n422_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n616_), .A2(new_n632_), .ZN(G1324gat));
  INV_X1    g432(.A(new_n462_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n612_), .A2(new_n397_), .A3(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n397_), .ZN(new_n636_));
  OAI21_X1  g435(.A(G8gat), .B1(new_n624_), .B2(new_n636_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n637_), .A2(KEYINPUT39), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(KEYINPUT39), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n635_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT40), .Z(G1325gat));
  NAND3_X1  g440(.A1(new_n612_), .A2(new_n323_), .A3(new_n456_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n630_), .A2(new_n456_), .ZN(new_n643_));
  AOI21_X1  g442(.A(KEYINPUT41), .B1(new_n643_), .B2(G15gat), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT41), .ZN(new_n645_));
  AOI211_X1 g444(.A(new_n645_), .B(new_n323_), .C1(new_n630_), .C2(new_n456_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n642_), .B1(new_n644_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT104), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  OAI211_X1 g448(.A(KEYINPUT104), .B(new_n642_), .C1(new_n644_), .C2(new_n646_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(G1326gat));
  INV_X1    g450(.A(G22gat), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n612_), .A2(new_n652_), .A3(new_n418_), .ZN(new_n653_));
  OAI21_X1  g452(.A(G22gat), .B1(new_n631_), .B2(new_n449_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n654_), .A2(KEYINPUT42), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n654_), .A2(KEYINPUT42), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n653_), .B1(new_n655_), .B2(new_n656_), .ZN(G1327gat));
  INV_X1    g456(.A(KEYINPUT106), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT43), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n607_), .A2(new_n610_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n456_), .B1(new_n452_), .B2(new_n454_), .ZN(new_n662_));
  OAI211_X1 g461(.A(new_n659_), .B(new_n661_), .C1(new_n662_), .C2(new_n421_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(KEYINPUT105), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT105), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n622_), .A2(new_n665_), .A3(new_n659_), .A4(new_n661_), .ZN(new_n666_));
  OAI21_X1  g465(.A(KEYINPUT43), .B1(new_n458_), .B2(new_n660_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n664_), .A2(new_n666_), .A3(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n582_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n617_), .A2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT44), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n668_), .A2(KEYINPUT44), .A3(new_n670_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n673_), .A2(new_n274_), .A3(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(G29gat), .ZN(new_n676_));
  INV_X1    g475(.A(new_n571_), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n677_), .A2(new_n623_), .A3(new_n669_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n495_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  NOR3_X1   g479(.A1(new_n680_), .A2(G29gat), .A3(new_n422_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n658_), .B1(new_n676_), .B2(new_n682_), .ZN(new_n683_));
  AOI211_X1 g482(.A(KEYINPUT106), .B(new_n681_), .C1(new_n675_), .C2(G29gat), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n683_), .A2(new_n684_), .ZN(G1328gat));
  INV_X1    g484(.A(G36gat), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n679_), .A2(new_n686_), .A3(new_n397_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT45), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n668_), .A2(KEYINPUT44), .A3(new_n670_), .ZN(new_n689_));
  AOI21_X1  g488(.A(KEYINPUT44), .B1(new_n668_), .B2(new_n670_), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n689_), .A2(new_n690_), .A3(new_n636_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n688_), .B1(new_n691_), .B2(new_n686_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT46), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  OAI211_X1 g493(.A(new_n688_), .B(KEYINPUT46), .C1(new_n691_), .C2(new_n686_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(G1329gat));
  AND4_X1   g495(.A1(G43gat), .A2(new_n673_), .A3(new_n456_), .A4(new_n674_), .ZN(new_n697_));
  AOI21_X1  g496(.A(G43gat), .B1(new_n679_), .B2(new_n456_), .ZN(new_n698_));
  OAI21_X1  g497(.A(KEYINPUT47), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n689_), .A2(new_n690_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n700_), .A2(G43gat), .A3(new_n456_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT47), .ZN(new_n702_));
  INV_X1    g501(.A(new_n698_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n701_), .A2(new_n702_), .A3(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n699_), .A2(new_n704_), .ZN(G1330gat));
  AOI21_X1  g504(.A(G50gat), .B1(new_n679_), .B2(new_n418_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n418_), .A2(G50gat), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n700_), .B2(new_n707_), .ZN(G1331gat));
  NOR3_X1   g507(.A1(new_n458_), .A2(new_n493_), .A3(new_n571_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n709_), .A2(new_n611_), .ZN(new_n710_));
  AOI21_X1  g509(.A(G57gat), .B1(new_n710_), .B2(new_n274_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT107), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n571_), .A2(new_n582_), .A3(new_n493_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n628_), .A2(new_n713_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n714_), .A2(G57gat), .A3(new_n274_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n712_), .A2(new_n715_), .ZN(G1332gat));
  INV_X1    g515(.A(G64gat), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n710_), .A2(new_n717_), .A3(new_n397_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n714_), .A2(new_n397_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(KEYINPUT108), .B(KEYINPUT48), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n719_), .A2(G64gat), .A3(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n719_), .B2(G64gat), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n718_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT109), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n723_), .B(new_n724_), .ZN(G1333gat));
  INV_X1    g524(.A(G71gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n726_), .B1(new_n714_), .B2(new_n456_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(KEYINPUT110), .B(KEYINPUT49), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n727_), .B(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n710_), .A2(new_n726_), .A3(new_n456_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1334gat));
  INV_X1    g530(.A(G78gat), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n732_), .B1(new_n714_), .B2(new_n418_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n733_), .B(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n710_), .A2(new_n732_), .A3(new_n418_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(G1335gat));
  AND3_X1   g536(.A1(new_n709_), .A2(new_n627_), .A3(new_n582_), .ZN(new_n738_));
  AOI21_X1  g537(.A(G85gat), .B1(new_n738_), .B2(new_n274_), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n571_), .A2(new_n669_), .A3(new_n493_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n668_), .A2(new_n740_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n274_), .A2(new_n505_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n739_), .B1(new_n741_), .B2(new_n742_), .ZN(G1336gat));
  INV_X1    g542(.A(G92gat), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n738_), .A2(new_n744_), .A3(new_n397_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n741_), .A2(new_n397_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n745_), .B1(new_n746_), .B2(new_n744_), .ZN(G1337gat));
  AOI21_X1  g546(.A(new_n515_), .B1(new_n741_), .B2(new_n456_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n738_), .A2(new_n456_), .A3(new_n502_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT112), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n748_), .A2(new_n750_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n751_), .B(new_n752_), .ZN(G1338gat));
  NAND3_X1  g552(.A1(new_n738_), .A2(new_n503_), .A3(new_n418_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n668_), .A2(new_n418_), .A3(new_n740_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT52), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n755_), .A2(new_n756_), .A3(G106gat), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n755_), .B2(G106gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n754_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(KEYINPUT53), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT53), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n761_), .B(new_n754_), .C1(new_n757_), .C2(new_n758_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(G1339gat));
  NAND4_X1  g562(.A1(new_n611_), .A2(new_n565_), .A3(new_n570_), .A4(new_n494_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT54), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n764_), .A2(KEYINPUT114), .A3(new_n765_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n766_), .B1(new_n764_), .B2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n493_), .A2(new_n562_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n552_), .A2(new_n771_), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n545_), .A2(new_n547_), .A3(KEYINPUT55), .A4(new_n551_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n547_), .A2(new_n538_), .A3(new_n551_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n543_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n772_), .A2(new_n773_), .A3(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n560_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT56), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n776_), .A2(KEYINPUT56), .A3(new_n560_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n770_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n485_), .A2(new_n478_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n476_), .A2(new_n479_), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n782_), .B(new_n491_), .C1(new_n783_), .C2(new_n478_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n490_), .A2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n786_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n623_), .B1(new_n781_), .B2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT57), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n623_), .A2(KEYINPUT57), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n792_), .B1(new_n781_), .B2(new_n787_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT116), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  AND3_X1   g594(.A1(new_n776_), .A2(KEYINPUT56), .A3(new_n560_), .ZN(new_n796_));
  AOI21_X1  g595(.A(KEYINPUT56), .B1(new_n776_), .B2(new_n560_), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n562_), .B(new_n785_), .C1(new_n796_), .C2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT58), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n660_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n785_), .A2(new_n562_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n801_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT58), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n800_), .A2(new_n803_), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n493_), .B(new_n562_), .C1(new_n796_), .C2(new_n797_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n785_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n807_), .A2(KEYINPUT116), .A3(new_n792_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n790_), .A2(new_n795_), .A3(new_n804_), .A4(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n769_), .B1(new_n809_), .B2(new_n582_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n456_), .A2(new_n274_), .A3(new_n419_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(G113gat), .B1(new_n812_), .B2(new_n493_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n813_), .B(KEYINPUT117), .ZN(new_n814_));
  OR2_X1    g613(.A1(new_n810_), .A2(new_n811_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT119), .ZN(new_n816_));
  OAI21_X1  g615(.A(KEYINPUT118), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT59), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT118), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n818_), .B1(new_n812_), .B2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n817_), .A2(new_n820_), .ZN(new_n821_));
  OAI211_X1 g620(.A(KEYINPUT118), .B(new_n818_), .C1(new_n815_), .C2(new_n816_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n494_), .A2(new_n229_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n814_), .B1(new_n823_), .B2(new_n824_), .ZN(G1340gat));
  INV_X1    g624(.A(KEYINPUT60), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT120), .B1(new_n826_), .B2(G120gat), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n227_), .B1(new_n571_), .B2(KEYINPUT60), .ZN(new_n828_));
  MUX2_X1   g627(.A(KEYINPUT120), .B(new_n827_), .S(new_n828_), .Z(new_n829_));
  NAND2_X1  g628(.A1(new_n812_), .A2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n571_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n830_), .B1(new_n831_), .B2(new_n227_), .ZN(G1341gat));
  NAND3_X1  g631(.A1(new_n812_), .A2(new_n224_), .A3(new_n669_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n582_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n833_), .B1(new_n834_), .B2(new_n224_), .ZN(G1342gat));
  NAND3_X1  g634(.A1(new_n812_), .A2(new_n222_), .A3(new_n627_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n660_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n836_), .B1(new_n837_), .B2(new_n222_), .ZN(G1343gat));
  INV_X1    g637(.A(KEYINPUT121), .ZN(new_n839_));
  NOR4_X1   g638(.A1(new_n456_), .A2(new_n422_), .A3(new_n449_), .A4(new_n397_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n839_), .B1(new_n810_), .B2(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(KEYINPUT116), .B1(new_n807_), .B2(new_n792_), .ZN(new_n843_));
  AOI211_X1 g642(.A(new_n794_), .B(new_n791_), .C1(new_n805_), .C2(new_n806_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  AOI22_X1  g644(.A1(new_n788_), .A2(new_n789_), .B1(new_n800_), .B2(new_n803_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n669_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  OAI211_X1 g646(.A(KEYINPUT121), .B(new_n840_), .C1(new_n847_), .C2(new_n769_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n842_), .A2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n493_), .ZN(new_n850_));
  XOR2_X1   g649(.A(KEYINPUT122), .B(G141gat), .Z(new_n851_));
  XNOR2_X1  g650(.A(new_n850_), .B(new_n851_), .ZN(G1344gat));
  NAND2_X1  g651(.A1(new_n849_), .A2(new_n677_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(KEYINPUT123), .B(G148gat), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n853_), .B(new_n854_), .ZN(G1345gat));
  NAND2_X1  g654(.A1(new_n795_), .A2(new_n808_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n798_), .A2(new_n799_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n661_), .B1(new_n802_), .B2(KEYINPUT58), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n627_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n859_));
  OAI22_X1  g658(.A1(new_n857_), .A2(new_n858_), .B1(new_n859_), .B2(KEYINPUT57), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n582_), .B1(new_n856_), .B2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n769_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(KEYINPUT121), .B1(new_n863_), .B2(new_n840_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n810_), .A2(new_n839_), .A3(new_n841_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n669_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(KEYINPUT124), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT124), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n849_), .A2(new_n868_), .A3(new_n669_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(KEYINPUT61), .B(G155gat), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n867_), .A2(new_n869_), .A3(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n870_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n868_), .B1(new_n849_), .B2(new_n669_), .ZN(new_n873_));
  AOI211_X1 g672(.A(KEYINPUT124), .B(new_n582_), .C1(new_n842_), .C2(new_n848_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n872_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n875_));
  AND2_X1   g674(.A1(new_n871_), .A2(new_n875_), .ZN(G1346gat));
  INV_X1    g675(.A(new_n849_), .ZN(new_n877_));
  OR3_X1    g676(.A1(new_n877_), .A2(G162gat), .A3(new_n623_), .ZN(new_n878_));
  OAI21_X1  g677(.A(G162gat), .B1(new_n877_), .B2(new_n660_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1347gat));
  NAND3_X1  g679(.A1(new_n336_), .A2(new_n449_), .A3(new_n397_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n881_), .A2(new_n494_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n863_), .A2(KEYINPUT125), .A3(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT125), .ZN(new_n884_));
  INV_X1    g683(.A(new_n882_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n810_), .B2(new_n885_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n883_), .A2(new_n886_), .A3(G169gat), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT62), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n863_), .A2(new_n342_), .A3(new_n345_), .A4(new_n882_), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n883_), .A2(new_n886_), .A3(KEYINPUT62), .A4(G169gat), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n889_), .A2(new_n890_), .A3(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT126), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n889_), .A2(KEYINPUT126), .A3(new_n890_), .A4(new_n891_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1348gat));
  NOR2_X1   g695(.A1(new_n810_), .A2(new_n881_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n677_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n898_), .B1(KEYINPUT127), .B2(new_n287_), .ZN(new_n899_));
  XOR2_X1   g698(.A(KEYINPUT127), .B(G176gat), .Z(new_n900_));
  AOI21_X1  g699(.A(new_n899_), .B1(new_n898_), .B2(new_n900_), .ZN(G1349gat));
  NAND2_X1  g700(.A1(new_n897_), .A2(new_n669_), .ZN(new_n902_));
  MUX2_X1   g701(.A(new_n361_), .B(new_n283_), .S(new_n902_), .Z(G1350gat));
  NAND3_X1  g702(.A1(new_n897_), .A2(new_n297_), .A3(new_n627_), .ZN(new_n904_));
  NOR3_X1   g703(.A1(new_n810_), .A2(new_n660_), .A3(new_n881_), .ZN(new_n905_));
  INV_X1    g704(.A(G190gat), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n904_), .B1(new_n905_), .B2(new_n906_), .ZN(G1351gat));
  NOR4_X1   g706(.A1(new_n810_), .A2(new_n456_), .A3(new_n424_), .A4(new_n636_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(new_n493_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g709(.A1(new_n908_), .A2(new_n677_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g711(.A1(new_n908_), .A2(new_n669_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n914_));
  AND2_X1   g713(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n915_));
  NOR3_X1   g714(.A1(new_n913_), .A2(new_n914_), .A3(new_n915_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n916_), .B1(new_n913_), .B2(new_n914_), .ZN(G1354gat));
  INV_X1    g716(.A(G218gat), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n908_), .A2(new_n918_), .A3(new_n627_), .ZN(new_n919_));
  AND2_X1   g718(.A1(new_n908_), .A2(new_n661_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n919_), .B1(new_n920_), .B2(new_n918_), .ZN(G1355gat));
endmodule


