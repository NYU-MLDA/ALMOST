//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 0 0 1 0 1 1 1 0 1 0 0 0 1 0 0 0 1 0 0 0 1 0 0 0 0 1 1 0 1 0 0 1 1 0 1 1 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n677_, new_n678_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n841_, new_n842_, new_n844_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n872_, new_n873_, new_n875_, new_n876_,
    new_n878_, new_n879_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n891_, new_n892_;
  NOR3_X1   g000(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n202_));
  NOR2_X1   g001(.A1(G141gat), .A2(G148gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT3), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G141gat), .A2(G148gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT2), .ZN(new_n206_));
  OAI22_X1  g005(.A1(new_n203_), .A2(new_n204_), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n205_), .B(KEYINPUT92), .ZN(new_n208_));
  AND2_X1   g007(.A1(new_n208_), .A2(new_n206_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT93), .ZN(new_n210_));
  AOI211_X1 g009(.A(new_n202_), .B(new_n207_), .C1(new_n209_), .C2(new_n210_), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n211_), .B1(new_n210_), .B2(new_n209_), .ZN(new_n212_));
  AND2_X1   g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n212_), .A2(new_n215_), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n203_), .B1(new_n213_), .B2(KEYINPUT1), .ZN(new_n217_));
  INV_X1    g016(.A(new_n215_), .ZN(new_n218_));
  OAI211_X1 g017(.A(new_n208_), .B(new_n217_), .C1(new_n218_), .C2(KEYINPUT1), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n216_), .A2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G113gat), .B(G120gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n221_), .B(KEYINPUT89), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G127gat), .B(G134gat), .ZN(new_n223_));
  XOR2_X1   g022(.A(new_n222_), .B(new_n223_), .Z(new_n224_));
  NOR2_X1   g023(.A1(new_n220_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(KEYINPUT90), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT90), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n222_), .A2(new_n227_), .A3(new_n223_), .ZN(new_n228_));
  AOI22_X1  g027(.A1(new_n216_), .A2(new_n219_), .B1(new_n226_), .B2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT4), .B1(new_n225_), .B2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G225gat), .A2(G233gat), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n229_), .A2(KEYINPUT4), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n230_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT98), .B(KEYINPUT0), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT99), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G1gat), .B(G29gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G57gat), .B(G85gat), .ZN(new_n239_));
  XOR2_X1   g038(.A(new_n238_), .B(new_n239_), .Z(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n231_), .B1(new_n225_), .B2(new_n229_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n234_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT101), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT101), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n234_), .A2(new_n245_), .A3(new_n241_), .A4(new_n242_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n234_), .A2(new_n242_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(new_n240_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n244_), .A2(new_n246_), .A3(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  XOR2_X1   g049(.A(G211gat), .B(G218gat), .Z(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT95), .B(G204gat), .ZN(new_n252_));
  INV_X1    g051(.A(G197gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT21), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n255_), .B1(G197gat), .B2(G204gat), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n251_), .B1(new_n254_), .B2(new_n256_), .ZN(new_n257_));
  MUX2_X1   g056(.A(G204gat), .B(new_n252_), .S(G197gat), .Z(new_n258_));
  OAI21_X1  g057(.A(new_n257_), .B1(new_n258_), .B2(KEYINPUT21), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n258_), .A2(KEYINPUT21), .A3(new_n251_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G169gat), .A2(G176gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT87), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G183gat), .A2(G190gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT23), .ZN(new_n266_));
  INV_X1    g065(.A(G183gat), .ZN(new_n267_));
  INV_X1    g066(.A(G190gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n264_), .B1(new_n266_), .B2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT22), .B(G169gat), .ZN(new_n271_));
  INV_X1    g070(.A(G176gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT24), .ZN(new_n274_));
  INV_X1    g073(.A(G169gat), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n274_), .A2(new_n275_), .A3(new_n272_), .ZN(new_n276_));
  AND2_X1   g075(.A1(new_n266_), .A2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT26), .B(G190gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT25), .B(G183gat), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  AOI22_X1  g080(.A1(new_n278_), .A2(new_n279_), .B1(new_n281_), .B2(new_n263_), .ZN(new_n282_));
  AOI22_X1  g081(.A1(new_n270_), .A2(new_n273_), .B1(new_n277_), .B2(new_n282_), .ZN(new_n283_));
  OR3_X1    g082(.A1(new_n262_), .A2(KEYINPUT97), .A3(new_n283_), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT97), .B1(new_n262_), .B2(new_n283_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT86), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n278_), .A2(new_n286_), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n268_), .A2(KEYINPUT26), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n279_), .B1(KEYINPUT86), .B2(new_n288_), .ZN(new_n289_));
  OAI221_X1 g088(.A(new_n277_), .B1(new_n264_), .B2(new_n280_), .C1(new_n287_), .C2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n273_), .B(KEYINPUT88), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(new_n270_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n262_), .A2(new_n290_), .A3(new_n292_), .ZN(new_n293_));
  NAND4_X1  g092(.A1(new_n284_), .A2(KEYINPUT20), .A3(new_n285_), .A4(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G226gat), .A2(G233gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT19), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n290_), .A2(new_n292_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(new_n261_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n262_), .A2(new_n283_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n299_), .A2(new_n300_), .A3(KEYINPUT20), .ZN(new_n301_));
  OR2_X1    g100(.A1(new_n301_), .A2(new_n296_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n297_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G8gat), .B(G36gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT18), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(G64gat), .ZN(new_n306_));
  INV_X1    g105(.A(G92gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n303_), .A2(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n297_), .A2(new_n308_), .A3(new_n302_), .ZN(new_n311_));
  AND2_X1   g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  OR2_X1    g111(.A1(new_n312_), .A2(KEYINPUT27), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n301_), .A2(new_n296_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n314_), .B1(new_n294_), .B2(new_n296_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(new_n309_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n316_), .A2(KEYINPUT27), .A3(new_n311_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n250_), .A2(new_n313_), .A3(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n226_), .A2(new_n228_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G71gat), .B(G99gat), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  AND3_X1   g120(.A1(new_n290_), .A2(new_n292_), .A3(KEYINPUT30), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(KEYINPUT30), .B1(new_n290_), .B2(new_n292_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G227gat), .A2(G233gat), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n323_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n326_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n328_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G15gat), .B(G43gat), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n327_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n330_), .B1(new_n327_), .B2(new_n329_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n321_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n333_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n335_), .A2(new_n320_), .A3(new_n331_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT91), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n334_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n338_));
  AND2_X1   g137(.A1(new_n338_), .A2(KEYINPUT31), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT31), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n334_), .A2(new_n336_), .A3(new_n337_), .A4(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n319_), .B1(new_n339_), .B2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT94), .B(KEYINPUT28), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  AND2_X1   g144(.A1(new_n216_), .A2(new_n219_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT29), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n345_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  NOR3_X1   g147(.A1(new_n220_), .A2(KEYINPUT29), .A3(new_n344_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G22gat), .B(G50gat), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NOR3_X1   g150(.A1(new_n348_), .A2(new_n349_), .A3(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n346_), .A2(new_n347_), .A3(new_n345_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n344_), .B1(new_n220_), .B2(KEYINPUT29), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n350_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT96), .ZN(new_n356_));
  NOR3_X1   g155(.A1(new_n352_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(G228gat), .ZN(new_n358_));
  INV_X1    g157(.A(G233gat), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  OAI211_X1 g160(.A(new_n361_), .B(new_n261_), .C1(new_n346_), .C2(new_n347_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n347_), .B1(new_n216_), .B2(new_n219_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n360_), .B1(new_n363_), .B2(new_n262_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G78gat), .B(G106gat), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n362_), .A2(new_n364_), .A3(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n362_), .A2(new_n364_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(new_n365_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n357_), .A2(new_n367_), .A3(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n367_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n356_), .B1(new_n352_), .B2(new_n355_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n351_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n353_), .A2(new_n350_), .A3(new_n354_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n373_), .A2(KEYINPUT96), .A3(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n371_), .A2(new_n372_), .A3(new_n375_), .ZN(new_n376_));
  AND2_X1   g175(.A1(new_n370_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n338_), .A2(KEYINPUT31), .ZN(new_n378_));
  INV_X1    g177(.A(new_n319_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n378_), .A2(new_n379_), .A3(new_n341_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n343_), .A2(new_n377_), .A3(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n370_), .A2(new_n376_), .ZN(new_n382_));
  AND3_X1   g181(.A1(new_n378_), .A2(new_n379_), .A3(new_n341_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n379_), .B1(new_n378_), .B2(new_n341_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n382_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n318_), .B1(new_n381_), .B2(new_n385_), .ZN(new_n386_));
  NOR3_X1   g185(.A1(new_n225_), .A2(new_n229_), .A3(new_n231_), .ZN(new_n387_));
  OR2_X1    g186(.A1(new_n387_), .A2(new_n240_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n232_), .B1(new_n230_), .B2(new_n233_), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n311_), .B(new_n310_), .C1(new_n388_), .C2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT100), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n391_), .A2(KEYINPUT33), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n390_), .B1(new_n248_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n392_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n247_), .A2(new_n240_), .A3(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n303_), .B1(KEYINPUT32), .B2(new_n308_), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n308_), .A2(KEYINPUT32), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n396_), .B1(new_n315_), .B2(new_n397_), .ZN(new_n398_));
  AOI22_X1  g197(.A1(new_n393_), .A2(new_n395_), .B1(new_n249_), .B2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n343_), .A2(new_n382_), .A3(new_n380_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  OR2_X1    g200(.A1(new_n386_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G230gat), .A2(G233gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(KEYINPUT64), .ZN(new_n404_));
  XNOR2_X1  g203(.A(KEYINPUT10), .B(G99gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(KEYINPUT65), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n406_), .A2(G106gat), .ZN(new_n407_));
  AND3_X1   g206(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n408_));
  AOI21_X1  g207(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT66), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G99gat), .A2(G106gat), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT6), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT66), .ZN(new_n414_));
  NAND3_X1  g213(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n413_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  AND2_X1   g215(.A1(new_n410_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G85gat), .A2(G92gat), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n418_), .A2(KEYINPUT9), .ZN(new_n419_));
  AND2_X1   g218(.A1(G85gat), .A2(G92gat), .ZN(new_n420_));
  NOR2_X1   g219(.A1(G85gat), .A2(G92gat), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n419_), .B1(new_n422_), .B2(KEYINPUT9), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n417_), .A2(new_n423_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n407_), .A2(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NOR3_X1   g226(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT69), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n413_), .A2(new_n430_), .A3(new_n415_), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT69), .B1(new_n408_), .B2(new_n409_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n429_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT67), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n434_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n435_));
  INV_X1    g234(.A(G85gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(new_n307_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n437_), .A2(KEYINPUT67), .A3(new_n418_), .ZN(new_n438_));
  AND2_X1   g237(.A1(new_n435_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n433_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT70), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n433_), .A2(new_n439_), .A3(KEYINPUT70), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(KEYINPUT8), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT8), .ZN(new_n445_));
  AND3_X1   g244(.A1(new_n435_), .A2(new_n438_), .A3(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n429_), .A2(new_n410_), .A3(new_n416_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT68), .ZN(new_n448_));
  AND3_X1   g247(.A1(new_n446_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n448_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n425_), .B1(new_n444_), .B2(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G57gat), .B(G64gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT11), .ZN(new_n454_));
  OR2_X1    g253(.A1(new_n453_), .A2(KEYINPUT11), .ZN(new_n455_));
  XNOR2_X1  g254(.A(KEYINPUT71), .B(G71gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(G78gat), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n456_), .A2(G78gat), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n454_), .B(new_n455_), .C1(new_n458_), .C2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n459_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n461_), .A2(KEYINPUT11), .A3(new_n453_), .A4(new_n457_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  AND2_X1   g262(.A1(new_n452_), .A2(new_n463_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n452_), .A2(new_n463_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n404_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT12), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n467_), .B1(new_n452_), .B2(new_n463_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n404_), .B1(new_n452_), .B2(new_n463_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n425_), .ZN(new_n470_));
  AND3_X1   g269(.A1(new_n433_), .A2(KEYINPUT70), .A3(new_n439_), .ZN(new_n471_));
  AOI21_X1  g270(.A(KEYINPUT70), .B1(new_n433_), .B2(new_n439_), .ZN(new_n472_));
  NOR3_X1   g271(.A1(new_n471_), .A2(new_n472_), .A3(new_n445_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n446_), .A2(new_n447_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(KEYINPUT68), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n446_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n470_), .B1(new_n473_), .B2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT72), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n463_), .A2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n460_), .A2(new_n462_), .A3(KEYINPUT72), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n467_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n478_), .A2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n468_), .A2(new_n469_), .A3(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n466_), .A2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G176gat), .B(G204gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT74), .ZN(new_n487_));
  XOR2_X1   g286(.A(G120gat), .B(G148gat), .Z(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n485_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n491_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n466_), .A2(new_n484_), .A3(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT13), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n492_), .A2(KEYINPUT13), .A3(new_n494_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G229gat), .A2(G233gat), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(KEYINPUT79), .B(G8gat), .ZN(new_n503_));
  INV_X1    g302(.A(G1gat), .ZN(new_n504_));
  OAI21_X1  g303(.A(KEYINPUT14), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G15gat), .B(G22gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  OR2_X1    g306(.A1(new_n507_), .A2(KEYINPUT80), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G1gat), .B(G8gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n507_), .A2(KEYINPUT80), .ZN(new_n510_));
  AND3_X1   g309(.A1(new_n508_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n509_), .B1(new_n508_), .B2(new_n510_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G29gat), .B(G36gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G43gat), .B(G50gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  NOR3_X1   g315(.A1(new_n511_), .A2(new_n512_), .A3(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n508_), .A2(new_n510_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n509_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n508_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n515_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n502_), .B1(new_n517_), .B2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n520_), .A2(new_n521_), .A3(new_n515_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT75), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n515_), .B(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT15), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT15), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n516_), .A2(new_n525_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n515_), .A2(KEYINPUT75), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n528_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n527_), .A2(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n511_), .A2(new_n512_), .ZN(new_n533_));
  OAI211_X1 g332(.A(new_n524_), .B(new_n501_), .C1(new_n532_), .C2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G113gat), .B(G141gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(G197gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(KEYINPUT82), .B(G169gat), .ZN(new_n537_));
  XOR2_X1   g336(.A(new_n536_), .B(new_n537_), .Z(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n523_), .A2(new_n534_), .A3(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT84), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n540_), .A2(new_n541_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT83), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n523_), .A2(new_n534_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n544_), .B1(new_n545_), .B2(new_n538_), .ZN(new_n546_));
  AOI211_X1 g345(.A(KEYINPUT83), .B(new_n539_), .C1(new_n523_), .C2(new_n534_), .ZN(new_n547_));
  OAI22_X1  g346(.A1(new_n542_), .A2(new_n543_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT85), .ZN(new_n549_));
  OR2_X1    g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n549_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  AND3_X1   g351(.A1(new_n402_), .A2(new_n500_), .A3(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G232gat), .A2(G233gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT34), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n555_), .A2(KEYINPUT35), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n556_), .B1(new_n452_), .B2(new_n515_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n557_), .B1(new_n452_), .B2(new_n532_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n558_), .A2(KEYINPUT35), .A3(new_n555_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G134gat), .B(G162gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT78), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G190gat), .B(G218gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n565_), .A2(KEYINPUT36), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n555_), .A2(KEYINPUT35), .ZN(new_n567_));
  OAI211_X1 g366(.A(new_n557_), .B(new_n567_), .C1(new_n452_), .C2(new_n532_), .ZN(new_n568_));
  AND3_X1   g367(.A1(new_n559_), .A2(new_n566_), .A3(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n565_), .B(KEYINPUT36), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n570_), .B1(new_n559_), .B2(new_n568_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  OR2_X1    g371(.A1(new_n572_), .A2(KEYINPUT37), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(KEYINPUT37), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G231gat), .A2(G233gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n533_), .B(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n480_), .A2(new_n481_), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n578_), .B(KEYINPUT81), .Z(new_n579_));
  AND2_X1   g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT17), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G127gat), .B(G155gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT16), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(G183gat), .ZN(new_n584_));
  INV_X1    g383(.A(G211gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  NOR3_X1   g385(.A1(new_n580_), .A2(new_n581_), .A3(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n587_), .B1(new_n577_), .B2(new_n579_), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n577_), .A2(new_n463_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n577_), .A2(new_n463_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n586_), .B(KEYINPUT17), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n589_), .A2(new_n590_), .A3(new_n591_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n588_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n575_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n553_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n597_), .A2(new_n504_), .A3(new_n249_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT38), .ZN(new_n599_));
  INV_X1    g398(.A(new_n572_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n402_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n500_), .A2(new_n548_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT102), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n603_), .A2(new_n593_), .ZN(new_n604_));
  OR2_X1    g403(.A1(new_n604_), .A2(KEYINPUT103), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(KEYINPUT103), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n601_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(G1gat), .B1(new_n607_), .B2(new_n250_), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n608_), .A2(KEYINPUT104), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n608_), .A2(KEYINPUT104), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n599_), .B1(new_n609_), .B2(new_n610_), .ZN(G1324gat));
  NAND2_X1  g410(.A1(new_n313_), .A2(new_n317_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n597_), .A2(new_n503_), .A3(new_n612_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n601_), .A2(new_n605_), .A3(new_n606_), .A4(new_n612_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT39), .ZN(new_n615_));
  AND3_X1   g414(.A1(new_n614_), .A2(new_n615_), .A3(G8gat), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n615_), .B1(new_n614_), .B2(G8gat), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n613_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n618_), .B(KEYINPUT40), .Z(G1325gat));
  NOR2_X1   g418(.A1(new_n383_), .A2(new_n384_), .ZN(new_n620_));
  NOR3_X1   g419(.A1(new_n596_), .A2(G15gat), .A3(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT105), .ZN(new_n622_));
  OAI21_X1  g421(.A(G15gat), .B1(new_n607_), .B2(new_n620_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(KEYINPUT41), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n623_), .A2(KEYINPUT41), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n622_), .A2(new_n624_), .A3(new_n625_), .ZN(G1326gat));
  OR3_X1    g425(.A1(new_n596_), .A2(G22gat), .A3(new_n382_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n601_), .A2(new_n605_), .A3(new_n606_), .A4(new_n377_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT42), .ZN(new_n629_));
  AND3_X1   g428(.A1(new_n628_), .A2(new_n629_), .A3(G22gat), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n629_), .B1(new_n628_), .B2(G22gat), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n627_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  XOR2_X1   g431(.A(new_n632_), .B(KEYINPUT106), .Z(G1327gat));
  NOR2_X1   g432(.A1(new_n593_), .A2(new_n600_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n553_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(G29gat), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n249_), .A2(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT108), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n636_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT107), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n575_), .B1(new_n386_), .B2(new_n401_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT43), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  OAI211_X1 g443(.A(KEYINPUT43), .B(new_n575_), .C1(new_n386_), .C2(new_n401_), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n644_), .A2(new_n594_), .A3(new_n603_), .A4(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT44), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n250_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n593_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n649_), .A2(KEYINPUT44), .A3(new_n603_), .A4(new_n645_), .ZN(new_n650_));
  AOI211_X1 g449(.A(new_n641_), .B(new_n637_), .C1(new_n648_), .C2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n646_), .A2(new_n647_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n652_), .A2(new_n249_), .A3(new_n650_), .ZN(new_n653_));
  AOI21_X1  g452(.A(KEYINPUT107), .B1(new_n653_), .B2(G29gat), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n640_), .B1(new_n651_), .B2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(KEYINPUT109), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT109), .ZN(new_n657_));
  OAI211_X1 g456(.A(new_n657_), .B(new_n640_), .C1(new_n651_), .C2(new_n654_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(G1328gat));
  INV_X1    g458(.A(KEYINPUT46), .ZN(new_n660_));
  XOR2_X1   g459(.A(new_n612_), .B(KEYINPUT110), .Z(new_n661_));
  NOR3_X1   g460(.A1(new_n635_), .A2(G36gat), .A3(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT45), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n652_), .A2(new_n612_), .A3(new_n650_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(G36gat), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n660_), .B1(new_n663_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT45), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n662_), .B(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n669_), .A2(KEYINPUT46), .A3(new_n665_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n667_), .A2(new_n670_), .ZN(G1329gat));
  INV_X1    g470(.A(new_n620_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n652_), .A2(G43gat), .A3(new_n672_), .A4(new_n650_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n635_), .A2(new_n620_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n673_), .B1(G43gat), .B2(new_n674_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g475(.A(G50gat), .B1(new_n636_), .B2(new_n377_), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n652_), .A2(G50gat), .A3(new_n377_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n677_), .B1(new_n678_), .B2(new_n650_), .ZN(G1331gat));
  INV_X1    g478(.A(new_n552_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(new_n593_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n681_), .A2(new_n500_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n601_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n684_), .A2(G57gat), .A3(new_n249_), .ZN(new_n685_));
  XOR2_X1   g484(.A(new_n685_), .B(KEYINPUT112), .Z(new_n686_));
  NOR2_X1   g485(.A1(new_n500_), .A2(new_n548_), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n402_), .A2(new_n595_), .A3(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(G57gat), .B1(new_n688_), .B2(new_n249_), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n689_), .B(KEYINPUT111), .Z(new_n690_));
  NOR2_X1   g489(.A1(new_n686_), .A2(new_n690_), .ZN(G1332gat));
  INV_X1    g490(.A(G64gat), .ZN(new_n692_));
  INV_X1    g491(.A(new_n661_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n688_), .A2(new_n692_), .A3(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(G64gat), .B1(new_n683_), .B2(new_n661_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT113), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n695_), .B(new_n696_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n697_), .A2(KEYINPUT48), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n697_), .A2(KEYINPUT48), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n694_), .B1(new_n698_), .B2(new_n699_), .ZN(G1333gat));
  INV_X1    g499(.A(G71gat), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n688_), .A2(new_n701_), .A3(new_n672_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT49), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n684_), .A2(new_n672_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n703_), .B1(new_n704_), .B2(G71gat), .ZN(new_n705_));
  OAI211_X1 g504(.A(new_n703_), .B(G71gat), .C1(new_n683_), .C2(new_n620_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n702_), .B1(new_n705_), .B2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT114), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  OAI211_X1 g509(.A(KEYINPUT114), .B(new_n702_), .C1(new_n705_), .C2(new_n707_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1334gat));
  OAI21_X1  g511(.A(G78gat), .B1(new_n683_), .B2(new_n382_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT50), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n382_), .A2(G78gat), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT115), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n688_), .A2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n714_), .A2(new_n717_), .ZN(G1335gat));
  NAND3_X1  g517(.A1(new_n649_), .A2(new_n645_), .A3(new_n687_), .ZN(new_n719_));
  OAI21_X1  g518(.A(G85gat), .B1(new_n719_), .B2(new_n250_), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n402_), .A2(new_n634_), .A3(new_n687_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n721_), .A2(new_n436_), .A3(new_n249_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(G1336gat));
  OAI21_X1  g522(.A(G92gat), .B1(new_n719_), .B2(new_n661_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n721_), .A2(new_n307_), .A3(new_n612_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(G1337gat));
  NOR2_X1   g525(.A1(new_n620_), .A2(new_n406_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n721_), .A2(new_n727_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT116), .ZN(new_n729_));
  OAI21_X1  g528(.A(G99gat), .B1(new_n719_), .B2(new_n620_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g531(.A(G106gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n721_), .A2(new_n733_), .A3(new_n377_), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n649_), .A2(new_n377_), .A3(new_n645_), .A4(new_n687_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(KEYINPUT117), .B(KEYINPUT52), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n735_), .A2(G106gat), .A3(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n735_), .B2(G106gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n734_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g539(.A(KEYINPUT122), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT57), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n572_), .A2(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n501_), .B1(new_n517_), .B2(new_n522_), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n524_), .B(new_n502_), .C1(new_n532_), .C2(new_n533_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n744_), .A2(new_n745_), .A3(new_n538_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT120), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n746_), .B(new_n747_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n540_), .B(new_n541_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n748_), .A2(new_n749_), .A3(new_n495_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n548_), .A2(new_n494_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT55), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n484_), .A2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n452_), .A2(new_n463_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n468_), .A2(new_n754_), .A3(new_n483_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(new_n404_), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n468_), .A2(new_n469_), .A3(KEYINPUT55), .A4(new_n483_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n753_), .A2(new_n756_), .A3(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT118), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n753_), .A2(new_n756_), .A3(KEYINPUT118), .A4(new_n757_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n760_), .A2(new_n491_), .A3(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT56), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n493_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n765_), .A2(KEYINPUT56), .A3(new_n761_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n751_), .B1(new_n764_), .B2(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n750_), .B1(new_n767_), .B2(KEYINPUT119), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT119), .ZN(new_n769_));
  AOI211_X1 g568(.A(new_n769_), .B(new_n751_), .C1(new_n764_), .C2(new_n766_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n743_), .B1(new_n768_), .B2(new_n770_), .ZN(new_n771_));
  AND3_X1   g570(.A1(new_n749_), .A2(new_n748_), .A3(new_n494_), .ZN(new_n772_));
  AND3_X1   g571(.A1(new_n765_), .A2(KEYINPUT56), .A3(new_n761_), .ZN(new_n773_));
  AOI21_X1  g572(.A(KEYINPUT56), .B1(new_n765_), .B2(new_n761_), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n772_), .B(KEYINPUT58), .C1(new_n773_), .C2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT121), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n772_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT58), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n764_), .A2(new_n766_), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n781_), .A2(KEYINPUT121), .A3(KEYINPUT58), .A4(new_n772_), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n777_), .A2(new_n780_), .A3(new_n782_), .A4(new_n575_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n771_), .A2(new_n783_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n548_), .A2(new_n494_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n785_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(new_n769_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n781_), .A2(KEYINPUT119), .A3(new_n785_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n787_), .A2(new_n788_), .A3(new_n750_), .ZN(new_n789_));
  AOI21_X1  g588(.A(KEYINPUT57), .B1(new_n789_), .B2(new_n600_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n741_), .B1(new_n784_), .B2(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n600_), .B1(new_n768_), .B2(new_n770_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(new_n742_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n793_), .A2(KEYINPUT122), .A3(new_n771_), .A4(new_n783_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n791_), .A2(new_n794_), .A3(new_n594_), .ZN(new_n795_));
  NOR3_X1   g594(.A1(new_n681_), .A2(new_n499_), .A3(new_n575_), .ZN(new_n796_));
  XOR2_X1   g595(.A(new_n796_), .B(KEYINPUT54), .Z(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT123), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n795_), .A2(KEYINPUT123), .A3(new_n797_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n612_), .A2(new_n250_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n672_), .A2(new_n382_), .A3(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n800_), .A2(new_n548_), .A3(new_n801_), .A4(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(G113gat), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(KEYINPUT124), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT124), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n805_), .A2(new_n809_), .A3(new_n806_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n594_), .B1(new_n784_), .B2(new_n790_), .ZN(new_n811_));
  AOI211_X1 g610(.A(KEYINPUT59), .B(new_n803_), .C1(new_n797_), .C2(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n800_), .A2(new_n801_), .A3(new_n804_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n812_), .B1(new_n813_), .B2(KEYINPUT59), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n680_), .A2(new_n806_), .ZN(new_n815_));
  AOI22_X1  g614(.A1(new_n808_), .A2(new_n810_), .B1(new_n814_), .B2(new_n815_), .ZN(G1340gat));
  INV_X1    g615(.A(KEYINPUT125), .ZN(new_n817_));
  INV_X1    g616(.A(G120gat), .ZN(new_n818_));
  AOI21_X1  g617(.A(KEYINPUT60), .B1(new_n499_), .B2(new_n818_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n818_), .A2(KEYINPUT60), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n817_), .B1(new_n813_), .B2(new_n822_), .ZN(new_n823_));
  AND3_X1   g622(.A1(new_n795_), .A2(KEYINPUT123), .A3(new_n797_), .ZN(new_n824_));
  AOI21_X1  g623(.A(KEYINPUT123), .B1(new_n795_), .B2(new_n797_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n826_), .A2(KEYINPUT125), .A3(new_n804_), .A4(new_n821_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n823_), .A2(new_n827_), .ZN(new_n828_));
  AOI211_X1 g627(.A(new_n500_), .B(new_n812_), .C1(new_n813_), .C2(KEYINPUT59), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n828_), .B1(new_n829_), .B2(new_n818_), .ZN(G1341gat));
  INV_X1    g629(.A(new_n813_), .ZN(new_n831_));
  INV_X1    g630(.A(G127gat), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n831_), .A2(new_n832_), .A3(new_n593_), .ZN(new_n833_));
  AOI211_X1 g632(.A(new_n594_), .B(new_n812_), .C1(new_n813_), .C2(KEYINPUT59), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n833_), .B1(new_n834_), .B2(new_n832_), .ZN(G1342gat));
  INV_X1    g634(.A(G134gat), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n831_), .A2(new_n836_), .A3(new_n572_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n575_), .ZN(new_n838_));
  AOI211_X1 g637(.A(new_n838_), .B(new_n812_), .C1(new_n813_), .C2(KEYINPUT59), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n837_), .B1(new_n839_), .B2(new_n836_), .ZN(G1343gat));
  NOR3_X1   g639(.A1(new_n693_), .A2(new_n250_), .A3(new_n381_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n826_), .A2(new_n548_), .A3(new_n841_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g642(.A1(new_n826_), .A2(new_n499_), .A3(new_n841_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g644(.A1(new_n826_), .A2(new_n593_), .A3(new_n841_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(KEYINPUT61), .B(G155gat), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n846_), .B(new_n847_), .ZN(G1346gat));
  NAND3_X1  g647(.A1(new_n826_), .A2(new_n575_), .A3(new_n841_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(G162gat), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n600_), .A2(G162gat), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n826_), .A2(new_n841_), .A3(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n852_), .ZN(G1347gat));
  NAND2_X1  g652(.A1(new_n797_), .A2(new_n811_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n661_), .A2(new_n249_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n672_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n856_), .A2(new_n377_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n854_), .A2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n548_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(G169gat), .ZN(new_n861_));
  XNOR2_X1  g660(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n863_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n860_), .A2(G169gat), .A3(new_n862_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n271_), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n864_), .B(new_n865_), .C1(new_n866_), .C2(new_n860_), .ZN(G1348gat));
  AOI21_X1  g666(.A(G176gat), .B1(new_n859_), .B2(new_n499_), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n824_), .A2(new_n825_), .A3(new_n377_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n856_), .A2(new_n272_), .A3(new_n500_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n868_), .B1(new_n869_), .B2(new_n870_), .ZN(G1349gat));
  NOR3_X1   g670(.A1(new_n858_), .A2(new_n594_), .A3(new_n279_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n869_), .A2(new_n593_), .A3(new_n672_), .A4(new_n855_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n872_), .B1(new_n873_), .B2(new_n267_), .ZN(G1350gat));
  OAI21_X1  g673(.A(G190gat), .B1(new_n858_), .B2(new_n838_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n572_), .A2(new_n278_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(new_n858_), .B2(new_n876_), .ZN(G1351gat));
  NOR3_X1   g676(.A1(new_n661_), .A2(new_n249_), .A3(new_n381_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n826_), .A2(new_n548_), .A3(new_n878_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(G197gat), .ZN(G1352gat));
  NAND4_X1  g679(.A1(new_n800_), .A2(new_n499_), .A3(new_n801_), .A4(new_n878_), .ZN(new_n881_));
  MUX2_X1   g680(.A(new_n252_), .B(G204gat), .S(new_n881_), .Z(G1353gat));
  INV_X1    g681(.A(KEYINPUT63), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n593_), .B1(new_n883_), .B2(new_n585_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(KEYINPUT127), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n826_), .A2(new_n878_), .A3(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n883_), .A2(new_n585_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n886_), .B(new_n887_), .ZN(G1354gat));
  NAND3_X1  g687(.A1(new_n826_), .A2(new_n575_), .A3(new_n878_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(G218gat), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n600_), .A2(G218gat), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n826_), .A2(new_n878_), .A3(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n890_), .A2(new_n892_), .ZN(G1355gat));
endmodule


