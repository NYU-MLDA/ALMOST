//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 0 0 1 1 0 1 0 1 1 0 1 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 1 0 1 1 0 0 1 0 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n588_, new_n589_, new_n590_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n645_, new_n646_,
    new_n647_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n657_, new_n658_, new_n659_, new_n661_,
    new_n662_, new_n663_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n768_, new_n769_, new_n770_, new_n771_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n779_, new_n780_,
    new_n782_, new_n783_, new_n784_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n806_, new_n807_, new_n809_,
    new_n810_, new_n812_, new_n813_, new_n814_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n834_, new_n835_;
  INV_X1    g000(.A(G169gat), .ZN(new_n202_));
  INV_X1    g001(.A(G176gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n205_), .A2(KEYINPUT24), .A3(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT25), .B(G183gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT26), .B(G190gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT23), .ZN(new_n212_));
  INV_X1    g011(.A(G183gat), .ZN(new_n213_));
  INV_X1    g012(.A(G190gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n212_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n216_));
  AND2_X1   g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT24), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n206_), .A2(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(KEYINPUT74), .B1(new_n217_), .B2(new_n219_), .ZN(new_n220_));
  AND4_X1   g019(.A1(KEYINPUT74), .A2(new_n215_), .A3(new_n219_), .A4(new_n216_), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n208_), .B(new_n211_), .C1(new_n220_), .C2(new_n221_), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n215_), .B(new_n216_), .C1(G183gat), .C2(G190gat), .ZN(new_n223_));
  OR2_X1    g022(.A1(new_n223_), .A2(KEYINPUT75), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT22), .B(G169gat), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n204_), .B1(new_n225_), .B2(new_n203_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n223_), .A2(KEYINPUT75), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n224_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n222_), .A2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT30), .ZN(new_n230_));
  OR2_X1    g029(.A1(G127gat), .A2(G134gat), .ZN(new_n231_));
  INV_X1    g030(.A(G113gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G127gat), .A2(G134gat), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n231_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  AND2_X1   g033(.A1(G127gat), .A2(G134gat), .ZN(new_n235_));
  NOR2_X1   g034(.A1(G127gat), .A2(G134gat), .ZN(new_n236_));
  OAI21_X1  g035(.A(G113gat), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  AND3_X1   g036(.A1(new_n234_), .A2(new_n237_), .A3(G120gat), .ZN(new_n238_));
  AOI21_X1  g037(.A(G120gat), .B1(new_n234_), .B2(new_n237_), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n230_), .B(new_n240_), .ZN(new_n241_));
  XOR2_X1   g040(.A(G15gat), .B(G43gat), .Z(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT31), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n241_), .B(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G71gat), .B(G99gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G227gat), .A2(G233gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n244_), .B(new_n247_), .ZN(new_n248_));
  AND2_X1   g047(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n249_));
  NOR2_X1   g048(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n250_));
  OAI22_X1  g049(.A1(new_n249_), .A2(new_n250_), .B1(G141gat), .B2(G148gat), .ZN(new_n251_));
  AND3_X1   g050(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n252_));
  AOI21_X1  g051(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n255_));
  INV_X1    g054(.A(G141gat), .ZN(new_n256_));
  INV_X1    g055(.A(G148gat), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n255_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n251_), .A2(new_n254_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT77), .ZN(new_n260_));
  INV_X1    g059(.A(G155gat), .ZN(new_n261_));
  INV_X1    g060(.A(G162gat), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n260_), .A2(new_n261_), .A3(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT77), .B1(G155gat), .B2(G162gat), .ZN(new_n264_));
  AND2_X1   g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G155gat), .A2(G162gat), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n259_), .A2(new_n265_), .A3(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(KEYINPUT1), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT1), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n269_), .A2(G155gat), .A3(G162gat), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n263_), .A2(new_n268_), .A3(new_n270_), .A4(new_n264_), .ZN(new_n271_));
  AND2_X1   g070(.A1(G141gat), .A2(G148gat), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT76), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n273_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n274_));
  OAI21_X1  g073(.A(KEYINPUT76), .B1(G141gat), .B2(G148gat), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n272_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT78), .ZN(new_n277_));
  AND3_X1   g076(.A1(new_n271_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n277_), .B1(new_n271_), .B2(new_n276_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n267_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(KEYINPUT29), .ZN(new_n281_));
  INV_X1    g080(.A(G197gat), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n282_), .A2(G204gat), .ZN(new_n283_));
  OR2_X1    g082(.A1(new_n283_), .A2(KEYINPUT81), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G211gat), .B(G218gat), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n284_), .A2(KEYINPUT21), .A3(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G197gat), .B(G204gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  OR2_X1    g087(.A1(new_n285_), .A2(KEYINPUT21), .ZN(new_n289_));
  INV_X1    g088(.A(new_n287_), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n284_), .A2(new_n290_), .A3(KEYINPUT21), .A4(new_n285_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n288_), .A2(new_n289_), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n281_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(G228gat), .ZN(new_n295_));
  INV_X1    g094(.A(G233gat), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n294_), .A2(new_n297_), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n281_), .B(new_n293_), .C1(new_n295_), .C2(new_n296_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  XOR2_X1   g099(.A(G78gat), .B(G106gat), .Z(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n298_), .A2(new_n299_), .A3(new_n301_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  XOR2_X1   g104(.A(G22gat), .B(G50gat), .Z(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT28), .ZN(new_n307_));
  OR3_X1    g106(.A1(new_n280_), .A2(KEYINPUT29), .A3(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n307_), .B1(new_n280_), .B2(KEYINPUT29), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  AND2_X1   g110(.A1(new_n311_), .A2(KEYINPUT80), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n311_), .A2(KEYINPUT80), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n305_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT82), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n304_), .A2(new_n315_), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n298_), .A2(new_n299_), .A3(KEYINPUT82), .A4(new_n301_), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n316_), .A2(new_n303_), .A3(new_n311_), .A4(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n314_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT91), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n280_), .A2(new_n240_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n238_), .A2(new_n239_), .ZN(new_n322_));
  OAI211_X1 g121(.A(new_n322_), .B(new_n267_), .C1(new_n279_), .C2(new_n278_), .ZN(new_n323_));
  AND3_X1   g122(.A1(new_n321_), .A2(KEYINPUT4), .A3(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT4), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n280_), .A2(new_n325_), .A3(new_n240_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G225gat), .A2(G233gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT90), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n326_), .A2(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n320_), .B1(new_n324_), .B2(new_n330_), .ZN(new_n331_));
  AND2_X1   g130(.A1(new_n321_), .A2(new_n323_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(new_n327_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n271_), .A2(new_n276_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(KEYINPUT78), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n271_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n322_), .B1(new_n337_), .B2(new_n267_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n328_), .B1(new_n338_), .B2(new_n325_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n321_), .A2(KEYINPUT4), .A3(new_n323_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n339_), .A2(KEYINPUT91), .A3(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n331_), .A2(new_n333_), .A3(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G1gat), .B(G29gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(KEYINPUT93), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G57gat), .B(G85gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT92), .B(KEYINPUT0), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n346_), .B(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n342_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT98), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n342_), .A2(KEYINPUT98), .A3(new_n350_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n331_), .A2(new_n333_), .A3(new_n341_), .A4(new_n349_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT97), .ZN(new_n356_));
  NOR3_X1   g155(.A1(new_n324_), .A2(new_n320_), .A3(new_n330_), .ZN(new_n357_));
  AOI21_X1  g156(.A(KEYINPUT91), .B1(new_n339_), .B2(new_n340_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT97), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n359_), .A2(new_n360_), .A3(new_n333_), .A4(new_n349_), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n353_), .A2(new_n354_), .A3(new_n356_), .A4(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT20), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n363_), .B1(new_n229_), .B2(new_n293_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT87), .ZN(new_n365_));
  XOR2_X1   g164(.A(KEYINPUT84), .B(KEYINPUT24), .Z(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(new_n206_), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n367_), .A2(new_n211_), .A3(new_n217_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT85), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n369_), .B1(new_n366_), .B2(new_n204_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(KEYINPUT84), .B(KEYINPUT24), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n205_), .A2(new_n371_), .A3(KEYINPUT85), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n370_), .A2(new_n207_), .A3(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n368_), .A2(new_n373_), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n217_), .B(KEYINPUT86), .C1(G183gat), .C2(G190gat), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT86), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n223_), .A2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n375_), .A2(new_n226_), .A3(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n374_), .A2(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n365_), .B1(new_n379_), .B2(new_n293_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n223_), .B(KEYINPUT86), .ZN(new_n381_));
  AOI22_X1  g180(.A1(new_n381_), .A2(new_n226_), .B1(new_n373_), .B2(new_n368_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n382_), .A2(KEYINPUT87), .A3(new_n292_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n364_), .A2(new_n380_), .A3(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G226gat), .A2(G233gat), .ZN(new_n385_));
  XOR2_X1   g184(.A(new_n385_), .B(KEYINPUT83), .Z(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT19), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n384_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n379_), .A2(new_n293_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n222_), .A2(new_n292_), .A3(new_n228_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n390_), .A2(KEYINPUT20), .A3(new_n387_), .A4(new_n391_), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n389_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n382_), .A2(KEYINPUT96), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT96), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n379_), .A2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n394_), .A2(new_n396_), .A3(new_n292_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n388_), .B1(new_n397_), .B2(new_n364_), .ZN(new_n398_));
  AND4_X1   g197(.A1(KEYINPUT20), .A2(new_n390_), .A3(new_n388_), .A4(new_n391_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G64gat), .B(G92gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(G36gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(KEYINPUT88), .B(KEYINPUT18), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(KEYINPUT89), .B(G8gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT32), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  MUX2_X1   g207(.A(new_n393_), .B(new_n400_), .S(new_n408_), .Z(new_n409_));
  NAND2_X1  g208(.A1(new_n362_), .A2(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n349_), .B1(new_n332_), .B2(new_n329_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n340_), .A2(new_n327_), .A3(new_n326_), .ZN(new_n412_));
  AND3_X1   g211(.A1(new_n411_), .A2(KEYINPUT95), .A3(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(KEYINPUT95), .B1(new_n411_), .B2(new_n412_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  AND3_X1   g214(.A1(new_n389_), .A2(new_n392_), .A3(new_n406_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n406_), .B1(new_n389_), .B2(new_n392_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT33), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n355_), .B1(KEYINPUT94), .B2(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(KEYINPUT94), .B(KEYINPUT33), .ZN(new_n421_));
  OR2_X1    g220(.A1(new_n355_), .A2(new_n421_), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n415_), .A2(new_n418_), .A3(new_n420_), .A4(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n319_), .B1(new_n410_), .B2(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n406_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n425_));
  OAI211_X1 g224(.A(KEYINPUT27), .B(new_n425_), .C1(new_n393_), .C2(new_n406_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT27), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n427_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n426_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n319_), .ZN(new_n430_));
  NOR3_X1   g229(.A1(new_n429_), .A2(new_n430_), .A3(new_n362_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n248_), .B1(new_n424_), .B2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(KEYINPUT99), .ZN(new_n433_));
  INV_X1    g232(.A(new_n248_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n362_), .ZN(new_n435_));
  OR3_X1    g234(.A1(new_n429_), .A2(KEYINPUT100), .A3(new_n319_), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT100), .B1(new_n429_), .B2(new_n319_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n434_), .A2(new_n435_), .A3(new_n436_), .A4(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT99), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n439_), .B(new_n248_), .C1(new_n424_), .C2(new_n431_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n433_), .A2(new_n438_), .A3(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G57gat), .B(G64gat), .ZN(new_n443_));
  OR2_X1    g242(.A1(new_n443_), .A2(KEYINPUT11), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(KEYINPUT11), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G71gat), .B(G78gat), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n444_), .A2(new_n445_), .A3(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n443_), .A2(new_n446_), .A3(KEYINPUT11), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G15gat), .B(G22gat), .ZN(new_n451_));
  INV_X1    g250(.A(G1gat), .ZN(new_n452_));
  INV_X1    g251(.A(G8gat), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT14), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n451_), .A2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G1gat), .B(G8gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n455_), .B(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n450_), .B(new_n457_), .ZN(new_n458_));
  AND2_X1   g257(.A1(G231gat), .A2(G233gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  XOR2_X1   g260(.A(G127gat), .B(G155gat), .Z(new_n462_));
  XNOR2_X1  g261(.A(G183gat), .B(G211gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  XOR2_X1   g263(.A(KEYINPUT69), .B(KEYINPUT16), .Z(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n467_), .A2(KEYINPUT68), .A3(KEYINPUT17), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n461_), .A2(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n468_), .B1(KEYINPUT17), .B2(new_n467_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n460_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G29gat), .B(G36gat), .ZN(new_n474_));
  INV_X1    g273(.A(G43gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(G50gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT15), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G99gat), .A2(G106gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT6), .ZN(new_n481_));
  OAI21_X1  g280(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n482_));
  OR3_X1    g281(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n481_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n484_));
  XOR2_X1   g283(.A(G85gat), .B(G92gat), .Z(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT8), .ZN(new_n487_));
  XOR2_X1   g286(.A(KEYINPUT10), .B(G99gat), .Z(new_n488_));
  INV_X1    g287(.A(G106gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n485_), .A2(KEYINPUT9), .ZN(new_n491_));
  NAND2_X1  g290(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n492_), .A2(KEYINPUT9), .ZN(new_n493_));
  NOR2_X1   g292(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n494_));
  OAI21_X1  g293(.A(G92gat), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n490_), .A2(new_n491_), .A3(new_n495_), .A4(new_n481_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n487_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n479_), .A2(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n487_), .A2(new_n478_), .A3(new_n496_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G232gat), .A2(G233gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT34), .ZN(new_n501_));
  OAI211_X1 g300(.A(new_n498_), .B(new_n499_), .C1(KEYINPUT35), .C2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(KEYINPUT35), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n502_), .B(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G190gat), .B(G218gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(G134gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(new_n262_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT36), .ZN(new_n508_));
  OR2_X1    g307(.A1(new_n504_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT36), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n507_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n504_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n509_), .A2(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n513_), .A2(KEYINPUT37), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT37), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n515_), .B1(new_n509_), .B2(new_n512_), .ZN(new_n516_));
  OR2_X1    g315(.A1(new_n514_), .A2(new_n516_), .ZN(new_n517_));
  NOR3_X1   g316(.A1(new_n442_), .A2(new_n473_), .A3(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n478_), .B(new_n457_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G229gat), .A2(G233gat), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n478_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n522_), .A2(new_n457_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n523_), .B1(new_n479_), .B2(new_n457_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n521_), .B1(new_n524_), .B2(new_n520_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G113gat), .B(G141gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(new_n202_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(new_n282_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT70), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n525_), .A2(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT71), .ZN(new_n531_));
  INV_X1    g330(.A(new_n528_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n525_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n531_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT72), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n531_), .A2(KEYINPUT72), .A3(new_n533_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT73), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n497_), .A2(new_n450_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT12), .ZN(new_n542_));
  INV_X1    g341(.A(new_n450_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n487_), .A2(new_n496_), .A3(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(G230gat), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n544_), .B1(new_n545_), .B2(new_n296_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT65), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n546_), .A2(new_n547_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n542_), .A2(new_n548_), .A3(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n541_), .A2(new_n544_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n551_), .A2(G230gat), .A3(G233gat), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G176gat), .B(G204gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(G148gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(KEYINPUT66), .B(KEYINPUT5), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  XOR2_X1   g356(.A(KEYINPUT67), .B(G120gat), .Z(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n553_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n553_), .A2(new_n559_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(KEYINPUT13), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n560_), .A2(new_n561_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT13), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  AND2_X1   g365(.A1(new_n563_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n540_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n518_), .A2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT101), .ZN(new_n571_));
  NOR3_X1   g370(.A1(new_n571_), .A2(G1gat), .A3(new_n435_), .ZN(new_n572_));
  OR2_X1    g371(.A1(new_n572_), .A2(KEYINPUT38), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(KEYINPUT38), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n442_), .A2(new_n473_), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n513_), .B(KEYINPUT102), .Z(new_n576_));
  INV_X1    g375(.A(new_n538_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n568_), .A2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n575_), .A2(new_n576_), .A3(new_n578_), .ZN(new_n579_));
  OAI21_X1  g378(.A(G1gat), .B1(new_n579_), .B2(new_n435_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n573_), .A2(new_n574_), .A3(new_n580_), .ZN(G1324gat));
  INV_X1    g380(.A(new_n429_), .ZN(new_n582_));
  OAI21_X1  g381(.A(G8gat), .B1(new_n579_), .B2(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT39), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n429_), .A2(new_n453_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n584_), .B1(new_n571_), .B2(new_n585_), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n586_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g386(.A(G15gat), .B1(new_n579_), .B2(new_n248_), .ZN(new_n588_));
  XOR2_X1   g387(.A(new_n588_), .B(KEYINPUT41), .Z(new_n589_));
  OR2_X1    g388(.A1(new_n248_), .A2(G15gat), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n589_), .B1(new_n571_), .B2(new_n590_), .ZN(G1326gat));
  XOR2_X1   g390(.A(new_n319_), .B(KEYINPUT103), .Z(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(G22gat), .B1(new_n579_), .B2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT42), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n593_), .A2(G22gat), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n595_), .B1(new_n571_), .B2(new_n596_), .ZN(G1327gat));
  NAND2_X1  g396(.A1(new_n578_), .A2(new_n473_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n441_), .A2(new_n517_), .ZN(new_n599_));
  OAI21_X1  g398(.A(KEYINPUT104), .B1(new_n514_), .B2(new_n516_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(KEYINPUT43), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n599_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n441_), .A2(new_n517_), .A3(new_n601_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n598_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(KEYINPUT105), .B(KEYINPUT44), .ZN(new_n606_));
  OAI21_X1  g405(.A(KEYINPUT106), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  NOR3_X1   g406(.A1(new_n568_), .A2(new_n577_), .A3(new_n472_), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n441_), .A2(new_n517_), .A3(new_n601_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n601_), .B1(new_n441_), .B2(new_n517_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n608_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT106), .ZN(new_n612_));
  INV_X1    g411(.A(new_n606_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n611_), .A2(new_n612_), .A3(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n607_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n605_), .A2(KEYINPUT44), .ZN(new_n616_));
  AND3_X1   g415(.A1(new_n615_), .A2(new_n362_), .A3(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(G29gat), .ZN(new_n618_));
  INV_X1    g417(.A(new_n513_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n442_), .A2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n620_), .A2(new_n569_), .A3(new_n473_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n362_), .A2(new_n618_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT107), .ZN(new_n623_));
  OAI22_X1  g422(.A1(new_n617_), .A2(new_n618_), .B1(new_n621_), .B2(new_n623_), .ZN(G1328gat));
  NOR3_X1   g423(.A1(new_n621_), .A2(G36gat), .A3(new_n582_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT45), .Z(new_n626_));
  INV_X1    g425(.A(G36gat), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n582_), .B1(new_n605_), .B2(KEYINPUT44), .ZN(new_n628_));
  AOI211_X1 g427(.A(KEYINPUT108), .B(new_n627_), .C1(new_n615_), .C2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT108), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n611_), .A2(new_n612_), .A3(new_n613_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n612_), .B1(new_n611_), .B2(new_n613_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n628_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n630_), .B1(new_n633_), .B2(G36gat), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n626_), .B1(new_n629_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT46), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  OAI211_X1 g436(.A(KEYINPUT46), .B(new_n626_), .C1(new_n629_), .C2(new_n634_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(G1329gat));
  NAND4_X1  g438(.A1(new_n615_), .A2(G43gat), .A3(new_n434_), .A4(new_n616_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(KEYINPUT109), .B(G43gat), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n641_), .B1(new_n621_), .B2(new_n248_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g443(.A(new_n430_), .B1(new_n607_), .B2(new_n614_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n477_), .B1(new_n605_), .B2(KEYINPUT44), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n621_), .A2(new_n593_), .ZN(new_n647_));
  AOI22_X1  g446(.A1(new_n645_), .A2(new_n646_), .B1(new_n477_), .B2(new_n647_), .ZN(G1331gat));
  NAND4_X1  g447(.A1(new_n575_), .A2(new_n576_), .A3(new_n568_), .A4(new_n540_), .ZN(new_n649_));
  INV_X1    g448(.A(G57gat), .ZN(new_n650_));
  NOR3_X1   g449(.A1(new_n649_), .A2(new_n650_), .A3(new_n435_), .ZN(new_n651_));
  XOR2_X1   g450(.A(new_n651_), .B(KEYINPUT110), .Z(new_n652_));
  NOR2_X1   g451(.A1(new_n567_), .A2(new_n538_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n518_), .A2(new_n653_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n650_), .B1(new_n654_), .B2(new_n435_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n652_), .A2(new_n655_), .ZN(G1332gat));
  OAI21_X1  g455(.A(G64gat), .B1(new_n649_), .B2(new_n582_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT48), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n582_), .A2(G64gat), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n658_), .B1(new_n654_), .B2(new_n659_), .ZN(G1333gat));
  OAI21_X1  g459(.A(G71gat), .B1(new_n649_), .B2(new_n248_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT49), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n248_), .A2(G71gat), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n662_), .B1(new_n654_), .B2(new_n663_), .ZN(G1334gat));
  OAI21_X1  g463(.A(G78gat), .B1(new_n649_), .B2(new_n593_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT50), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n593_), .A2(G78gat), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT111), .Z(new_n668_));
  OAI21_X1  g467(.A(new_n666_), .B1(new_n654_), .B2(new_n668_), .ZN(G1335gat));
  NAND3_X1  g468(.A1(new_n620_), .A2(new_n473_), .A3(new_n653_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(G85gat), .B1(new_n671_), .B2(new_n362_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT112), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n653_), .A2(new_n473_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n674_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n494_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n435_), .B1(new_n676_), .B2(new_n492_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n673_), .B1(new_n675_), .B2(new_n677_), .ZN(G1336gat));
  AOI21_X1  g477(.A(G92gat), .B1(new_n671_), .B2(new_n429_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n429_), .A2(G92gat), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n679_), .B1(new_n675_), .B2(new_n680_), .ZN(G1337gat));
  NAND2_X1  g480(.A1(new_n675_), .A2(new_n434_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(G99gat), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT113), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n671_), .A2(new_n488_), .A3(new_n434_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n683_), .A2(new_n684_), .A3(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g486(.A1(new_n671_), .A2(new_n489_), .A3(new_n319_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT52), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n675_), .A2(new_n319_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n689_), .B1(new_n690_), .B2(G106gat), .ZN(new_n691_));
  AOI211_X1 g490(.A(KEYINPUT52), .B(new_n489_), .C1(new_n675_), .C2(new_n319_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n688_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g493(.A(new_n540_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT57), .ZN(new_n696_));
  INV_X1    g495(.A(new_n519_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(new_n520_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n524_), .B(KEYINPUT115), .Z(new_n699_));
  OAI21_X1  g498(.A(new_n698_), .B1(new_n699_), .B2(new_n520_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n533_), .B1(new_n700_), .B2(new_n532_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n562_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT55), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n550_), .A2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n542_), .A2(new_n544_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n705_), .A2(G230gat), .A3(G233gat), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n550_), .A2(new_n703_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n704_), .A2(new_n706_), .A3(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(new_n559_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT56), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n560_), .A2(KEYINPUT114), .A3(new_n710_), .ZN(new_n711_));
  AOI22_X1  g510(.A1(new_n536_), .A2(new_n537_), .B1(new_n709_), .B2(new_n711_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n708_), .A2(new_n559_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n713_), .A2(KEYINPUT114), .A3(new_n710_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n702_), .B1(new_n712_), .B2(new_n714_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n696_), .B1(new_n715_), .B2(new_n513_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n709_), .A2(new_n711_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n538_), .A2(new_n714_), .A3(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n702_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n720_), .A2(KEYINPUT57), .A3(new_n619_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n560_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n722_), .B1(new_n713_), .B2(new_n710_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n701_), .B1(new_n709_), .B2(KEYINPUT56), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(KEYINPUT116), .A2(KEYINPUT58), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n723_), .B(new_n724_), .C1(KEYINPUT116), .C2(KEYINPUT58), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n727_), .A2(new_n517_), .A3(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n716_), .A2(new_n721_), .A3(new_n729_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n517_), .A2(new_n473_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n540_), .A2(new_n731_), .A3(new_n567_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(KEYINPUT54), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT54), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n540_), .A2(new_n731_), .A3(new_n734_), .A4(new_n567_), .ZN(new_n735_));
  AOI22_X1  g534(.A1(new_n730_), .A2(new_n473_), .B1(new_n733_), .B2(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n434_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT117), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(KEYINPUT59), .ZN(new_n739_));
  NOR4_X1   g538(.A1(new_n736_), .A2(new_n435_), .A3(new_n737_), .A4(new_n739_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(KEYINPUT117), .B(KEYINPUT59), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n730_), .A2(new_n473_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n733_), .A2(new_n735_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n737_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n742_), .B1(new_n745_), .B2(new_n362_), .ZN(new_n746_));
  OAI211_X1 g545(.A(G113gat), .B(new_n695_), .C1(new_n740_), .C2(new_n746_), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n736_), .A2(new_n435_), .A3(new_n737_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(new_n538_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(new_n232_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n747_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT118), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n747_), .A2(KEYINPUT118), .A3(new_n750_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(G1340gat));
  INV_X1    g554(.A(G120gat), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n756_), .B1(new_n567_), .B2(KEYINPUT60), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n748_), .B(new_n757_), .C1(KEYINPUT60), .C2(new_n756_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n740_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n746_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n567_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n758_), .B1(new_n761_), .B2(new_n756_), .ZN(G1341gat));
  AOI21_X1  g561(.A(G127gat), .B1(new_n748_), .B2(new_n472_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n759_), .A2(new_n760_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n472_), .A2(G127gat), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT119), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n763_), .B1(new_n764_), .B2(new_n766_), .ZN(G1342gat));
  INV_X1    g566(.A(new_n576_), .ZN(new_n768_));
  AOI21_X1  g567(.A(G134gat), .B1(new_n748_), .B2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n517_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n770_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n769_), .B1(new_n771_), .B2(G134gat), .ZN(G1343gat));
  NAND2_X1  g571(.A1(new_n743_), .A2(new_n744_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n429_), .A2(new_n430_), .ZN(new_n774_));
  AND3_X1   g573(.A1(new_n773_), .A2(new_n248_), .A3(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n362_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n776_), .A2(new_n577_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(new_n256_), .ZN(G1344gat));
  NOR2_X1   g577(.A1(new_n776_), .A2(new_n567_), .ZN(new_n779_));
  XOR2_X1   g578(.A(KEYINPUT120), .B(G148gat), .Z(new_n780_));
  XNOR2_X1  g579(.A(new_n779_), .B(new_n780_), .ZN(G1345gat));
  NOR2_X1   g580(.A1(new_n776_), .A2(new_n473_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(G155gat), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n782_), .B(new_n784_), .ZN(G1346gat));
  NOR2_X1   g584(.A1(new_n736_), .A2(new_n434_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n786_), .A2(new_n362_), .A3(new_n774_), .A4(new_n517_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(G162gat), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT122), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n775_), .A2(new_n262_), .A3(new_n362_), .A4(new_n768_), .ZN(new_n790_));
  AND3_X1   g589(.A1(new_n788_), .A2(new_n789_), .A3(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n789_), .B1(new_n788_), .B2(new_n790_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n791_), .A2(new_n792_), .ZN(G1347gat));
  NAND2_X1  g592(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n582_), .A2(new_n362_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n434_), .A2(new_n795_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT123), .ZN(new_n797_));
  NOR3_X1   g596(.A1(new_n736_), .A2(new_n592_), .A3(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  OAI211_X1 g598(.A(G169gat), .B(new_n794_), .C1(new_n799_), .C2(new_n577_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n801_));
  OR2_X1    g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n798_), .A2(new_n538_), .A3(new_n225_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n800_), .A2(new_n801_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n802_), .A2(new_n803_), .A3(new_n804_), .ZN(G1348gat));
  NAND3_X1  g604(.A1(new_n798_), .A2(new_n203_), .A3(new_n568_), .ZN(new_n806_));
  NOR4_X1   g605(.A1(new_n736_), .A2(new_n567_), .A3(new_n319_), .A4(new_n797_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n806_), .B1(new_n807_), .B2(new_n203_), .ZN(G1349gat));
  NOR3_X1   g607(.A1(new_n799_), .A2(new_n209_), .A3(new_n473_), .ZN(new_n809_));
  OR4_X1    g608(.A1(new_n319_), .A2(new_n736_), .A3(new_n473_), .A4(new_n797_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n809_), .B1(new_n213_), .B2(new_n810_), .ZN(G1350gat));
  OAI21_X1  g610(.A(G190gat), .B1(new_n799_), .B2(new_n770_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n768_), .A2(new_n210_), .ZN(new_n813_));
  XOR2_X1   g612(.A(new_n813_), .B(KEYINPUT125), .Z(new_n814_));
  OAI21_X1  g613(.A(new_n812_), .B1(new_n799_), .B2(new_n814_), .ZN(G1351gat));
  NAND4_X1  g614(.A1(new_n786_), .A2(KEYINPUT126), .A3(new_n319_), .A4(new_n795_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n773_), .A2(new_n248_), .A3(new_n319_), .A4(new_n795_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT126), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n577_), .B1(new_n816_), .B2(new_n819_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n820_), .B(new_n282_), .ZN(G1352gat));
  INV_X1    g620(.A(KEYINPUT127), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(G204gat), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n567_), .B1(new_n816_), .B2(new_n819_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n822_), .A2(G204gat), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n823_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(new_n824_), .B2(new_n823_), .ZN(G1353gat));
  XNOR2_X1  g626(.A(KEYINPUT63), .B(G211gat), .ZN(new_n828_));
  AOI211_X1 g627(.A(new_n473_), .B(new_n828_), .C1(new_n816_), .C2(new_n819_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n816_), .A2(new_n819_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n472_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n829_), .B1(new_n831_), .B2(new_n832_), .ZN(G1354gat));
  AOI21_X1  g632(.A(G218gat), .B1(new_n830_), .B2(new_n768_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n770_), .B1(new_n816_), .B2(new_n819_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n834_), .B1(G218gat), .B2(new_n835_), .ZN(G1355gat));
endmodule


