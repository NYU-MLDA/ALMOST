//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0 0 0 1 0 1 1 0 1 0 0 1 1 1 0 1 1 0 0 0 1 1 1 0 1 0 1 1 0 1 0 0 0 0 0 0 0 0 1 1 0 0 1 1 1 0 0 1 0 1 0 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n742_,
    new_n743_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n872_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n879_, new_n880_, new_n882_, new_n883_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_, new_n902_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n910_, new_n911_, new_n913_,
    new_n914_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_;
  INV_X1    g000(.A(KEYINPUT20), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G183gat), .A2(G190gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT81), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n203_), .A2(KEYINPUT23), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n209_), .B1(G183gat), .B2(G190gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT22), .B(G169gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT92), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(G176gat), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n212_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n210_), .A2(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n205_), .A2(new_n206_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n203_), .A2(KEYINPUT23), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(KEYINPUT82), .ZN(new_n221_));
  OR2_X1    g020(.A1(new_n219_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(G169gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(new_n216_), .ZN(new_n224_));
  OR2_X1    g023(.A1(new_n224_), .A2(KEYINPUT24), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(KEYINPUT24), .A3(new_n211_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT25), .B(G183gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT26), .B(G190gat), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n227_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n222_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n218_), .A2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G211gat), .B(G218gat), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT88), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(G197gat), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT87), .B1(new_n236_), .B2(G204gat), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT87), .ZN(new_n238_));
  INV_X1    g037(.A(G204gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n238_), .A2(new_n239_), .A3(G197gat), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n237_), .B(new_n240_), .C1(G197gat), .C2(new_n239_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n233_), .A2(new_n234_), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n235_), .A2(KEYINPUT21), .A3(new_n241_), .A4(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n236_), .A2(G204gat), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n239_), .A2(G197gat), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT21), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  OAI211_X1 g045(.A(new_n246_), .B(new_n233_), .C1(new_n241_), .C2(KEYINPUT21), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n243_), .A2(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n202_), .B1(new_n232_), .B2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G226gat), .A2(G233gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT19), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT91), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(G183gat), .ZN(new_n254_));
  OAI21_X1  g053(.A(KEYINPUT79), .B1(new_n254_), .B2(KEYINPUT25), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n229_), .B(new_n255_), .C1(new_n228_), .C2(KEYINPUT79), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT80), .ZN(new_n257_));
  AND2_X1   g056(.A1(new_n225_), .A2(new_n226_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n257_), .A2(new_n209_), .A3(new_n258_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(G169gat), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n219_), .A2(new_n221_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(G183gat), .A2(G190gat), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n261_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n259_), .A2(new_n264_), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n249_), .B(new_n253_), .C1(new_n248_), .C2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n248_), .ZN(new_n267_));
  AOI22_X1  g066(.A1(new_n210_), .A2(new_n217_), .B1(new_n222_), .B2(new_n230_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n248_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  AND3_X1   g069(.A1(new_n267_), .A2(KEYINPUT20), .A3(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n251_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n266_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G8gat), .B(G36gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT18), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G64gat), .B(G92gat), .ZN(new_n276_));
  XOR2_X1   g075(.A(new_n275_), .B(new_n276_), .Z(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n273_), .A2(new_n278_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n265_), .A2(new_n248_), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT20), .B1(new_n268_), .B2(new_n269_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n252_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n267_), .A2(KEYINPUT20), .A3(new_n272_), .A4(new_n270_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT97), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n282_), .A2(new_n283_), .A3(new_n284_), .A4(new_n277_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n282_), .A2(new_n277_), .A3(new_n283_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT97), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n279_), .A2(new_n285_), .A3(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT27), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT93), .ZN(new_n290_));
  OR2_X1    g089(.A1(new_n286_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT27), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n282_), .A2(new_n283_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(new_n278_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n286_), .A2(new_n290_), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n291_), .A2(new_n292_), .A3(new_n294_), .A4(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n289_), .A2(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(G141gat), .A2(G148gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT3), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G141gat), .A2(G148gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT2), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G155gat), .A2(G162gat), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(G155gat), .A2(G162gat), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n305_), .B1(KEYINPUT1), .B2(new_n303_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n307_), .B1(KEYINPUT1), .B2(new_n303_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n298_), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n309_), .A2(new_n300_), .ZN(new_n310_));
  AOI22_X1  g109(.A1(new_n302_), .A2(new_n306_), .B1(new_n308_), .B2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT29), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  XOR2_X1   g112(.A(G22gat), .B(G50gat), .Z(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT28), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n313_), .B(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G78gat), .B(G106gat), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G228gat), .A2(G233gat), .ZN(new_n319_));
  OAI211_X1 g118(.A(new_n248_), .B(new_n319_), .C1(new_n312_), .C2(new_n311_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n302_), .A2(new_n306_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n308_), .A2(new_n310_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(KEYINPUT89), .B(KEYINPUT29), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n269_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n318_), .B(new_n320_), .C1(new_n325_), .C2(new_n319_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n316_), .B1(new_n327_), .B2(KEYINPUT90), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n320_), .B1(new_n325_), .B2(new_n319_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(new_n317_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(new_n326_), .ZN(new_n331_));
  OR2_X1    g130(.A1(new_n328_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n328_), .A2(new_n331_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G71gat), .B(G99gat), .ZN(new_n335_));
  INV_X1    g134(.A(G43gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT30), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n265_), .A2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT83), .B(G15gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G227gat), .A2(G233gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n338_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n344_), .A2(new_n259_), .A3(new_n264_), .ZN(new_n345_));
  AND3_X1   g144(.A1(new_n339_), .A2(new_n343_), .A3(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n343_), .B1(new_n339_), .B2(new_n345_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G127gat), .B(G134gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G113gat), .B(G120gat), .ZN(new_n349_));
  XOR2_X1   g148(.A(new_n348_), .B(new_n349_), .Z(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT84), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n348_), .B(new_n349_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT84), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n351_), .A2(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT31), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(KEYINPUT85), .ZN(new_n357_));
  OR3_X1    g156(.A1(new_n346_), .A2(new_n347_), .A3(new_n357_), .ZN(new_n358_));
  OR2_X1    g157(.A1(new_n356_), .A2(KEYINPUT85), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n359_), .B(new_n357_), .C1(new_n346_), .C2(new_n347_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n355_), .A2(new_n323_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n323_), .A2(new_n350_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n362_), .A2(new_n364_), .A3(KEYINPUT4), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G225gat), .A2(G233gat), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n311_), .B1(new_n351_), .B2(new_n354_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(KEYINPUT94), .B(KEYINPUT4), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n365_), .A2(new_n367_), .A3(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n362_), .A2(new_n364_), .A3(new_n366_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G1gat), .B(G29gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(G85gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT0), .B(G57gat), .ZN(new_n376_));
  XOR2_X1   g175(.A(new_n375_), .B(new_n376_), .Z(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n373_), .A2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n371_), .A2(new_n377_), .A3(new_n372_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n361_), .A2(new_n381_), .ZN(new_n382_));
  AND3_X1   g181(.A1(new_n297_), .A2(new_n334_), .A3(new_n382_), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n277_), .A2(KEYINPUT32), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n273_), .A2(new_n384_), .ZN(new_n385_));
  OAI211_X1 g184(.A(new_n385_), .B(new_n381_), .C1(new_n384_), .C2(new_n293_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n380_), .B(KEYINPUT33), .ZN(new_n387_));
  NOR3_X1   g186(.A1(new_n368_), .A2(new_n363_), .A3(new_n366_), .ZN(new_n388_));
  OAI21_X1  g187(.A(KEYINPUT95), .B1(new_n388_), .B2(new_n377_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n362_), .A2(new_n364_), .A3(new_n367_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT95), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n390_), .A2(new_n391_), .A3(new_n378_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n365_), .A2(new_n366_), .A3(new_n370_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n389_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(KEYINPUT96), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT96), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n392_), .A2(new_n389_), .A3(new_n393_), .A4(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n395_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n387_), .A2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n291_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n386_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(new_n334_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n381_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n403_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n297_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n402_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT86), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n361_), .B(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n383_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G43gat), .B(G50gat), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(G36gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(G29gat), .ZN(new_n414_));
  INV_X1    g213(.A(G29gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(G36gat), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n414_), .A2(new_n416_), .A3(KEYINPUT67), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(KEYINPUT67), .B1(new_n414_), .B2(new_n416_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n412_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n414_), .A2(new_n416_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT67), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n423_), .A2(new_n417_), .A3(new_n411_), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n420_), .A2(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G15gat), .B(G22gat), .ZN(new_n426_));
  INV_X1    g225(.A(G1gat), .ZN(new_n427_));
  INV_X1    g226(.A(G8gat), .ZN(new_n428_));
  OAI21_X1  g227(.A(KEYINPUT14), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n426_), .A2(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G1gat), .B(G8gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n430_), .B(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n425_), .B(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G229gat), .A2(G233gat), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  AND3_X1   g235(.A1(new_n420_), .A2(new_n424_), .A3(KEYINPUT15), .ZN(new_n437_));
  AOI21_X1  g236(.A(KEYINPUT15), .B1(new_n420_), .B2(new_n424_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(new_n432_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n425_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n432_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n440_), .A2(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n436_), .B1(new_n444_), .B2(new_n435_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT77), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G113gat), .B(G141gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G169gat), .B(G197gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n447_), .B(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(KEYINPUT75), .B(KEYINPUT76), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n449_), .B(new_n450_), .ZN(new_n451_));
  XOR2_X1   g250(.A(new_n451_), .B(KEYINPUT78), .Z(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n446_), .A2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n445_), .A2(KEYINPUT77), .A3(new_n452_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n410_), .A2(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G57gat), .B(G64gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G71gat), .B(G78gat), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n458_), .A2(new_n459_), .A3(KEYINPUT11), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n458_), .A2(KEYINPUT11), .ZN(new_n461_));
  INV_X1    g260(.A(new_n459_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n458_), .A2(KEYINPUT11), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n460_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  AND2_X1   g264(.A1(G231gat), .A2(G233gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n465_), .B(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(KEYINPUT72), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(new_n432_), .ZN(new_n469_));
  XOR2_X1   g268(.A(G127gat), .B(G155gat), .Z(new_n470_));
  XNOR2_X1  g269(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n470_), .B(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G183gat), .B(G211gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n474_), .A2(KEYINPUT17), .ZN(new_n475_));
  AND2_X1   g274(.A1(new_n469_), .A2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n474_), .B(KEYINPUT17), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n469_), .A2(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT74), .B1(new_n476_), .B2(new_n478_), .ZN(new_n479_));
  OR2_X1    g278(.A1(new_n478_), .A2(KEYINPUT74), .ZN(new_n480_));
  AND2_X1   g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(G85gat), .ZN(new_n483_));
  INV_X1    g282(.A(G92gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G85gat), .A2(G92gat), .ZN(new_n486_));
  AND2_X1   g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G99gat), .A2(G106gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT6), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT6), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n490_), .A2(G99gat), .A3(G106gat), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n489_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT7), .ZN(new_n493_));
  INV_X1    g292(.A(G99gat), .ZN(new_n494_));
  INV_X1    g293(.A(G106gat), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n493_), .A2(new_n494_), .A3(new_n495_), .A4(KEYINPUT65), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT65), .ZN(new_n497_));
  OAI22_X1  g296(.A1(new_n497_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n487_), .B1(new_n492_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT8), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  OAI211_X1 g301(.A(KEYINPUT8), .B(new_n487_), .C1(new_n492_), .C2(new_n499_), .ZN(new_n503_));
  OR2_X1    g302(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n504_), .A2(new_n495_), .A3(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n485_), .A2(KEYINPUT9), .A3(new_n486_), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n486_), .A2(KEYINPUT9), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n509_), .B1(new_n489_), .B2(new_n491_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n502_), .A2(new_n503_), .A3(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT66), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  AOI22_X1  g313(.A1(new_n500_), .A2(new_n501_), .B1(new_n508_), .B2(new_n510_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n515_), .A2(KEYINPUT66), .A3(new_n503_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n514_), .A2(new_n439_), .A3(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G232gat), .A2(G233gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT34), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n519_), .A2(KEYINPUT35), .ZN(new_n520_));
  AND3_X1   g319(.A1(new_n502_), .A2(new_n503_), .A3(new_n511_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n520_), .B1(new_n521_), .B2(new_n441_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n517_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n519_), .A2(KEYINPUT35), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n524_), .A2(KEYINPUT68), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n524_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT68), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n523_), .A2(new_n526_), .A3(new_n530_), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n517_), .A2(new_n522_), .A3(new_n528_), .A4(new_n527_), .ZN(new_n532_));
  XOR2_X1   g331(.A(G190gat), .B(G218gat), .Z(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT69), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G134gat), .B(G162gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  XOR2_X1   g335(.A(new_n536_), .B(KEYINPUT36), .Z(new_n537_));
  NAND3_X1  g336(.A1(new_n531_), .A2(new_n532_), .A3(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT71), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT71), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n531_), .A2(new_n532_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n536_), .A2(KEYINPUT36), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(new_n538_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n540_), .B1(new_n541_), .B2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT37), .ZN(new_n547_));
  AND3_X1   g346(.A1(new_n531_), .A2(new_n532_), .A3(new_n537_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n543_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n549_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n550_));
  OAI21_X1  g349(.A(KEYINPUT37), .B1(new_n548_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT70), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n545_), .A2(KEYINPUT70), .A3(KEYINPUT37), .ZN(new_n554_));
  AOI22_X1  g353(.A1(new_n546_), .A2(new_n547_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n482_), .A2(new_n555_), .ZN(new_n556_));
  OAI211_X1 g355(.A(KEYINPUT12), .B(new_n460_), .C1(new_n463_), .C2(new_n464_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n514_), .A2(new_n516_), .A3(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT12), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n560_), .B1(new_n521_), .B2(new_n465_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G230gat), .A2(G233gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT64), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n515_), .A2(new_n503_), .A3(new_n465_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n559_), .A2(new_n561_), .A3(new_n564_), .A4(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n565_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n465_), .B1(new_n515_), .B2(new_n503_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n563_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n566_), .A2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G120gat), .B(G148gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT5), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G176gat), .B(G204gat), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n572_), .B(new_n573_), .Z(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n570_), .A2(new_n575_), .ZN(new_n576_));
  AND3_X1   g375(.A1(new_n566_), .A2(new_n569_), .A3(new_n575_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT13), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n457_), .A2(new_n556_), .A3(new_n580_), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n381_), .A2(KEYINPUT98), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n381_), .A2(KEYINPUT98), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n581_), .A2(new_n427_), .A3(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT38), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT100), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n410_), .A2(new_n546_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n456_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n580_), .A2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT99), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n591_), .A2(new_n481_), .A3(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(G1gat), .B1(new_n595_), .B2(new_n403_), .ZN(new_n596_));
  OAI211_X1 g395(.A(new_n590_), .B(new_n596_), .C1(new_n587_), .C2(new_n586_), .ZN(G1324gat));
  INV_X1    g396(.A(new_n297_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n581_), .A2(new_n428_), .A3(new_n598_), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n595_), .A2(new_n297_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT39), .ZN(new_n601_));
  AND3_X1   g400(.A1(new_n600_), .A2(new_n601_), .A3(G8gat), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n601_), .B1(new_n600_), .B2(G8gat), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n599_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT40), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  OAI211_X1 g405(.A(KEYINPUT40), .B(new_n599_), .C1(new_n602_), .C2(new_n603_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(G1325gat));
  OAI21_X1  g407(.A(G15gat), .B1(new_n595_), .B2(new_n409_), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n609_), .B(KEYINPUT101), .Z(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(KEYINPUT41), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n609_), .B(KEYINPUT101), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT41), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(G15gat), .ZN(new_n615_));
  INV_X1    g414(.A(new_n409_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n581_), .A2(new_n615_), .A3(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n611_), .A2(new_n614_), .A3(new_n617_), .ZN(G1326gat));
  OAI21_X1  g417(.A(G22gat), .B1(new_n595_), .B2(new_n334_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT42), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n334_), .A2(G22gat), .ZN(new_n621_));
  XOR2_X1   g420(.A(new_n621_), .B(KEYINPUT102), .Z(new_n622_));
  NAND2_X1  g421(.A1(new_n581_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n620_), .A2(new_n623_), .ZN(G1327gat));
  NAND2_X1  g423(.A1(new_n482_), .A2(new_n546_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n580_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n457_), .A2(new_n415_), .A3(new_n381_), .A4(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT104), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n594_), .A2(new_n482_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n555_), .A2(KEYINPUT103), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(KEYINPUT43), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n541_), .B1(new_n548_), .B2(new_n550_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n634_), .A2(new_n547_), .A3(new_n539_), .ZN(new_n635_));
  AOI21_X1  g434(.A(KEYINPUT70), .B1(new_n545_), .B2(KEYINPUT37), .ZN(new_n636_));
  AOI211_X1 g435(.A(new_n552_), .B(new_n547_), .C1(new_n544_), .C2(new_n538_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n635_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n633_), .B1(new_n410_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n334_), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n295_), .A2(new_n294_), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n641_), .A2(new_n291_), .A3(new_n398_), .A4(new_n387_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n640_), .B1(new_n642_), .B2(new_n386_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n404_), .B1(new_n289_), .B2(new_n296_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n409_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n297_), .A2(new_n334_), .A3(new_n382_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n647_), .A2(new_n555_), .A3(new_n632_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n630_), .B1(new_n639_), .B2(new_n648_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n629_), .B1(new_n649_), .B2(KEYINPUT44), .ZN(new_n650_));
  INV_X1    g449(.A(new_n630_), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n647_), .A2(new_n555_), .A3(new_n632_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n632_), .B1(new_n647_), .B2(new_n555_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n651_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT44), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n654_), .A2(KEYINPUT104), .A3(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n650_), .A2(new_n656_), .ZN(new_n657_));
  OAI211_X1 g456(.A(KEYINPUT44), .B(new_n651_), .C1(new_n652_), .C2(new_n653_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(new_n585_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n657_), .A2(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(KEYINPUT105), .B1(new_n661_), .B2(G29gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n659_), .B1(new_n650_), .B2(new_n656_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT105), .ZN(new_n664_));
  NOR3_X1   g463(.A1(new_n663_), .A2(new_n664_), .A3(new_n415_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n628_), .B1(new_n662_), .B2(new_n665_), .ZN(G1328gat));
  INV_X1    g465(.A(KEYINPUT46), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n658_), .A2(new_n598_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n413_), .B1(new_n657_), .B2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n457_), .A2(new_n627_), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n297_), .A2(KEYINPUT106), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n297_), .A2(KEYINPUT106), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n671_), .A2(G36gat), .A3(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT45), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n667_), .B1(new_n670_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT45), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n676_), .B(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n668_), .B1(new_n650_), .B2(new_n656_), .ZN(new_n681_));
  OAI211_X1 g480(.A(new_n680_), .B(KEYINPUT46), .C1(new_n413_), .C2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n678_), .A2(new_n682_), .ZN(G1329gat));
  NAND3_X1  g482(.A1(new_n358_), .A2(G43gat), .A3(new_n360_), .ZN(new_n684_));
  AOI211_X1 g483(.A(new_n655_), .B(new_n630_), .C1(new_n639_), .C2(new_n648_), .ZN(new_n685_));
  AOI211_X1 g484(.A(new_n684_), .B(new_n685_), .C1(new_n650_), .C2(new_n656_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n336_), .B1(new_n671_), .B2(new_n409_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(KEYINPUT47), .B1(new_n686_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT47), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n657_), .A2(new_n658_), .ZN(new_n691_));
  OAI211_X1 g490(.A(new_n690_), .B(new_n687_), .C1(new_n691_), .C2(new_n684_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n689_), .A2(new_n692_), .ZN(G1330gat));
  INV_X1    g492(.A(KEYINPUT107), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n640_), .A2(G50gat), .ZN(new_n695_));
  AOI211_X1 g494(.A(new_n695_), .B(new_n685_), .C1(new_n650_), .C2(new_n656_), .ZN(new_n696_));
  INV_X1    g495(.A(G50gat), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n697_), .B1(new_n671_), .B2(new_n334_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n694_), .B1(new_n696_), .B2(new_n699_), .ZN(new_n700_));
  OAI211_X1 g499(.A(KEYINPUT107), .B(new_n698_), .C1(new_n691_), .C2(new_n695_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(G1331gat));
  NOR2_X1   g501(.A1(new_n410_), .A2(new_n592_), .ZN(new_n703_));
  AND3_X1   g502(.A1(new_n703_), .A2(new_n556_), .A3(new_n626_), .ZN(new_n704_));
  AOI21_X1  g503(.A(G57gat), .B1(new_n704_), .B2(new_n585_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT108), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n626_), .A2(new_n456_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n707_), .A2(new_n482_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n591_), .A2(new_n708_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT109), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n381_), .A2(G57gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n706_), .B1(new_n710_), .B2(new_n711_), .ZN(G1332gat));
  INV_X1    g511(.A(G64gat), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n704_), .A2(new_n713_), .A3(new_n674_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n710_), .B2(new_n674_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT48), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n715_), .A2(new_n716_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n714_), .B1(new_n717_), .B2(new_n718_), .ZN(G1333gat));
  INV_X1    g518(.A(G71gat), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n704_), .A2(new_n720_), .A3(new_n616_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n710_), .B2(new_n616_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT49), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n722_), .A2(new_n723_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n721_), .B1(new_n724_), .B2(new_n725_), .ZN(G1334gat));
  INV_X1    g525(.A(G78gat), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n704_), .A2(new_n727_), .A3(new_n640_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n727_), .B1(new_n710_), .B2(new_n640_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n729_), .A2(new_n730_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n728_), .B1(new_n731_), .B2(new_n732_), .ZN(G1335gat));
  NOR2_X1   g532(.A1(new_n707_), .A2(new_n481_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n734_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n735_));
  OAI21_X1  g534(.A(G85gat), .B1(new_n735_), .B2(new_n403_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n625_), .A2(new_n580_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n703_), .A2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n739_), .A2(new_n483_), .A3(new_n585_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n736_), .A2(new_n740_), .ZN(G1336gat));
  OAI21_X1  g540(.A(G92gat), .B1(new_n735_), .B2(new_n675_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n739_), .A2(new_n484_), .A3(new_n598_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(G1337gat));
  NAND2_X1  g543(.A1(new_n504_), .A2(new_n505_), .ZN(new_n745_));
  OR3_X1    g544(.A1(new_n738_), .A2(new_n361_), .A3(new_n745_), .ZN(new_n746_));
  OAI211_X1 g545(.A(new_n616_), .B(new_n734_), .C1(new_n652_), .C2(new_n653_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT111), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n747_), .A2(new_n748_), .A3(G99gat), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n747_), .B2(G99gat), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n746_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT51), .ZN(G1338gat));
  NOR2_X1   g551(.A1(new_n334_), .A2(G106gat), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  OR3_X1    g553(.A1(new_n738_), .A2(KEYINPUT112), .A3(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(KEYINPUT112), .B1(new_n738_), .B2(new_n754_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n640_), .B(new_n734_), .C1(new_n652_), .C2(new_n653_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(G106gat), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT52), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n758_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n757_), .A2(new_n761_), .A3(new_n762_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n763_), .B(new_n764_), .ZN(G1339gat));
  NAND4_X1  g564(.A1(new_n481_), .A2(new_n456_), .A3(new_n638_), .A4(new_n580_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT54), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n766_), .B(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT117), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n514_), .A2(new_n516_), .A3(new_n558_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n565_), .B1(new_n568_), .B2(KEYINPUT12), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n563_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n772_), .A2(KEYINPUT55), .A3(new_n566_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n770_), .A2(new_n771_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT55), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n774_), .A2(new_n775_), .A3(new_n564_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n773_), .A2(new_n776_), .A3(new_n574_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT56), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n575_), .A2(new_n778_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n773_), .A2(new_n776_), .A3(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT115), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT115), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n773_), .A2(new_n776_), .A3(new_n783_), .A4(new_n780_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n779_), .A2(new_n782_), .A3(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n451_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT114), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n444_), .A2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n440_), .A2(KEYINPUT114), .A3(new_n443_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n434_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n433_), .A2(new_n435_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n786_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n577_), .ZN(new_n793_));
  OR2_X1    g592(.A1(new_n445_), .A2(new_n786_), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n792_), .A2(new_n793_), .A3(new_n794_), .ZN(new_n795_));
  AND3_X1   g594(.A1(new_n785_), .A2(KEYINPUT58), .A3(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(KEYINPUT58), .B1(new_n785_), .B2(new_n795_), .ZN(new_n797_));
  NOR3_X1   g596(.A1(new_n796_), .A2(new_n797_), .A3(new_n638_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n634_), .A2(new_n539_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n454_), .A2(new_n793_), .A3(new_n455_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n800_), .B1(new_n779_), .B2(new_n781_), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n792_), .B(new_n794_), .C1(new_n576_), .C2(new_n577_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n799_), .B1(new_n801_), .B2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT57), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n769_), .B1(new_n798_), .B2(new_n806_), .ZN(new_n807_));
  OAI211_X1 g606(.A(KEYINPUT57), .B(new_n799_), .C1(new_n801_), .C2(new_n803_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n785_), .A2(new_n795_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT58), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n785_), .A2(KEYINPUT58), .A3(new_n795_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n811_), .A2(new_n555_), .A3(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n804_), .A2(new_n805_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n813_), .A2(KEYINPUT117), .A3(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n807_), .A2(new_n808_), .A3(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n768_), .B1(new_n816_), .B2(new_n482_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n598_), .A2(new_n640_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n584_), .A2(new_n361_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n820_), .A2(KEYINPUT59), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(KEYINPUT118), .B1(new_n817_), .B2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT118), .ZN(new_n824_));
  INV_X1    g623(.A(new_n808_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n813_), .A2(new_n814_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n825_), .B1(new_n826_), .B2(new_n769_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n481_), .B1(new_n827_), .B2(new_n815_), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n824_), .B(new_n821_), .C1(new_n828_), .C2(new_n768_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n823_), .A2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n813_), .A2(new_n808_), .A3(new_n814_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n813_), .A2(new_n814_), .A3(KEYINPUT116), .A4(new_n808_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n833_), .A2(new_n482_), .A3(new_n834_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n766_), .B(KEYINPUT54), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n820_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(KEYINPUT59), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n830_), .A2(new_n592_), .A3(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(G113gat), .ZN(new_n842_));
  OR2_X1    g641(.A1(new_n456_), .A2(G113gat), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n839_), .B2(new_n843_), .ZN(G1340gat));
  INV_X1    g643(.A(KEYINPUT121), .ZN(new_n845_));
  XNOR2_X1  g644(.A(KEYINPUT119), .B(G120gat), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n580_), .B1(new_n839_), .B2(KEYINPUT59), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n846_), .B1(new_n830_), .B2(new_n847_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n580_), .A2(KEYINPUT60), .ZN(new_n849_));
  MUX2_X1   g648(.A(KEYINPUT60), .B(new_n849_), .S(new_n846_), .Z(new_n850_));
  NAND3_X1  g649(.A1(new_n837_), .A2(new_n838_), .A3(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(KEYINPUT120), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n820_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT120), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(new_n854_), .A3(new_n850_), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n852_), .A2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n845_), .B1(new_n848_), .B2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n852_), .A2(new_n855_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT59), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n626_), .B1(new_n853_), .B2(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n860_), .B1(new_n823_), .B2(new_n829_), .ZN(new_n861_));
  OAI211_X1 g660(.A(KEYINPUT121), .B(new_n858_), .C1(new_n861_), .C2(new_n846_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n857_), .A2(new_n862_), .ZN(G1341gat));
  AOI21_X1  g662(.A(G127gat), .B1(new_n853_), .B2(new_n481_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n830_), .A2(new_n840_), .ZN(new_n865_));
  INV_X1    g664(.A(G127gat), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n866_), .B1(new_n481_), .B2(KEYINPUT122), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n867_), .B1(KEYINPUT122), .B2(new_n866_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n864_), .B1(new_n865_), .B2(new_n868_), .ZN(G1342gat));
  NAND3_X1  g668(.A1(new_n830_), .A2(new_n555_), .A3(new_n840_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(G134gat), .ZN(new_n871_));
  OR2_X1    g670(.A1(new_n799_), .A2(G134gat), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n871_), .B1(new_n839_), .B2(new_n872_), .ZN(G1343gat));
  AOI21_X1  g672(.A(new_n616_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n874_), .A2(new_n640_), .A3(new_n585_), .A4(new_n675_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n875_), .A2(new_n456_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(KEYINPUT123), .B(G141gat), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n876_), .B(new_n877_), .ZN(G1344gat));
  NOR2_X1   g677(.A1(new_n875_), .A2(new_n580_), .ZN(new_n879_));
  XOR2_X1   g678(.A(KEYINPUT124), .B(G148gat), .Z(new_n880_));
  XNOR2_X1  g679(.A(new_n879_), .B(new_n880_), .ZN(G1345gat));
  NOR2_X1   g680(.A1(new_n875_), .A2(new_n482_), .ZN(new_n882_));
  XOR2_X1   g681(.A(KEYINPUT61), .B(G155gat), .Z(new_n883_));
  XNOR2_X1  g682(.A(new_n882_), .B(new_n883_), .ZN(G1346gat));
  OAI21_X1  g683(.A(G162gat), .B1(new_n875_), .B2(new_n638_), .ZN(new_n885_));
  OR2_X1    g684(.A1(new_n799_), .A2(G162gat), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n885_), .B1(new_n875_), .B2(new_n886_), .ZN(G1347gat));
  NOR3_X1   g686(.A1(new_n675_), .A2(new_n409_), .A3(new_n585_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(new_n334_), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n817_), .A2(new_n456_), .A3(new_n889_), .ZN(new_n890_));
  OR3_X1    g689(.A1(new_n890_), .A2(KEYINPUT125), .A3(new_n223_), .ZN(new_n891_));
  OAI21_X1  g690(.A(KEYINPUT125), .B1(new_n890_), .B2(new_n223_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n891_), .A2(KEYINPUT62), .A3(new_n892_), .ZN(new_n893_));
  OR2_X1    g692(.A1(new_n892_), .A2(KEYINPUT62), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n817_), .A2(new_n889_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n592_), .A2(new_n215_), .ZN(new_n896_));
  XOR2_X1   g695(.A(new_n896_), .B(KEYINPUT126), .Z(new_n897_));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n897_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n893_), .A2(new_n894_), .A3(new_n898_), .ZN(G1348gat));
  AOI21_X1  g698(.A(G176gat), .B1(new_n895_), .B2(new_n626_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n640_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n901_));
  AND3_X1   g700(.A1(new_n888_), .A2(G176gat), .A3(new_n626_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n900_), .B1(new_n901_), .B2(new_n902_), .ZN(G1349gat));
  INV_X1    g702(.A(new_n895_), .ZN(new_n904_));
  NOR3_X1   g703(.A1(new_n904_), .A2(new_n228_), .A3(new_n482_), .ZN(new_n905_));
  AND3_X1   g704(.A1(new_n901_), .A2(new_n481_), .A3(new_n888_), .ZN(new_n906_));
  OR2_X1    g705(.A1(new_n906_), .A2(KEYINPUT127), .ZN(new_n907_));
  AOI21_X1  g706(.A(G183gat), .B1(new_n906_), .B2(KEYINPUT127), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n905_), .B1(new_n907_), .B2(new_n908_), .ZN(G1350gat));
  OAI21_X1  g708(.A(G190gat), .B1(new_n904_), .B2(new_n638_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n895_), .A2(new_n229_), .A3(new_n546_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(G1351gat));
  NAND3_X1  g711(.A1(new_n874_), .A2(new_n405_), .A3(new_n674_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n913_), .A2(new_n456_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(new_n236_), .ZN(G1352gat));
  NOR2_X1   g714(.A1(new_n913_), .A2(new_n580_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(new_n239_), .ZN(G1353gat));
  NOR2_X1   g716(.A1(new_n913_), .A2(new_n482_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n919_));
  AND2_X1   g718(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n918_), .B1(new_n919_), .B2(new_n920_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n921_), .B1(new_n918_), .B2(new_n919_), .ZN(G1354gat));
  OAI21_X1  g721(.A(G218gat), .B1(new_n913_), .B2(new_n638_), .ZN(new_n923_));
  OR2_X1    g722(.A1(new_n799_), .A2(G218gat), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n923_), .B1(new_n913_), .B2(new_n924_), .ZN(G1355gat));
endmodule


