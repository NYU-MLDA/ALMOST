//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 1 0 0 0 1 1 1 0 0 0 1 1 0 0 0 1 0 0 1 1 0 0 1 0 0 1 1 1 1 1 0 1 1 1 0 1 0 0 0 0 1 1 0 0 1 1 0 0 0 1 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n801_, new_n802_, new_n803_, new_n804_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n821_, new_n822_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n955_, new_n956_, new_n957_, new_n958_, new_n960_,
    new_n961_, new_n963_, new_n964_, new_n966_, new_n967_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n981_, new_n982_,
    new_n983_, new_n984_, new_n985_, new_n987_, new_n988_, new_n990_,
    new_n991_, new_n993_, new_n994_, new_n996_, new_n997_, new_n998_,
    new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1006_,
    new_n1007_;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G71gat), .B(G78gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n204_), .B1(KEYINPUT11), .B2(new_n202_), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n206_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT6), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  XOR2_X1   g013(.A(KEYINPUT10), .B(G99gat), .Z(new_n215_));
  INV_X1    g014(.A(G106gat), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n214_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(G85gat), .ZN(new_n218_));
  INV_X1    g017(.A(G92gat), .ZN(new_n219_));
  AOI21_X1  g018(.A(KEYINPUT65), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G85gat), .A2(G92gat), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n220_), .B1(new_n222_), .B2(KEYINPUT64), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT9), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT65), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n225_), .B1(G85gat), .B2(G92gat), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n224_), .B1(new_n226_), .B2(new_n221_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n223_), .A2(new_n227_), .ZN(new_n228_));
  OAI211_X1 g027(.A(new_n220_), .B(new_n224_), .C1(new_n222_), .C2(KEYINPUT64), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n217_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT7), .ZN(new_n231_));
  INV_X1    g030(.A(G99gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n231_), .A2(new_n232_), .A3(new_n216_), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n233_), .A2(new_n212_), .A3(new_n213_), .A4(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT66), .ZN(new_n236_));
  NOR2_X1   g035(.A1(G85gat), .A2(G92gat), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n222_), .A2(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n235_), .A2(new_n236_), .A3(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(KEYINPUT8), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n236_), .B1(new_n235_), .B2(new_n238_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n230_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  AOI211_X1 g041(.A(new_n236_), .B(KEYINPUT8), .C1(new_n235_), .C2(new_n238_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n209_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT12), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n243_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n235_), .A2(new_n238_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT66), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n249_), .A2(KEYINPUT8), .A3(new_n239_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n209_), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n247_), .A2(new_n250_), .A3(new_n251_), .A4(new_n230_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n250_), .A2(new_n247_), .A3(new_n230_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n253_), .A2(KEYINPUT12), .A3(new_n209_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G230gat), .A2(G233gat), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n246_), .A2(new_n252_), .A3(new_n254_), .A4(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT67), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NOR3_X1   g057(.A1(new_n242_), .A2(new_n243_), .A3(new_n209_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n259_), .B1(new_n245_), .B2(new_n244_), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n260_), .A2(KEYINPUT67), .A3(new_n255_), .A4(new_n254_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n252_), .A2(new_n244_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n255_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n258_), .A2(new_n261_), .A3(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G120gat), .B(G148gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT5), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT68), .ZN(new_n268_));
  XOR2_X1   g067(.A(G176gat), .B(G204gat), .Z(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(KEYINPUT69), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n268_), .B(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n265_), .A2(new_n272_), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n258_), .A2(new_n261_), .A3(new_n264_), .A4(new_n271_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n273_), .A2(KEYINPUT70), .A3(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT70), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n265_), .A2(new_n276_), .A3(new_n272_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  OR2_X1    g077(.A1(new_n278_), .A2(KEYINPUT13), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(KEYINPUT13), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G29gat), .B(G36gat), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n282_), .A2(KEYINPUT71), .ZN(new_n283_));
  INV_X1    g082(.A(G36gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(G29gat), .ZN(new_n285_));
  INV_X1    g084(.A(G29gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(G36gat), .ZN(new_n287_));
  AND3_X1   g086(.A1(new_n285_), .A2(new_n287_), .A3(KEYINPUT71), .ZN(new_n288_));
  INV_X1    g087(.A(G50gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(G43gat), .ZN(new_n290_));
  INV_X1    g089(.A(G43gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(G50gat), .ZN(new_n292_));
  AND3_X1   g091(.A1(new_n290_), .A2(new_n292_), .A3(KEYINPUT72), .ZN(new_n293_));
  AOI21_X1  g092(.A(KEYINPUT72), .B1(new_n290_), .B2(new_n292_), .ZN(new_n294_));
  OAI22_X1  g093(.A1(new_n283_), .A2(new_n288_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n285_), .A2(new_n287_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT71), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n282_), .A2(KEYINPUT71), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT72), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n291_), .A2(G50gat), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n289_), .A2(G43gat), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n300_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n290_), .A2(new_n292_), .A3(KEYINPUT72), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n298_), .A2(new_n299_), .A3(new_n303_), .A4(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n295_), .A2(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G15gat), .B(G22gat), .ZN(new_n307_));
  INV_X1    g106(.A(G1gat), .ZN(new_n308_));
  INV_X1    g107(.A(G8gat), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT14), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n307_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G1gat), .B(G8gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  XOR2_X1   g112(.A(new_n306_), .B(new_n313_), .Z(new_n314_));
  NAND2_X1  g113(.A1(G229gat), .A2(G233gat), .ZN(new_n315_));
  OR2_X1    g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n313_), .B1(new_n305_), .B2(new_n295_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n306_), .A2(KEYINPUT15), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT15), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n295_), .A2(new_n305_), .A3(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n317_), .B1(new_n321_), .B2(new_n313_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n315_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n316_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G113gat), .B(G141gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G169gat), .B(G197gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n324_), .B(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n330_), .A2(KEYINPUT78), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT78), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n329_), .A2(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n281_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(G169gat), .ZN(new_n336_));
  INV_X1    g135(.A(G176gat), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n336_), .A2(new_n337_), .A3(KEYINPUT81), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT81), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n339_), .B1(G169gat), .B2(G176gat), .ZN(new_n340_));
  AOI21_X1  g139(.A(KEYINPUT24), .B1(new_n338_), .B2(new_n340_), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n338_), .A2(new_n340_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G169gat), .A2(G176gat), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n343_), .A2(KEYINPUT24), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n341_), .B1(new_n342_), .B2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(G190gat), .ZN(new_n346_));
  AOI21_X1  g145(.A(KEYINPUT80), .B1(new_n346_), .B2(KEYINPUT26), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(KEYINPUT26), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT26), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(G190gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n347_), .B1(new_n351_), .B2(KEYINPUT80), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT25), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(G183gat), .ZN(new_n354_));
  INV_X1    g153(.A(G183gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT25), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT79), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n354_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n353_), .A2(KEYINPUT79), .A3(G183gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n352_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT23), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n362_), .A2(G183gat), .A3(G190gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(KEYINPUT82), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G183gat), .A2(G190gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(KEYINPUT23), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT82), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n367_), .A2(new_n362_), .A3(G183gat), .A4(G190gat), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n364_), .A2(new_n366_), .A3(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n345_), .A2(new_n361_), .A3(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n343_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT22), .B(G169gat), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n371_), .B1(new_n372_), .B2(new_n337_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n355_), .A2(KEYINPUT23), .ZN(new_n374_));
  AOI22_X1  g173(.A1(new_n374_), .A2(G190gat), .B1(KEYINPUT23), .B2(new_n365_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(G183gat), .A2(G190gat), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n373_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n370_), .A2(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(KEYINPUT83), .B(KEYINPUT30), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G227gat), .A2(G233gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(G15gat), .ZN(new_n382_));
  XOR2_X1   g181(.A(G71gat), .B(G99gat), .Z(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT84), .B(G43gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n380_), .B(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT85), .ZN(new_n388_));
  OR2_X1    g187(.A1(new_n380_), .A2(new_n386_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT85), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n380_), .A2(new_n386_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n389_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G127gat), .B(G134gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G113gat), .B(G120gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(KEYINPUT31), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n388_), .A2(new_n392_), .A3(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n396_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n387_), .A2(KEYINPUT85), .A3(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  AND3_X1   g200(.A1(KEYINPUT87), .A2(G155gat), .A3(G162gat), .ZN(new_n402_));
  AOI21_X1  g201(.A(KEYINPUT87), .B1(G155gat), .B2(G162gat), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT1), .ZN(new_n404_));
  NOR3_X1   g203(.A1(new_n402_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G155gat), .A2(G162gat), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT87), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(KEYINPUT87), .A2(G155gat), .A3(G162gat), .ZN(new_n409_));
  AOI21_X1  g208(.A(KEYINPUT1), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  OAI22_X1  g209(.A1(new_n405_), .A2(new_n410_), .B1(G155gat), .B2(G162gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G141gat), .A2(G148gat), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(G141gat), .A2(G148gat), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT2), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n416_), .B1(new_n412_), .B2(KEYINPUT88), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n412_), .A2(KEYINPUT88), .A3(new_n416_), .ZN(new_n419_));
  OAI21_X1  g218(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT3), .ZN(new_n421_));
  INV_X1    g220(.A(G141gat), .ZN(new_n422_));
  INV_X1    g221(.A(G148gat), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n421_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n418_), .A2(new_n419_), .A3(new_n420_), .A4(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(G155gat), .ZN(new_n426_));
  INV_X1    g225(.A(G162gat), .ZN(new_n427_));
  AOI22_X1  g226(.A1(new_n408_), .A2(new_n409_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  AOI22_X1  g227(.A1(new_n411_), .A2(new_n415_), .B1(new_n425_), .B2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(new_n395_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n404_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n408_), .A2(KEYINPUT1), .A3(new_n409_), .ZN(new_n432_));
  AOI22_X1  g231(.A1(new_n431_), .A2(new_n432_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n415_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n424_), .A2(new_n420_), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n412_), .A2(KEYINPUT88), .A3(new_n416_), .ZN(new_n436_));
  NOR3_X1   g235(.A1(new_n435_), .A2(new_n436_), .A3(new_n417_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n428_), .ZN(new_n438_));
  OAI22_X1  g237(.A1(new_n433_), .A2(new_n434_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n395_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G225gat), .A2(G233gat), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n430_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n430_), .A2(KEYINPUT4), .A3(new_n441_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n442_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n445_), .B1(new_n441_), .B2(KEYINPUT4), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n443_), .B1(new_n444_), .B2(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G1gat), .B(G29gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(KEYINPUT0), .ZN(new_n449_));
  INV_X1    g248(.A(G57gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n449_), .B(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(new_n218_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n447_), .A2(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n451_), .B(G85gat), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n454_), .B(new_n443_), .C1(new_n444_), .C2(new_n446_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT100), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT29), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n429_), .A2(new_n459_), .ZN(new_n460_));
  XOR2_X1   g259(.A(new_n460_), .B(KEYINPUT28), .Z(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G197gat), .B(G204gat), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT21), .ZN(new_n464_));
  INV_X1    g263(.A(G218gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(G211gat), .ZN(new_n466_));
  INV_X1    g265(.A(G211gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(G218gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n463_), .B1(new_n464_), .B2(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G211gat), .B(G218gat), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT21), .B1(new_n471_), .B2(KEYINPUT90), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(new_n472_), .ZN(new_n473_));
  OAI211_X1 g272(.A(KEYINPUT21), .B(new_n463_), .C1(new_n471_), .C2(KEYINPUT90), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n473_), .A2(KEYINPUT91), .A3(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(KEYINPUT91), .B1(new_n473_), .B2(new_n474_), .ZN(new_n476_));
  OAI22_X1  g275(.A1(new_n475_), .A2(new_n476_), .B1(new_n429_), .B2(new_n459_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G228gat), .A2(G233gat), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT89), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n481_), .B1(new_n429_), .B2(new_n459_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n439_), .A2(KEYINPUT89), .A3(KEYINPUT29), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n479_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n482_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G78gat), .B(G106gat), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  AND3_X1   g286(.A1(new_n480_), .A2(new_n485_), .A3(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n487_), .B1(new_n480_), .B2(new_n485_), .ZN(new_n489_));
  XOR2_X1   g288(.A(G22gat), .B(G50gat), .Z(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NOR3_X1   g290(.A1(new_n488_), .A2(new_n489_), .A3(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n483_), .A2(new_n484_), .ZN(new_n493_));
  AOI21_X1  g292(.A(KEYINPUT89), .B1(new_n439_), .B2(KEYINPUT29), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT91), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT90), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n464_), .B1(new_n469_), .B2(new_n497_), .ZN(new_n498_));
  AND2_X1   g297(.A1(G197gat), .A2(G204gat), .ZN(new_n499_));
  NOR2_X1   g298(.A1(G197gat), .A2(G204gat), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n501_), .B1(new_n471_), .B2(KEYINPUT21), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n498_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n474_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n496_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n473_), .A2(KEYINPUT91), .A3(new_n474_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n439_), .A2(KEYINPUT29), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n478_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n486_), .B1(new_n495_), .B2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n480_), .A2(new_n485_), .A3(new_n487_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n490_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n462_), .B1(new_n492_), .B2(new_n512_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n491_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n510_), .A2(new_n511_), .A3(new_n490_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n514_), .A2(new_n515_), .A3(new_n461_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n513_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT27), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G8gat), .B(G36gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT18), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT96), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G64gat), .B(G92gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n503_), .A2(new_n504_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n525_), .A2(new_n370_), .A3(new_n377_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT20), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT94), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n526_), .A2(KEYINPUT94), .A3(KEYINPUT20), .ZN(new_n530_));
  AND4_X1   g329(.A1(new_n354_), .A2(new_n356_), .A3(new_n348_), .A4(new_n350_), .ZN(new_n531_));
  NOR3_X1   g330(.A1(new_n531_), .A2(new_n341_), .A3(new_n375_), .ZN(new_n532_));
  AND3_X1   g331(.A1(new_n343_), .A2(KEYINPUT95), .A3(KEYINPUT24), .ZN(new_n533_));
  AOI21_X1  g332(.A(KEYINPUT95), .B1(new_n343_), .B2(KEYINPUT24), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n342_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n376_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n369_), .A2(new_n536_), .ZN(new_n537_));
  AOI22_X1  g336(.A1(new_n532_), .A2(new_n535_), .B1(new_n537_), .B2(new_n373_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n538_), .A2(new_n525_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n529_), .A2(new_n530_), .A3(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G226gat), .A2(G233gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT93), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n541_), .A2(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n544_), .B1(new_n538_), .B2(new_n525_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n525_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n378_), .A2(new_n549_), .ZN(new_n550_));
  AND3_X1   g349(.A1(new_n548_), .A2(new_n550_), .A3(KEYINPUT20), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n524_), .B1(new_n547_), .B2(new_n552_), .ZN(new_n553_));
  AOI211_X1 g352(.A(new_n523_), .B(new_n551_), .C1(new_n541_), .C2(new_n546_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n518_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n551_), .B1(new_n541_), .B2(new_n546_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n518_), .B1(new_n556_), .B2(new_n524_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n538_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n550_), .A2(new_n558_), .A3(KEYINPUT20), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(new_n544_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT98), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n529_), .A2(new_n530_), .A3(new_n540_), .A4(new_n545_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n559_), .A2(KEYINPUT98), .A3(new_n544_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n562_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(new_n523_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n557_), .A2(new_n566_), .ZN(new_n567_));
  AND4_X1   g366(.A1(new_n458_), .A2(new_n517_), .A3(new_n555_), .A4(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n539_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n545_), .B1(new_n569_), .B2(new_n530_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n523_), .B1(new_n570_), .B2(new_n551_), .ZN(new_n571_));
  AND3_X1   g370(.A1(new_n526_), .A2(KEYINPUT94), .A3(KEYINPUT20), .ZN(new_n572_));
  AOI21_X1  g371(.A(KEYINPUT94), .B1(new_n526_), .B2(KEYINPUT20), .ZN(new_n573_));
  NOR3_X1   g372(.A1(new_n572_), .A2(new_n573_), .A3(new_n539_), .ZN(new_n574_));
  OAI211_X1 g373(.A(new_n552_), .B(new_n524_), .C1(new_n574_), .C2(new_n545_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n571_), .A2(new_n575_), .ZN(new_n576_));
  AOI22_X1  g375(.A1(new_n518_), .A2(new_n576_), .B1(new_n557_), .B2(new_n566_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n458_), .B1(new_n577_), .B2(new_n517_), .ZN(new_n578_));
  OAI211_X1 g377(.A(new_n401_), .B(new_n457_), .C1(new_n568_), .C2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT86), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n397_), .A2(new_n580_), .A3(new_n399_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n580_), .B1(new_n397_), .B2(new_n399_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  AND3_X1   g383(.A1(new_n514_), .A2(new_n461_), .A3(new_n515_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n461_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(KEYINPUT97), .B1(new_n553_), .B2(new_n554_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT97), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n571_), .A2(new_n575_), .A3(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT33), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n455_), .A2(new_n591_), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n444_), .A2(new_n446_), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n593_), .A2(KEYINPUT33), .A3(new_n443_), .A4(new_n454_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n430_), .A2(new_n441_), .A3(new_n445_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n442_), .B1(new_n441_), .B2(KEYINPUT4), .ZN(new_n596_));
  OAI211_X1 g395(.A(new_n595_), .B(new_n452_), .C1(new_n444_), .C2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n592_), .A2(new_n594_), .A3(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n588_), .A2(new_n590_), .A3(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n524_), .A2(KEYINPUT32), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n565_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT99), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n565_), .A2(KEYINPUT99), .A3(new_n602_), .ZN(new_n606_));
  AOI22_X1  g405(.A1(new_n556_), .A2(new_n601_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n605_), .A2(new_n606_), .A3(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n587_), .B1(new_n600_), .B2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n555_), .A2(new_n567_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n513_), .A2(new_n516_), .A3(new_n457_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n584_), .B1(new_n609_), .B2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n579_), .A2(new_n613_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n335_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(G231gat), .A2(G233gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n313_), .B(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(new_n251_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT17), .ZN(new_n619_));
  XOR2_X1   g418(.A(G127gat), .B(G155gat), .Z(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT16), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G183gat), .B(G211gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  OR3_X1    g422(.A1(new_n618_), .A2(new_n619_), .A3(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(KEYINPUT17), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n618_), .A2(new_n625_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n624_), .A2(new_n626_), .ZN(new_n627_));
  XOR2_X1   g426(.A(new_n627_), .B(KEYINPUT77), .Z(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT37), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n321_), .A2(new_n253_), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n250_), .A2(new_n247_), .A3(new_n230_), .A4(new_n306_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(G232gat), .A2(G233gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT34), .ZN(new_n634_));
  OAI21_X1  g433(.A(KEYINPUT74), .B1(new_n634_), .B2(KEYINPUT35), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n631_), .A2(new_n632_), .A3(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n634_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT35), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n637_), .A2(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(G190gat), .B(G218gat), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT73), .ZN(new_n643_));
  XNOR2_X1  g442(.A(G134gat), .B(G162gat), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n643_), .B(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT36), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n635_), .B1(new_n321_), .B2(new_n253_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n640_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n648_), .A2(new_n649_), .A3(new_n632_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n641_), .A2(new_n647_), .A3(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT75), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n630_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n645_), .B(KEYINPUT36), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n648_), .A2(new_n649_), .A3(new_n632_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n649_), .B1(new_n648_), .B2(new_n632_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n654_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n657_), .A2(KEYINPUT76), .A3(new_n651_), .ZN(new_n658_));
  AOI21_X1  g457(.A(KEYINPUT76), .B1(new_n657_), .B2(new_n651_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n653_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT76), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n641_), .A2(new_n647_), .A3(new_n650_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n654_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n663_), .B1(new_n641_), .B2(new_n650_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n661_), .B1(new_n662_), .B2(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(KEYINPUT37), .B1(new_n662_), .B2(KEYINPUT75), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n657_), .A2(new_n651_), .A3(KEYINPUT76), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n665_), .A2(new_n666_), .A3(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n660_), .A2(new_n668_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n629_), .A2(new_n669_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n615_), .A2(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n671_), .A2(new_n308_), .A3(new_n456_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT38), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT101), .ZN(new_n675_));
  INV_X1    g474(.A(new_n627_), .ZN(new_n676_));
  NOR3_X1   g475(.A1(new_n281_), .A2(new_n676_), .A3(new_n330_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n657_), .A2(new_n651_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n679_), .B1(new_n579_), .B2(new_n613_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n677_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(G1gat), .B1(new_n682_), .B2(new_n457_), .ZN(new_n683_));
  OAI211_X1 g482(.A(new_n675_), .B(new_n683_), .C1(new_n673_), .C2(new_n672_), .ZN(G1324gat));
  AOI21_X1  g483(.A(new_n309_), .B1(new_n681_), .B2(new_n610_), .ZN(new_n685_));
  XOR2_X1   g484(.A(new_n685_), .B(KEYINPUT39), .Z(new_n686_));
  NAND3_X1  g485(.A1(new_n671_), .A2(new_n309_), .A3(new_n610_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  XOR2_X1   g487(.A(KEYINPUT102), .B(KEYINPUT40), .Z(new_n689_));
  XNOR2_X1  g488(.A(new_n688_), .B(new_n689_), .ZN(G1325gat));
  OAI21_X1  g489(.A(G15gat), .B1(new_n682_), .B2(new_n584_), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n691_), .A2(KEYINPUT41), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(KEYINPUT41), .ZN(new_n693_));
  INV_X1    g492(.A(G15gat), .ZN(new_n694_));
  INV_X1    g493(.A(new_n583_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(new_n581_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n671_), .A2(new_n694_), .A3(new_n696_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n692_), .A2(new_n693_), .A3(new_n697_), .ZN(G1326gat));
  INV_X1    g497(.A(G22gat), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n699_), .B1(new_n681_), .B2(new_n587_), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT42), .Z(new_n701_));
  NAND3_X1  g500(.A1(new_n671_), .A2(new_n699_), .A3(new_n587_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(G1327gat));
  NOR2_X1   g502(.A1(new_n628_), .A2(new_n678_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n615_), .A2(KEYINPUT106), .A3(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n335_), .A2(new_n614_), .A3(new_n704_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT106), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n705_), .A2(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(G29gat), .B1(new_n709_), .B2(new_n456_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT103), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n660_), .A2(new_n668_), .A3(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n711_), .B1(new_n660_), .B2(new_n668_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  OAI21_X1  g514(.A(KEYINPUT100), .B1(new_n610_), .B2(new_n587_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n577_), .A2(new_n458_), .A3(new_n517_), .ZN(new_n717_));
  AOI211_X1 g516(.A(new_n400_), .B(new_n456_), .C1(new_n716_), .C2(new_n717_), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n571_), .A2(new_n589_), .A3(new_n575_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n589_), .B1(new_n571_), .B2(new_n575_), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n719_), .A2(new_n720_), .A3(new_n598_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n606_), .A2(new_n607_), .ZN(new_n722_));
  AOI21_X1  g521(.A(KEYINPUT99), .B1(new_n565_), .B2(new_n602_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n517_), .B1(new_n721_), .B2(new_n724_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n577_), .A2(new_n587_), .A3(new_n457_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n696_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n715_), .B1(new_n718_), .B2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(KEYINPUT43), .ZN(new_n729_));
  INV_X1    g528(.A(new_n669_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n730_), .A2(KEYINPUT43), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n731_), .B1(new_n718_), .B2(new_n727_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n628_), .B1(new_n729_), .B2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT105), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n281_), .A2(new_n330_), .ZN(new_n735_));
  NAND4_X1  g534(.A1(new_n733_), .A2(new_n734_), .A3(KEYINPUT44), .A4(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT43), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n714_), .B1(new_n579_), .B2(new_n613_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n732_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n739_), .A2(KEYINPUT44), .A3(new_n629_), .A4(new_n735_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT105), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n736_), .A2(new_n741_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n739_), .A2(new_n629_), .A3(new_n735_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(KEYINPUT104), .B(KEYINPUT44), .ZN(new_n744_));
  AOI211_X1 g543(.A(new_n286_), .B(new_n457_), .C1(new_n743_), .C2(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n710_), .B1(new_n742_), .B2(new_n745_), .ZN(G1328gat));
  AOI21_X1  g545(.A(new_n577_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n740_), .A2(KEYINPUT105), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n740_), .A2(KEYINPUT105), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n747_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(G36gat), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT107), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT46), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n705_), .A2(new_n284_), .A3(new_n610_), .A4(new_n708_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT45), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n751_), .A2(new_n752_), .A3(new_n753_), .A4(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n752_), .A2(new_n753_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n284_), .B1(new_n742_), .B2(new_n747_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT45), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n754_), .B(new_n760_), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n757_), .B(new_n758_), .C1(new_n759_), .C2(new_n761_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n756_), .A2(new_n762_), .ZN(G1329gat));
  NAND2_X1  g562(.A1(new_n743_), .A2(new_n744_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n742_), .A2(G43gat), .A3(new_n401_), .A4(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n705_), .A2(new_n696_), .A3(new_n708_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(new_n291_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT108), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n766_), .A2(KEYINPUT108), .A3(new_n291_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n765_), .A2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT47), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT47), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n765_), .A2(new_n771_), .A3(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(G1330gat));
  NAND3_X1  g575(.A1(new_n709_), .A2(new_n289_), .A3(new_n587_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n742_), .A2(new_n587_), .A3(new_n764_), .ZN(new_n778_));
  AND3_X1   g577(.A1(new_n778_), .A2(KEYINPUT109), .A3(G50gat), .ZN(new_n779_));
  AOI21_X1  g578(.A(KEYINPUT109), .B1(new_n778_), .B2(G50gat), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n777_), .B1(new_n779_), .B2(new_n780_), .ZN(G1331gat));
  AND2_X1   g580(.A1(new_n279_), .A2(new_n280_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n782_), .A2(new_n329_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n783_), .A2(new_n614_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n784_), .A2(new_n670_), .ZN(new_n785_));
  AOI21_X1  g584(.A(G57gat), .B1(new_n785_), .B2(new_n456_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n786_), .A2(KEYINPUT110), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n786_), .A2(KEYINPUT110), .ZN(new_n788_));
  INV_X1    g587(.A(new_n334_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n789_), .A2(new_n629_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n680_), .A2(new_n281_), .A3(new_n790_), .ZN(new_n791_));
  XOR2_X1   g590(.A(KEYINPUT111), .B(G57gat), .Z(new_n792_));
  NOR3_X1   g591(.A1(new_n791_), .A2(new_n457_), .A3(new_n792_), .ZN(new_n793_));
  NOR3_X1   g592(.A1(new_n787_), .A2(new_n788_), .A3(new_n793_), .ZN(G1332gat));
  OAI21_X1  g593(.A(G64gat), .B1(new_n791_), .B2(new_n577_), .ZN(new_n795_));
  XOR2_X1   g594(.A(KEYINPUT112), .B(KEYINPUT48), .Z(new_n796_));
  XNOR2_X1  g595(.A(new_n795_), .B(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(G64gat), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n785_), .A2(new_n798_), .A3(new_n610_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n797_), .A2(new_n799_), .ZN(G1333gat));
  OAI21_X1  g599(.A(G71gat), .B1(new_n791_), .B2(new_n584_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n801_), .B(KEYINPUT49), .ZN(new_n802_));
  INV_X1    g601(.A(G71gat), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n785_), .A2(new_n803_), .A3(new_n696_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n802_), .A2(new_n804_), .ZN(G1334gat));
  OAI21_X1  g604(.A(G78gat), .B1(new_n791_), .B2(new_n517_), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n806_), .B(KEYINPUT50), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n517_), .A2(G78gat), .ZN(new_n808_));
  XOR2_X1   g607(.A(new_n808_), .B(KEYINPUT113), .Z(new_n809_));
  NAND2_X1  g608(.A1(new_n785_), .A2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n807_), .A2(new_n810_), .ZN(G1335gat));
  NAND2_X1  g610(.A1(new_n733_), .A2(new_n783_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT114), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n733_), .A2(KEYINPUT114), .A3(new_n783_), .ZN(new_n815_));
  AND2_X1   g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(G85gat), .B1(new_n816_), .B2(new_n457_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n784_), .A2(new_n704_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n818_), .A2(new_n218_), .A3(new_n456_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n817_), .A2(new_n819_), .ZN(G1336gat));
  OAI21_X1  g619(.A(G92gat), .B1(new_n816_), .B2(new_n577_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n818_), .A2(new_n219_), .A3(new_n610_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(G1337gat));
  OAI21_X1  g622(.A(G99gat), .B1(new_n816_), .B2(new_n584_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT51), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n818_), .A2(new_n215_), .A3(new_n401_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n824_), .A2(new_n825_), .A3(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n814_), .A2(new_n815_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n232_), .B1(new_n828_), .B2(new_n696_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n826_), .ZN(new_n830_));
  OAI21_X1  g629(.A(KEYINPUT51), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n827_), .A2(new_n831_), .ZN(G1338gat));
  INV_X1    g631(.A(KEYINPUT52), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n739_), .A2(new_n629_), .A3(new_n587_), .A4(new_n783_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT115), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n834_), .A2(new_n835_), .A3(G106gat), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n835_), .B1(new_n834_), .B2(G106gat), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n833_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n838_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n840_), .A2(KEYINPUT52), .A3(new_n836_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n818_), .A2(new_n216_), .A3(new_n587_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n839_), .A2(new_n841_), .A3(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(KEYINPUT53), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n839_), .A2(new_n841_), .A3(new_n845_), .A4(new_n842_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n846_), .ZN(G1339gat));
  AOI21_X1  g646(.A(new_n400_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n456_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT121), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n322_), .A2(new_n323_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n328_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n853_));
  AOI22_X1  g652(.A1(new_n324_), .A2(new_n328_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  AND2_X1   g653(.A1(new_n854_), .A2(new_n274_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT55), .ZN(new_n856_));
  OR2_X1    g655(.A1(new_n256_), .A2(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n246_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n858_));
  AND3_X1   g657(.A1(new_n858_), .A2(KEYINPUT117), .A3(new_n263_), .ZN(new_n859_));
  AOI21_X1  g658(.A(KEYINPUT117), .B1(new_n858_), .B2(new_n263_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n857_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  AND3_X1   g660(.A1(new_n258_), .A2(new_n261_), .A3(new_n856_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n272_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT56), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n258_), .A2(new_n261_), .A3(new_n856_), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n866_), .B(new_n857_), .C1(new_n860_), .C2(new_n859_), .ZN(new_n867_));
  AOI21_X1  g666(.A(KEYINPUT56), .B1(new_n867_), .B2(new_n272_), .ZN(new_n868_));
  OAI211_X1 g667(.A(KEYINPUT58), .B(new_n855_), .C1(new_n865_), .C2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n669_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n863_), .A2(new_n864_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n867_), .A2(KEYINPUT56), .A3(new_n272_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(KEYINPUT58), .B1(new_n873_), .B2(new_n855_), .ZN(new_n874_));
  OR2_X1    g673(.A1(new_n870_), .A2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n329_), .A2(new_n274_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  XOR2_X1   g676(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n878_));
  AOI21_X1  g677(.A(new_n878_), .B1(new_n867_), .B2(new_n272_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n877_), .B1(new_n865_), .B2(new_n879_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n275_), .A2(new_n277_), .A3(new_n854_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n679_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(KEYINPUT120), .B1(new_n882_), .B2(KEYINPUT57), .ZN(new_n883_));
  INV_X1    g682(.A(new_n878_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n863_), .A2(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n876_), .B1(new_n885_), .B2(new_n872_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n881_), .ZN(new_n887_));
  OAI211_X1 g686(.A(KEYINPUT57), .B(new_n678_), .C1(new_n886_), .C2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT120), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n875_), .B1(new_n883_), .B2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT119), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n882_), .A2(new_n892_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n678_), .B1(new_n886_), .B2(new_n887_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(KEYINPUT119), .ZN(new_n895_));
  AOI21_X1  g694(.A(KEYINPUT57), .B1(new_n893_), .B2(new_n895_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n851_), .B1(new_n891_), .B2(new_n896_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n870_), .A2(new_n874_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n882_), .A2(KEYINPUT120), .A3(KEYINPUT57), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n888_), .A2(new_n889_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n898_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT57), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n882_), .A2(new_n892_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n894_), .A2(KEYINPUT119), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n902_), .B1(new_n903_), .B2(new_n904_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n901_), .A2(new_n905_), .A3(KEYINPUT121), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n627_), .B1(new_n897_), .B2(new_n906_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n790_), .A2(new_n782_), .A3(new_n730_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT116), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n908_), .A2(new_n909_), .A3(KEYINPUT54), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n910_), .B1(KEYINPUT54), .B2(new_n908_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n909_), .B1(new_n908_), .B2(KEYINPUT54), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n911_), .A2(new_n912_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n850_), .B1(new_n907_), .B2(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT122), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n891_), .A2(new_n851_), .A3(new_n896_), .ZN(new_n917_));
  AOI21_X1  g716(.A(KEYINPUT121), .B1(new_n901_), .B2(new_n905_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n676_), .B1(new_n917_), .B2(new_n918_), .ZN(new_n919_));
  OR2_X1    g718(.A1(new_n911_), .A2(new_n912_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n921_), .A2(KEYINPUT122), .A3(new_n850_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n916_), .A2(new_n922_), .A3(new_n329_), .ZN(new_n923_));
  INV_X1    g722(.A(G113gat), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n628_), .B1(new_n901_), .B2(new_n905_), .ZN(new_n925_));
  OR2_X1    g724(.A1(new_n913_), .A2(new_n925_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n849_), .B(KEYINPUT123), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n927_), .A2(KEYINPUT59), .ZN(new_n928_));
  AOI22_X1  g727(.A1(new_n914_), .A2(KEYINPUT59), .B1(new_n926_), .B2(new_n928_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(KEYINPUT124), .B(G113gat), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n789_), .A2(new_n930_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(KEYINPUT125), .ZN(new_n932_));
  AOI22_X1  g731(.A1(new_n923_), .A2(new_n924_), .B1(new_n929_), .B2(new_n932_), .ZN(G1340gat));
  OAI21_X1  g732(.A(new_n928_), .B1(new_n913_), .B2(new_n925_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n849_), .B1(new_n919_), .B2(new_n920_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT59), .ZN(new_n936_));
  OAI211_X1 g735(.A(new_n281_), .B(new_n934_), .C1(new_n935_), .C2(new_n936_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n937_), .A2(G120gat), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT60), .ZN(new_n939_));
  INV_X1    g738(.A(G120gat), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n281_), .A2(new_n939_), .A3(new_n940_), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n941_), .B1(new_n939_), .B2(new_n940_), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n916_), .A2(new_n922_), .A3(new_n942_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n938_), .A2(new_n943_), .ZN(G1341gat));
  OAI211_X1 g743(.A(new_n627_), .B(new_n934_), .C1(new_n935_), .C2(new_n936_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n945_), .A2(G127gat), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n629_), .A2(G127gat), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n916_), .A2(new_n922_), .A3(new_n947_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n946_), .A2(new_n948_), .ZN(G1342gat));
  OAI211_X1 g748(.A(new_n669_), .B(new_n934_), .C1(new_n935_), .C2(new_n936_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n950_), .A2(G134gat), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n678_), .A2(G134gat), .ZN(new_n952_));
  NAND3_X1  g751(.A1(new_n916_), .A2(new_n922_), .A3(new_n952_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n951_), .A2(new_n953_), .ZN(G1343gat));
  NAND2_X1  g753(.A1(new_n584_), .A2(new_n587_), .ZN(new_n955_));
  NOR3_X1   g754(.A1(new_n955_), .A2(new_n457_), .A3(new_n610_), .ZN(new_n956_));
  NAND3_X1  g755(.A1(new_n921_), .A2(new_n329_), .A3(new_n956_), .ZN(new_n957_));
  XOR2_X1   g756(.A(KEYINPUT126), .B(G141gat), .Z(new_n958_));
  XNOR2_X1  g757(.A(new_n957_), .B(new_n958_), .ZN(G1344gat));
  NAND3_X1  g758(.A1(new_n921_), .A2(new_n281_), .A3(new_n956_), .ZN(new_n960_));
  XOR2_X1   g759(.A(KEYINPUT127), .B(G148gat), .Z(new_n961_));
  XNOR2_X1  g760(.A(new_n960_), .B(new_n961_), .ZN(G1345gat));
  NAND3_X1  g761(.A1(new_n921_), .A2(new_n628_), .A3(new_n956_), .ZN(new_n963_));
  XNOR2_X1  g762(.A(KEYINPUT61), .B(G155gat), .ZN(new_n964_));
  XNOR2_X1  g763(.A(new_n963_), .B(new_n964_), .ZN(G1346gat));
  AND4_X1   g764(.A1(G162gat), .A2(new_n921_), .A3(new_n715_), .A4(new_n956_), .ZN(new_n966_));
  NAND3_X1  g765(.A1(new_n921_), .A2(new_n679_), .A3(new_n956_), .ZN(new_n967_));
  AOI21_X1  g766(.A(new_n966_), .B1(new_n427_), .B2(new_n967_), .ZN(G1347gat));
  INV_X1    g767(.A(KEYINPUT62), .ZN(new_n969_));
  NOR2_X1   g768(.A1(new_n577_), .A2(new_n456_), .ZN(new_n970_));
  INV_X1    g769(.A(new_n970_), .ZN(new_n971_));
  NOR2_X1   g770(.A1(new_n971_), .A2(new_n584_), .ZN(new_n972_));
  INV_X1    g771(.A(new_n972_), .ZN(new_n973_));
  NOR2_X1   g772(.A1(new_n973_), .A2(new_n587_), .ZN(new_n974_));
  OAI211_X1 g773(.A(new_n329_), .B(new_n974_), .C1(new_n913_), .C2(new_n925_), .ZN(new_n975_));
  INV_X1    g774(.A(new_n975_), .ZN(new_n976_));
  OAI21_X1  g775(.A(new_n969_), .B1(new_n976_), .B2(new_n336_), .ZN(new_n977_));
  NAND3_X1  g776(.A1(new_n975_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n978_));
  NAND2_X1  g777(.A1(new_n976_), .A2(new_n372_), .ZN(new_n979_));
  NAND3_X1  g778(.A1(new_n977_), .A2(new_n978_), .A3(new_n979_), .ZN(G1348gat));
  NAND2_X1  g779(.A1(new_n926_), .A2(new_n974_), .ZN(new_n981_));
  INV_X1    g780(.A(new_n981_), .ZN(new_n982_));
  NAND2_X1  g781(.A1(new_n982_), .A2(new_n281_), .ZN(new_n983_));
  AOI21_X1  g782(.A(new_n587_), .B1(new_n919_), .B2(new_n920_), .ZN(new_n984_));
  NOR3_X1   g783(.A1(new_n973_), .A2(new_n782_), .A3(new_n337_), .ZN(new_n985_));
  AOI22_X1  g784(.A1(new_n983_), .A2(new_n337_), .B1(new_n984_), .B2(new_n985_), .ZN(G1349gat));
  NAND3_X1  g785(.A1(new_n984_), .A2(new_n628_), .A3(new_n972_), .ZN(new_n987_));
  AOI21_X1  g786(.A(new_n676_), .B1(new_n354_), .B2(new_n356_), .ZN(new_n988_));
  AOI22_X1  g787(.A1(new_n355_), .A2(new_n987_), .B1(new_n982_), .B2(new_n988_), .ZN(G1350gat));
  OAI21_X1  g788(.A(G190gat), .B1(new_n981_), .B2(new_n730_), .ZN(new_n990_));
  OR2_X1    g789(.A1(new_n678_), .A2(new_n351_), .ZN(new_n991_));
  OAI21_X1  g790(.A(new_n990_), .B1(new_n981_), .B2(new_n991_), .ZN(G1351gat));
  NOR2_X1   g791(.A1(new_n955_), .A2(new_n971_), .ZN(new_n993_));
  NAND3_X1  g792(.A1(new_n921_), .A2(new_n329_), .A3(new_n993_), .ZN(new_n994_));
  XNOR2_X1  g793(.A(new_n994_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g794(.A1(new_n921_), .A2(new_n993_), .ZN(new_n996_));
  OR3_X1    g795(.A1(new_n996_), .A2(G204gat), .A3(new_n782_), .ZN(new_n997_));
  OAI21_X1  g796(.A(G204gat), .B1(new_n996_), .B2(new_n782_), .ZN(new_n998_));
  NAND2_X1  g797(.A1(new_n997_), .A2(new_n998_), .ZN(G1353gat));
  INV_X1    g798(.A(new_n996_), .ZN(new_n1000_));
  XNOR2_X1  g799(.A(KEYINPUT63), .B(G211gat), .ZN(new_n1001_));
  NAND3_X1  g800(.A1(new_n1000_), .A2(new_n627_), .A3(new_n1001_), .ZN(new_n1002_));
  NOR2_X1   g801(.A1(new_n996_), .A2(new_n676_), .ZN(new_n1003_));
  NOR2_X1   g802(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1004_));
  OAI21_X1  g803(.A(new_n1002_), .B1(new_n1003_), .B2(new_n1004_), .ZN(G1354gat));
  OAI21_X1  g804(.A(G218gat), .B1(new_n996_), .B2(new_n730_), .ZN(new_n1006_));
  NAND2_X1  g805(.A1(new_n679_), .A2(new_n465_), .ZN(new_n1007_));
  OAI21_X1  g806(.A(new_n1006_), .B1(new_n996_), .B2(new_n1007_), .ZN(G1355gat));
endmodule


