//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 1 0 0 1 1 1 0 0 0 1 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 0 0 0 1 1 1 0 1 0 0 1 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n615_, new_n616_, new_n617_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n814_, new_n815_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n823_, new_n824_, new_n825_, new_n826_, new_n828_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n863_,
    new_n864_, new_n866_, new_n867_, new_n869_, new_n870_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n885_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT31), .ZN(new_n205_));
  INV_X1    g004(.A(G183gat), .ZN(new_n206_));
  INV_X1    g005(.A(G190gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT23), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT77), .B(KEYINPUT23), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n208_), .B(new_n211_), .C1(new_n212_), .C2(new_n209_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT79), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n209_), .ZN(new_n216_));
  AND2_X1   g015(.A1(new_n210_), .A2(KEYINPUT77), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n210_), .A2(KEYINPUT77), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n216_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n219_), .A2(KEYINPUT79), .A3(new_n208_), .A4(new_n211_), .ZN(new_n220_));
  INV_X1    g019(.A(G169gat), .ZN(new_n221_));
  INV_X1    g020(.A(G176gat), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT78), .ZN(new_n224_));
  AND2_X1   g023(.A1(new_n221_), .A2(KEYINPUT22), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n221_), .A2(KEYINPUT22), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n224_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n221_), .A2(KEYINPUT22), .ZN(new_n228_));
  AOI21_X1  g027(.A(G176gat), .B1(new_n228_), .B2(KEYINPUT78), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n223_), .B1(new_n227_), .B2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n215_), .A2(new_n220_), .A3(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n207_), .A2(KEYINPUT26), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT26), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(G190gat), .ZN(new_n234_));
  AND2_X1   g033(.A1(new_n232_), .A2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT25), .B(G183gat), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT24), .ZN(new_n237_));
  NOR2_X1   g036(.A1(G169gat), .A2(G176gat), .ZN(new_n238_));
  AOI22_X1  g037(.A1(new_n235_), .A2(new_n236_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n216_), .A2(new_n210_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n240_), .B1(new_n212_), .B2(new_n216_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n223_), .A2(new_n238_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT24), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n239_), .A2(new_n241_), .A3(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n231_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G227gat), .A2(G233gat), .ZN(new_n246_));
  INV_X1    g045(.A(G71gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(G99gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n245_), .B(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G15gat), .B(G43gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT80), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT30), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n250_), .B(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT81), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n205_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n256_), .B1(new_n255_), .B2(new_n254_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n254_), .A2(new_n255_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(new_n205_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G155gat), .A2(G162gat), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(G155gat), .A2(G162gat), .ZN(new_n263_));
  NOR3_X1   g062(.A1(new_n262_), .A2(new_n263_), .A3(KEYINPUT1), .ZN(new_n264_));
  OR2_X1    g063(.A1(G141gat), .A2(G148gat), .ZN(new_n265_));
  NAND3_X1  g064(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G141gat), .A2(G148gat), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n265_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  OAI21_X1  g067(.A(KEYINPUT82), .B1(new_n264_), .B2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n263_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT1), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n270_), .A2(new_n271_), .A3(new_n261_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n267_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(G141gat), .A2(G148gat), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT82), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n272_), .A2(new_n275_), .A3(new_n276_), .A4(new_n266_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n269_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT83), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n267_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(KEYINPUT2), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT2), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n267_), .A2(new_n279_), .A3(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT3), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n274_), .A2(new_n284_), .ZN(new_n285_));
  OAI21_X1  g084(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n281_), .A2(new_n283_), .A3(new_n285_), .A4(new_n286_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n262_), .A2(new_n263_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n278_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n204_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  AOI22_X1  g091(.A1(new_n269_), .A2(new_n277_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(new_n204_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n292_), .A2(KEYINPUT4), .A3(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G225gat), .A2(G233gat), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT98), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n204_), .B1(new_n278_), .B2(new_n289_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT4), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n298_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  NOR4_X1   g100(.A1(new_n293_), .A2(KEYINPUT98), .A3(KEYINPUT4), .A4(new_n204_), .ZN(new_n302_));
  OAI211_X1 g101(.A(new_n295_), .B(new_n297_), .C1(new_n301_), .C2(new_n302_), .ZN(new_n303_));
  AND2_X1   g102(.A1(new_n292_), .A2(new_n294_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(new_n296_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G1gat), .B(G29gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(G85gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(KEYINPUT0), .B(G57gat), .ZN(new_n309_));
  XOR2_X1   g108(.A(new_n308_), .B(new_n309_), .Z(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n306_), .A2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n303_), .A2(new_n305_), .A3(new_n310_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n260_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(G204gat), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT87), .B1(new_n316_), .B2(G197gat), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT87), .ZN(new_n318_));
  INV_X1    g117(.A(G197gat), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n318_), .A2(new_n319_), .A3(G204gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n316_), .A2(G197gat), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n317_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(KEYINPUT88), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT88), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n317_), .A2(new_n320_), .A3(new_n324_), .A4(new_n321_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G211gat), .B(G218gat), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT21), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n323_), .A2(new_n325_), .A3(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n316_), .A2(G197gat), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n319_), .A2(G204gat), .ZN(new_n331_));
  OAI21_X1  g130(.A(KEYINPUT21), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  OAI211_X1 g131(.A(new_n332_), .B(new_n326_), .C1(new_n322_), .C2(KEYINPUT21), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n329_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT29), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n334_), .B1(new_n293_), .B2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT86), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT89), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT89), .ZN(new_n339_));
  OAI211_X1 g138(.A(new_n334_), .B(new_n339_), .C1(new_n293_), .C2(new_n335_), .ZN(new_n340_));
  INV_X1    g139(.A(G228gat), .ZN(new_n341_));
  INV_X1    g140(.A(G233gat), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n338_), .A2(new_n340_), .A3(new_n343_), .ZN(new_n344_));
  OAI221_X1 g143(.A(KEYINPUT89), .B1(new_n341_), .B2(new_n342_), .C1(new_n336_), .C2(new_n337_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G78gat), .B(G106gat), .ZN(new_n347_));
  XOR2_X1   g146(.A(new_n347_), .B(KEYINPUT90), .Z(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(new_n348_), .ZN(new_n349_));
  XOR2_X1   g148(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n350_));
  INV_X1    g149(.A(KEYINPUT84), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n293_), .A2(new_n351_), .A3(new_n335_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n351_), .B1(new_n293_), .B2(new_n335_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n350_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n354_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n350_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n356_), .A2(new_n352_), .A3(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G22gat), .B(G50gat), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n355_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n359_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n357_), .B1(new_n356_), .B2(new_n352_), .ZN(new_n362_));
  NOR3_X1   g161(.A1(new_n353_), .A2(new_n354_), .A3(new_n350_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n361_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n344_), .A2(new_n345_), .A3(new_n347_), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n349_), .A2(new_n360_), .A3(new_n364_), .A4(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT91), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  AND2_X1   g167(.A1(new_n364_), .A2(new_n360_), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n369_), .A2(KEYINPUT91), .A3(new_n349_), .A4(new_n365_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n346_), .B(new_n348_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n369_), .ZN(new_n372_));
  AOI22_X1  g171(.A1(new_n368_), .A2(new_n370_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  XOR2_X1   g172(.A(G8gat), .B(G36gat), .Z(new_n374_));
  XNOR2_X1  g173(.A(G64gat), .B(G92gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT96), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G226gat), .A2(G233gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT19), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n231_), .A2(new_n244_), .A3(new_n333_), .A4(new_n329_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT92), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n382_), .A2(new_n383_), .A3(KEYINPUT20), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n232_), .A2(new_n234_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT93), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n232_), .A2(new_n234_), .A3(KEYINPUT93), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n387_), .A2(new_n236_), .A3(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT94), .B(KEYINPUT24), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n242_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n238_), .ZN(new_n393_));
  OR2_X1    g192(.A1(new_n390_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT95), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n394_), .A2(new_n395_), .A3(new_n219_), .A4(new_n211_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n211_), .B1(new_n212_), .B2(new_n209_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n390_), .A2(new_n393_), .ZN(new_n398_));
  OAI21_X1  g197(.A(KEYINPUT95), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n392_), .B1(new_n396_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n223_), .ZN(new_n401_));
  XOR2_X1   g200(.A(KEYINPUT22), .B(G169gat), .Z(new_n402_));
  OAI21_X1  g201(.A(new_n401_), .B1(new_n402_), .B2(G176gat), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n403_), .B1(new_n241_), .B2(new_n208_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n334_), .B1(new_n400_), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n384_), .A2(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n383_), .B1(new_n382_), .B2(KEYINPUT20), .ZN(new_n407_));
  OAI211_X1 g206(.A(new_n379_), .B(new_n381_), .C1(new_n406_), .C2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n396_), .A2(new_n399_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n392_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n404_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n411_), .A2(new_n333_), .A3(new_n329_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n381_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n245_), .A2(new_n334_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n412_), .A2(KEYINPUT20), .A3(new_n413_), .A4(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n408_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n382_), .A2(KEYINPUT20), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT92), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n418_), .A2(new_n405_), .A3(new_n384_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n379_), .B1(new_n419_), .B2(new_n381_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n378_), .B1(new_n416_), .B2(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n381_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT96), .ZN(new_n423_));
  INV_X1    g222(.A(new_n378_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n423_), .A2(new_n424_), .A3(new_n415_), .A4(new_n408_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n421_), .A2(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(KEYINPUT102), .B(KEYINPUT27), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT27), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n412_), .A2(KEYINPUT20), .A3(new_n414_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(new_n381_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n431_), .B1(new_n419_), .B2(new_n381_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n429_), .B1(new_n432_), .B2(new_n378_), .ZN(new_n433_));
  AOI22_X1  g232(.A1(new_n426_), .A2(new_n428_), .B1(new_n425_), .B2(new_n433_), .ZN(new_n434_));
  AND3_X1   g233(.A1(new_n315_), .A2(new_n373_), .A3(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n424_), .A2(KEYINPUT32), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n423_), .A2(new_n415_), .A3(new_n408_), .A4(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n436_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n432_), .A2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n437_), .A2(new_n439_), .A3(new_n314_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n304_), .A2(new_n297_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(new_n311_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT100), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n295_), .B(new_n296_), .C1(new_n301_), .C2(new_n302_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT100), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n441_), .A2(new_n445_), .A3(new_n311_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n443_), .A2(new_n444_), .A3(new_n446_), .ZN(new_n447_));
  AND3_X1   g246(.A1(new_n313_), .A2(KEYINPUT99), .A3(KEYINPUT33), .ZN(new_n448_));
  AOI21_X1  g247(.A(KEYINPUT33), .B1(new_n313_), .B2(KEYINPUT99), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n447_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n440_), .B1(new_n426_), .B2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(new_n373_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT101), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT101), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n451_), .A2(new_n373_), .A3(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n368_), .A2(new_n370_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n371_), .A2(new_n372_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n314_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(new_n434_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n453_), .A2(new_n455_), .A3(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n435_), .B1(new_n460_), .B2(new_n260_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G85gat), .B(G92gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(KEYINPUT66), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT8), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G99gat), .A2(G106gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(KEYINPUT6), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(G99gat), .A2(G106gat), .ZN(new_n468_));
  XOR2_X1   g267(.A(new_n468_), .B(KEYINPUT7), .Z(new_n469_));
  OAI211_X1 g268(.A(new_n463_), .B(new_n464_), .C1(new_n467_), .C2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT67), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  OR2_X1    g271(.A1(new_n469_), .A2(new_n467_), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n473_), .A2(KEYINPUT67), .A3(new_n464_), .A4(new_n463_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n463_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT68), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n469_), .B1(new_n476_), .B2(new_n466_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n467_), .A2(KEYINPUT68), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n475_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n472_), .B(new_n474_), .C1(new_n479_), .C2(new_n464_), .ZN(new_n480_));
  XOR2_X1   g279(.A(KEYINPUT10), .B(G99gat), .Z(new_n481_));
  XNOR2_X1  g280(.A(KEYINPUT64), .B(G106gat), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n467_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT9), .ZN(new_n484_));
  XOR2_X1   g283(.A(KEYINPUT65), .B(G85gat), .Z(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(G92gat), .ZN(new_n486_));
  OAI221_X1 g285(.A(new_n483_), .B1(new_n484_), .B2(new_n462_), .C1(new_n485_), .C2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n480_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT70), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n480_), .A2(KEYINPUT70), .A3(new_n487_), .ZN(new_n491_));
  XOR2_X1   g290(.A(G29gat), .B(G36gat), .Z(new_n492_));
  XOR2_X1   g291(.A(G43gat), .B(G50gat), .Z(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT15), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n490_), .A2(new_n491_), .A3(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n480_), .A2(new_n487_), .A3(new_n494_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G232gat), .A2(G233gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT34), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G190gat), .B(G218gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G134gat), .B(G162gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n502_), .B(new_n503_), .ZN(new_n504_));
  AOI22_X1  g303(.A1(new_n498_), .A2(new_n501_), .B1(KEYINPUT36), .B2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n500_), .B(KEYINPUT71), .ZN(new_n506_));
  XOR2_X1   g305(.A(new_n506_), .B(KEYINPUT35), .Z(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n508_), .B1(new_n498_), .B2(KEYINPUT72), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT72), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n496_), .A2(new_n510_), .A3(new_n497_), .A4(new_n507_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n505_), .A2(new_n509_), .A3(new_n511_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n504_), .A2(KEYINPUT36), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n513_), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n505_), .A2(new_n509_), .A3(new_n515_), .A4(new_n511_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n514_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n461_), .A2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G57gat), .B(G64gat), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n520_), .A2(KEYINPUT11), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(KEYINPUT11), .ZN(new_n522_));
  XOR2_X1   g321(.A(G71gat), .B(G78gat), .Z(new_n523_));
  NAND3_X1  g322(.A1(new_n521_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  OR2_X1    g323(.A1(new_n522_), .A2(new_n523_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n488_), .A2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n480_), .A2(new_n487_), .A3(new_n526_), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT69), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G230gat), .A2(G233gat), .ZN(new_n532_));
  OR3_X1    g331(.A1(new_n530_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n529_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT12), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n534_), .B1(new_n535_), .B2(new_n528_), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n490_), .A2(KEYINPUT12), .A3(new_n491_), .A4(new_n527_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n536_), .A2(new_n532_), .A3(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n531_), .B1(new_n530_), .B2(new_n532_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n533_), .A2(new_n538_), .A3(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G120gat), .B(G148gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT5), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G176gat), .B(G204gat), .ZN(new_n543_));
  XOR2_X1   g342(.A(new_n542_), .B(new_n543_), .Z(new_n544_));
  NAND2_X1  g343(.A1(new_n540_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n544_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n533_), .A2(new_n538_), .A3(new_n539_), .A4(new_n546_), .ZN(new_n547_));
  AND3_X1   g346(.A1(new_n545_), .A2(KEYINPUT13), .A3(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(KEYINPUT13), .B1(new_n545_), .B2(new_n547_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G231gat), .A2(G233gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n526_), .B(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G1gat), .B(G8gat), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT73), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  OR2_X1    g355(.A1(G15gat), .A2(G22gat), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G15gat), .A2(G22gat), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G1gat), .A2(G8gat), .ZN(new_n559_));
  AOI22_X1  g358(.A1(new_n557_), .A2(new_n558_), .B1(KEYINPUT14), .B2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n556_), .B(new_n560_), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n553_), .B(new_n561_), .Z(new_n562_));
  XOR2_X1   g361(.A(G127gat), .B(G155gat), .Z(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT16), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G183gat), .B(G211gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT17), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  AND2_X1   g367(.A1(new_n566_), .A2(new_n567_), .ZN(new_n569_));
  NOR3_X1   g368(.A1(new_n562_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n562_), .A2(new_n568_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n494_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n561_), .A2(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n575_), .B1(new_n495_), .B2(new_n561_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G229gat), .A2(G233gat), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n561_), .B(new_n574_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n577_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n578_), .A2(KEYINPUT74), .A3(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n582_), .B1(KEYINPUT74), .B2(new_n578_), .ZN(new_n583_));
  XOR2_X1   g382(.A(G113gat), .B(G141gat), .Z(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT75), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G169gat), .B(G197gat), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n585_), .B(new_n586_), .Z(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n583_), .A2(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(KEYINPUT76), .B1(new_n583_), .B2(new_n588_), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n589_), .A2(new_n590_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NOR3_X1   g392(.A1(new_n551_), .A2(new_n573_), .A3(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n519_), .A2(new_n594_), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n595_), .B(KEYINPUT103), .Z(new_n596_));
  INV_X1    g395(.A(new_n314_), .ZN(new_n597_));
  OAI21_X1  g396(.A(G1gat), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n598_), .B(KEYINPUT104), .Z(new_n599_));
  NOR2_X1   g398(.A1(new_n461_), .A2(new_n593_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT37), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n517_), .A2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n514_), .A2(KEYINPUT37), .A3(new_n516_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n604_), .A2(new_n573_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n600_), .A2(new_n550_), .A3(new_n605_), .ZN(new_n606_));
  NOR3_X1   g405(.A1(new_n606_), .A2(G1gat), .A3(new_n597_), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n607_), .B(KEYINPUT38), .Z(new_n608_));
  NAND2_X1  g407(.A1(new_n599_), .A2(new_n608_), .ZN(G1324gat));
  OAI21_X1  g408(.A(G8gat), .B1(new_n595_), .B2(new_n434_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT39), .ZN(new_n611_));
  OR2_X1    g410(.A1(new_n434_), .A2(G8gat), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n611_), .B1(new_n606_), .B2(new_n612_), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n613_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g413(.A(G15gat), .B1(new_n596_), .B2(new_n260_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT41), .ZN(new_n616_));
  NOR3_X1   g415(.A1(new_n606_), .A2(G15gat), .A3(new_n260_), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n616_), .A2(new_n617_), .ZN(G1326gat));
  OAI21_X1  g417(.A(G22gat), .B1(new_n596_), .B2(new_n373_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n373_), .A2(G22gat), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n621_), .B1(new_n606_), .B2(new_n622_), .ZN(G1327gat));
  XOR2_X1   g422(.A(KEYINPUT108), .B(KEYINPUT44), .Z(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n603_), .ZN(new_n626_));
  AOI21_X1  g425(.A(KEYINPUT37), .B1(new_n514_), .B2(new_n516_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n460_), .A2(new_n260_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n435_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n628_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT43), .ZN(new_n632_));
  OAI21_X1  g431(.A(KEYINPUT106), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT106), .ZN(new_n634_));
  OAI211_X1 g433(.A(new_n634_), .B(KEYINPUT43), .C1(new_n461_), .C2(new_n628_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n260_), .ZN(new_n636_));
  AOI22_X1  g435(.A1(new_n452_), .A2(KEYINPUT101), .B1(new_n458_), .B2(new_n434_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n636_), .B1(new_n637_), .B2(new_n455_), .ZN(new_n638_));
  OAI211_X1 g437(.A(new_n632_), .B(new_n604_), .C1(new_n638_), .C2(new_n435_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(KEYINPUT107), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n629_), .A2(new_n630_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT107), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n641_), .A2(new_n642_), .A3(new_n632_), .A4(new_n604_), .ZN(new_n643_));
  AOI22_X1  g442(.A1(new_n633_), .A2(new_n635_), .B1(new_n640_), .B2(new_n643_), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n551_), .A2(new_n572_), .A3(new_n593_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n625_), .B1(new_n644_), .B2(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n604_), .B1(new_n638_), .B2(new_n435_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n634_), .B1(new_n648_), .B2(KEYINPUT43), .ZN(new_n649_));
  INV_X1    g448(.A(new_n635_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n642_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n651_));
  NOR4_X1   g450(.A1(new_n461_), .A2(KEYINPUT107), .A3(new_n628_), .A4(KEYINPUT43), .ZN(new_n652_));
  OAI22_X1  g451(.A1(new_n649_), .A2(new_n650_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n653_), .A2(KEYINPUT44), .A3(new_n645_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n647_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(G29gat), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n597_), .A2(new_n656_), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n600_), .A2(new_n518_), .A3(new_n573_), .A4(new_n550_), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n658_), .A2(new_n597_), .ZN(new_n659_));
  AOI22_X1  g458(.A1(new_n655_), .A2(new_n657_), .B1(new_n656_), .B2(new_n659_), .ZN(G1328gat));
  OR2_X1    g459(.A1(new_n434_), .A2(G36gat), .ZN(new_n661_));
  OR3_X1    g460(.A1(new_n658_), .A2(KEYINPUT110), .A3(new_n661_), .ZN(new_n662_));
  OAI21_X1  g461(.A(KEYINPUT110), .B1(new_n658_), .B2(new_n661_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT45), .ZN(new_n665_));
  INV_X1    g464(.A(new_n434_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n647_), .A2(new_n654_), .A3(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT109), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n667_), .A2(new_n668_), .A3(G36gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n668_), .B1(new_n667_), .B2(G36gat), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n665_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT46), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  OAI211_X1 g472(.A(KEYINPUT46), .B(new_n665_), .C1(new_n669_), .C2(new_n670_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(G1329gat));
  INV_X1    g474(.A(G43gat), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n260_), .A2(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n647_), .A2(new_n654_), .A3(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(KEYINPUT111), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT111), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n647_), .A2(new_n654_), .A3(new_n680_), .A4(new_n677_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n676_), .B1(new_n658_), .B2(new_n260_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT112), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(KEYINPUT47), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT47), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n682_), .A2(new_n687_), .A3(new_n684_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n688_), .ZN(G1330gat));
  INV_X1    g488(.A(new_n373_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n655_), .A2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(G50gat), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n373_), .A2(G50gat), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT113), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n692_), .B1(new_n658_), .B2(new_n694_), .ZN(G1331gat));
  INV_X1    g494(.A(new_n593_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n461_), .A2(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT114), .ZN(new_n698_));
  NOR4_X1   g497(.A1(new_n698_), .A2(new_n573_), .A3(new_n550_), .A4(new_n604_), .ZN(new_n699_));
  INV_X1    g498(.A(G57gat), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n699_), .A2(new_n700_), .A3(new_n314_), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n550_), .A2(new_n573_), .A3(new_n696_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n519_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(G57gat), .B1(new_n704_), .B2(new_n597_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n701_), .A2(new_n705_), .ZN(G1332gat));
  INV_X1    g505(.A(G64gat), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n707_), .B1(new_n703_), .B2(new_n666_), .ZN(new_n708_));
  XOR2_X1   g507(.A(new_n708_), .B(KEYINPUT48), .Z(new_n709_));
  NAND3_X1  g508(.A1(new_n699_), .A2(new_n707_), .A3(new_n666_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1333gat));
  AOI21_X1  g510(.A(new_n247_), .B1(new_n703_), .B2(new_n636_), .ZN(new_n712_));
  XOR2_X1   g511(.A(new_n712_), .B(KEYINPUT49), .Z(new_n713_));
  NAND3_X1  g512(.A1(new_n699_), .A2(new_n247_), .A3(new_n636_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(G1334gat));
  INV_X1    g514(.A(G78gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n716_), .B1(new_n703_), .B2(new_n690_), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT50), .Z(new_n718_));
  NAND3_X1  g517(.A1(new_n699_), .A2(new_n716_), .A3(new_n690_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n720_), .B(KEYINPUT115), .Z(G1335gat));
  NOR4_X1   g520(.A1(new_n698_), .A2(new_n517_), .A3(new_n572_), .A4(new_n550_), .ZN(new_n722_));
  AOI21_X1  g521(.A(G85gat), .B1(new_n722_), .B2(new_n314_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n551_), .A2(new_n573_), .A3(new_n593_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n644_), .A2(new_n724_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n597_), .A2(new_n485_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n723_), .B1(new_n725_), .B2(new_n726_), .ZN(G1336gat));
  AOI21_X1  g526(.A(G92gat), .B1(new_n722_), .B2(new_n666_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n666_), .A2(G92gat), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT116), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n728_), .B1(new_n725_), .B2(new_n730_), .ZN(G1337gat));
  NAND2_X1  g530(.A1(new_n725_), .A2(new_n636_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n636_), .A2(new_n481_), .ZN(new_n733_));
  AOI22_X1  g532(.A1(new_n732_), .A2(G99gat), .B1(new_n722_), .B2(new_n733_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g534(.A1(new_n722_), .A2(new_n690_), .A3(new_n482_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n725_), .A2(new_n690_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(KEYINPUT117), .A2(KEYINPUT52), .ZN(new_n738_));
  INV_X1    g537(.A(G106gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n739_), .B1(KEYINPUT117), .B2(KEYINPUT52), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n737_), .A2(new_n738_), .A3(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n738_), .B1(new_n737_), .B2(new_n740_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n736_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g543(.A(KEYINPUT58), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n532_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT55), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n538_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n536_), .A2(new_n537_), .A3(KEYINPUT55), .A4(new_n532_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n546_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n583_), .A2(new_n588_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n576_), .A2(new_n580_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n579_), .A2(new_n577_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n754_), .A2(new_n587_), .A3(new_n755_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n753_), .A2(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n752_), .A2(new_n547_), .A3(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT56), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n750_), .A2(KEYINPUT119), .A3(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n745_), .B1(new_n758_), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT120), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n761_), .A2(new_n762_), .A3(new_n604_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n757_), .A2(new_n547_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n764_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n748_), .A2(new_n749_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(new_n544_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT119), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n767_), .A2(new_n768_), .A3(KEYINPUT56), .ZN(new_n769_));
  AOI21_X1  g568(.A(KEYINPUT58), .B1(new_n765_), .B2(new_n769_), .ZN(new_n770_));
  OAI21_X1  g569(.A(KEYINPUT120), .B1(new_n770_), .B2(new_n628_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n765_), .A2(new_n769_), .A3(KEYINPUT58), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n763_), .A2(new_n771_), .A3(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT57), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT121), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n591_), .A2(new_n592_), .A3(new_n547_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT118), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n767_), .A2(new_n777_), .A3(new_n759_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n750_), .B1(KEYINPUT118), .B2(KEYINPUT56), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n776_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n757_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n781_), .B1(new_n545_), .B2(new_n547_), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n517_), .B(new_n775_), .C1(new_n780_), .C2(new_n782_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n774_), .A2(KEYINPUT121), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n785_), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n517_), .B(new_n784_), .C1(new_n780_), .C2(new_n782_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n773_), .A2(new_n786_), .A3(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n605_), .A2(new_n550_), .ZN(new_n789_));
  OR3_X1    g588(.A1(new_n789_), .A2(KEYINPUT54), .A3(new_n696_), .ZN(new_n790_));
  OAI21_X1  g589(.A(KEYINPUT54), .B1(new_n789_), .B2(new_n696_), .ZN(new_n791_));
  AOI22_X1  g590(.A1(new_n788_), .A2(new_n573_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n666_), .A2(new_n690_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n793_), .A2(new_n314_), .A3(new_n636_), .ZN(new_n794_));
  XOR2_X1   g593(.A(KEYINPUT123), .B(KEYINPUT59), .Z(new_n795_));
  OR3_X1    g594(.A1(new_n792_), .A2(new_n794_), .A3(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT122), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n788_), .A2(new_n797_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n773_), .A2(new_n786_), .A3(KEYINPUT122), .A4(new_n787_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n798_), .A2(new_n573_), .A3(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n790_), .A2(new_n791_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n794_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT59), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n796_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(G113gat), .B1(new_n804_), .B2(new_n593_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n802_), .ZN(new_n806_));
  OR2_X1    g605(.A1(new_n593_), .A2(G113gat), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n805_), .B1(new_n806_), .B2(new_n807_), .ZN(G1340gat));
  OAI21_X1  g607(.A(G120gat), .B1(new_n804_), .B2(new_n550_), .ZN(new_n809_));
  INV_X1    g608(.A(G120gat), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n810_), .B1(new_n550_), .B2(KEYINPUT60), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n811_), .B1(KEYINPUT60), .B2(new_n810_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n809_), .B1(new_n806_), .B2(new_n812_), .ZN(G1341gat));
  OAI21_X1  g612(.A(G127gat), .B1(new_n804_), .B2(new_n573_), .ZN(new_n814_));
  OR2_X1    g613(.A1(new_n573_), .A2(G127gat), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n814_), .B1(new_n806_), .B2(new_n815_), .ZN(G1342gat));
  XNOR2_X1  g615(.A(KEYINPUT124), .B(G134gat), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n604_), .A2(new_n817_), .ZN(new_n818_));
  OR2_X1    g617(.A1(new_n804_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(G134gat), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n820_), .B1(new_n806_), .B2(new_n517_), .ZN(new_n821_));
  AND2_X1   g620(.A1(new_n819_), .A2(new_n821_), .ZN(G1343gat));
  NOR3_X1   g621(.A1(new_n666_), .A2(new_n597_), .A3(new_n373_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  AOI211_X1 g623(.A(new_n636_), .B(new_n824_), .C1(new_n800_), .C2(new_n801_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n696_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n826_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g626(.A1(new_n825_), .A2(new_n551_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n828_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g628(.A(KEYINPUT125), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n825_), .A2(new_n830_), .A3(new_n572_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n800_), .A2(new_n801_), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n832_), .A2(new_n260_), .A3(new_n572_), .A4(new_n823_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(KEYINPUT125), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n831_), .A2(new_n834_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(KEYINPUT61), .B(G155gat), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n835_), .A2(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n831_), .A2(new_n834_), .A3(new_n836_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(G1346gat));
  INV_X1    g639(.A(G162gat), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n825_), .A2(new_n841_), .A3(new_n518_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n832_), .A2(new_n260_), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n843_), .A2(new_n628_), .A3(new_n824_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n842_), .B1(new_n844_), .B2(new_n841_), .ZN(G1347gat));
  NAND2_X1  g644(.A1(new_n666_), .A2(new_n315_), .ZN(new_n846_));
  NOR3_X1   g645(.A1(new_n792_), .A2(new_n690_), .A3(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n696_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n848_), .A2(new_n402_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n221_), .B1(new_n847_), .B2(new_n696_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n849_), .B1(KEYINPUT62), .B2(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n851_), .B1(KEYINPUT62), .B2(new_n850_), .ZN(G1348gat));
  AOI21_X1  g651(.A(new_n690_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n846_), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n853_), .A2(G176gat), .A3(new_n551_), .A4(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n847_), .A2(new_n551_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n855_), .B1(new_n857_), .B2(G176gat), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT126), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n855_), .B(KEYINPUT126), .C1(new_n857_), .C2(G176gat), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(G1349gat));
  NAND3_X1  g661(.A1(new_n853_), .A2(new_n572_), .A3(new_n854_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n573_), .A2(new_n236_), .ZN(new_n864_));
  AOI22_X1  g663(.A1(new_n863_), .A2(new_n206_), .B1(new_n847_), .B2(new_n864_), .ZN(G1350gat));
  NAND4_X1  g664(.A1(new_n847_), .A2(new_n387_), .A3(new_n388_), .A4(new_n518_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n847_), .A2(new_n604_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n866_), .B1(new_n867_), .B2(new_n207_), .ZN(G1351gat));
  NAND2_X1  g667(.A1(new_n666_), .A2(new_n458_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n843_), .A2(new_n593_), .A3(new_n869_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(new_n319_), .ZN(G1352gat));
  NOR3_X1   g670(.A1(new_n843_), .A2(new_n550_), .A3(new_n869_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(new_n316_), .ZN(G1353gat));
  NOR2_X1   g672(.A1(new_n843_), .A2(new_n869_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n573_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(KEYINPUT127), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n876_), .A2(new_n879_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n874_), .A2(new_n878_), .A3(new_n875_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(G1354gat));
  INV_X1    g681(.A(G218gat), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n874_), .A2(new_n883_), .A3(new_n518_), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n843_), .A2(new_n628_), .A3(new_n869_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n885_), .B2(new_n883_), .ZN(G1355gat));
endmodule


