//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 1 1 0 1 0 1 0 0 0 1 0 0 1 1 1 0 0 0 0 1 1 0 0 0 1 0 1 1 1 1 1 1 0 0 1 1 1 1 1 0 1 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n634_, new_n635_,
    new_n636_, new_n638_, new_n639_, new_n640_, new_n641_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n726_, new_n727_, new_n728_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n762_, new_n763_, new_n765_, new_n766_, new_n767_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n838_, new_n839_, new_n840_, new_n841_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n848_, new_n849_, new_n850_,
    new_n852_, new_n853_, new_n854_, new_n856_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n901_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_;
  XNOR2_X1  g000(.A(G22gat), .B(G50gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G78gat), .B(G106gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G228gat), .A2(G233gat), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(G141gat), .ZN(new_n208_));
  INV_X1    g007(.A(G148gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G141gat), .A2(G148gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n212_));
  AND3_X1   g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G155gat), .B(G162gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n213_), .B1(KEYINPUT1), .B2(new_n214_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT84), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n208_), .A2(new_n209_), .A3(KEYINPUT3), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT3), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n219_), .B1(G141gat), .B2(G148gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT2), .ZN(new_n221_));
  AOI22_X1  g020(.A1(new_n218_), .A2(new_n220_), .B1(new_n221_), .B2(new_n211_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n214_), .B1(new_n217_), .B2(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n215_), .B1(new_n223_), .B2(KEYINPUT85), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT85), .ZN(new_n225_));
  AOI211_X1 g024(.A(new_n225_), .B(new_n214_), .C1(new_n217_), .C2(new_n222_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT29), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(G197gat), .A2(G204gat), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT87), .B(G197gat), .ZN(new_n232_));
  INV_X1    g031(.A(G204gat), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n231_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT21), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G211gat), .B(G218gat), .ZN(new_n236_));
  NOR3_X1   g035(.A1(new_n234_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(G197gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT87), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT87), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(G197gat), .ZN(new_n241_));
  AOI21_X1  g040(.A(G204gat), .B1(new_n239_), .B2(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT88), .B1(new_n233_), .B2(G197gat), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT88), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n244_), .A2(new_n238_), .A3(G204gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT21), .B1(new_n242_), .B2(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n233_), .B1(new_n239_), .B2(new_n241_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n235_), .B1(new_n248_), .B2(new_n230_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n247_), .A2(new_n249_), .A3(new_n236_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT89), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n236_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n253_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n254_), .A2(KEYINPUT89), .A3(new_n247_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n237_), .B1(new_n252_), .B2(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n207_), .B1(new_n229_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT86), .ZN(new_n258_));
  INV_X1    g057(.A(new_n237_), .ZN(new_n259_));
  AOI21_X1  g058(.A(KEYINPUT89), .B1(new_n254_), .B2(new_n247_), .ZN(new_n260_));
  AND4_X1   g059(.A1(KEYINPUT89), .A2(new_n247_), .A3(new_n249_), .A4(new_n236_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n259_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n262_), .B(new_n206_), .C1(new_n228_), .C2(new_n227_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n257_), .A2(new_n258_), .A3(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT90), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n227_), .A2(new_n228_), .ZN(new_n266_));
  XOR2_X1   g065(.A(new_n266_), .B(KEYINPUT28), .Z(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT90), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n257_), .A2(new_n258_), .A3(new_n263_), .A4(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n265_), .A2(new_n268_), .A3(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n268_), .B1(new_n265_), .B2(new_n270_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n203_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n265_), .A2(new_n270_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(new_n267_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n276_), .A2(new_n202_), .A3(new_n271_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n274_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT97), .ZN(new_n280_));
  AND2_X1   g079(.A1(KEYINPUT78), .A2(G169gat), .ZN(new_n281_));
  NOR2_X1   g080(.A1(KEYINPUT78), .A2(G169gat), .ZN(new_n282_));
  OAI21_X1  g081(.A(KEYINPUT22), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT79), .ZN(new_n284_));
  XNOR2_X1  g083(.A(KEYINPUT80), .B(G176gat), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT22), .ZN(new_n286_));
  AND2_X1   g085(.A1(new_n286_), .A2(G169gat), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT79), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n289_), .B(KEYINPUT22), .C1(new_n281_), .C2(new_n282_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n284_), .A2(new_n288_), .A3(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(G183gat), .ZN(new_n292_));
  INV_X1    g091(.A(G190gat), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT23), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT23), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n295_), .A2(G183gat), .A3(G190gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n292_), .A2(new_n293_), .ZN(new_n298_));
  AOI22_X1  g097(.A1(new_n297_), .A2(new_n298_), .B1(G169gat), .B2(G176gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n293_), .A2(KEYINPUT26), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT26), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(G190gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n292_), .A2(KEYINPUT25), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT25), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(G183gat), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n300_), .A2(new_n302_), .A3(new_n303_), .A4(new_n305_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(G169gat), .A2(G176gat), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G169gat), .A2(G176gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n308_), .A2(KEYINPUT24), .A3(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT24), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n307_), .A2(new_n311_), .ZN(new_n312_));
  AND3_X1   g111(.A1(new_n306_), .A2(new_n310_), .A3(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT77), .ZN(new_n314_));
  AND2_X1   g113(.A1(new_n296_), .A2(new_n314_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n296_), .A2(new_n314_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n294_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  AOI22_X1  g116(.A1(new_n291_), .A2(new_n299_), .B1(new_n313_), .B2(new_n317_), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n259_), .B(new_n318_), .C1(new_n260_), .C2(new_n261_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(new_n298_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n288_), .B1(new_n286_), .B2(G169gat), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n320_), .A2(new_n309_), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n303_), .A2(new_n305_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT91), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT91), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n303_), .A2(new_n305_), .A3(new_n325_), .ZN(new_n326_));
  AND2_X1   g125(.A1(new_n300_), .A2(new_n302_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n324_), .A2(new_n326_), .A3(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n309_), .A2(KEYINPUT24), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT92), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n307_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n331_), .B1(new_n330_), .B2(new_n329_), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n328_), .A2(new_n332_), .A3(new_n297_), .A4(new_n312_), .ZN(new_n333_));
  AND2_X1   g132(.A1(new_n322_), .A2(new_n333_), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n319_), .B(KEYINPUT20), .C1(new_n256_), .C2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G226gat), .A2(G233gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT19), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n280_), .B1(new_n335_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT20), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n339_), .B1(new_n256_), .B2(new_n318_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n322_), .A2(new_n333_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n262_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n337_), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n340_), .A2(KEYINPUT97), .A3(new_n342_), .A4(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(KEYINPUT20), .B1(new_n262_), .B2(new_n341_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT93), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n346_), .B1(new_n256_), .B2(new_n318_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n318_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n262_), .A2(KEYINPUT93), .A3(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n345_), .B1(new_n347_), .B2(new_n349_), .ZN(new_n350_));
  OAI211_X1 g149(.A(new_n338_), .B(new_n344_), .C1(new_n350_), .C2(new_n343_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G8gat), .B(G36gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT18), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G64gat), .B(G92gat), .ZN(new_n354_));
  XOR2_X1   g153(.A(new_n353_), .B(new_n354_), .Z(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n351_), .A2(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n339_), .B1(new_n334_), .B2(new_n256_), .ZN(new_n358_));
  NOR3_X1   g157(.A1(new_n256_), .A2(new_n346_), .A3(new_n318_), .ZN(new_n359_));
  AOI21_X1  g158(.A(KEYINPUT93), .B1(new_n262_), .B2(new_n348_), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n343_), .B(new_n358_), .C1(new_n359_), .C2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n335_), .A2(new_n337_), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n361_), .A2(KEYINPUT99), .A3(new_n355_), .A4(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n361_), .A2(new_n355_), .A3(new_n362_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT99), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n357_), .A2(new_n363_), .A3(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT27), .ZN(new_n368_));
  INV_X1    g167(.A(new_n364_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n355_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n370_));
  OR3_X1    g169(.A1(new_n369_), .A2(KEYINPUT27), .A3(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n368_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G225gat), .A2(G233gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G127gat), .B(G134gat), .ZN(new_n374_));
  OR2_X1    g173(.A1(new_n374_), .A2(KEYINPUT81), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(KEYINPUT81), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G113gat), .B(G120gat), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n375_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n377_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n374_), .A2(KEYINPUT81), .ZN(new_n380_));
  INV_X1    g179(.A(G134gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(G127gat), .ZN(new_n382_));
  INV_X1    g181(.A(G127gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(G134gat), .ZN(new_n384_));
  AND3_X1   g183(.A1(new_n382_), .A2(new_n384_), .A3(KEYINPUT81), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n379_), .B1(new_n380_), .B2(new_n385_), .ZN(new_n386_));
  AND2_X1   g185(.A1(new_n378_), .A2(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n387_), .B1(new_n224_), .B2(new_n226_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n218_), .A2(new_n220_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n211_), .A2(new_n221_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT84), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n216_), .B(new_n392_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n391_), .A2(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n225_), .B1(new_n394_), .B2(new_n214_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n378_), .A2(new_n386_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n223_), .A2(KEYINPUT85), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n395_), .A2(new_n396_), .A3(new_n397_), .A4(new_n215_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n388_), .A2(KEYINPUT4), .A3(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT4), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n387_), .B(new_n400_), .C1(new_n224_), .C2(new_n226_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n373_), .B1(new_n399_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n388_), .A2(new_n398_), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n404_), .A2(new_n373_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G1gat), .B(G29gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(G85gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(KEYINPUT0), .B(G57gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n408_), .B(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n403_), .A2(new_n406_), .A3(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n410_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n412_), .B1(new_n402_), .B2(new_n405_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n411_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G71gat), .B(G99gat), .ZN(new_n416_));
  INV_X1    g215(.A(G43gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n318_), .B(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G227gat), .A2(G233gat), .ZN(new_n420_));
  INV_X1    g219(.A(G15gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(KEYINPUT30), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n419_), .B(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n396_), .B(KEYINPUT31), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT83), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n426_), .B(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n424_), .A2(new_n425_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT82), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n429_), .B(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n428_), .A2(new_n431_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n279_), .A2(new_n372_), .A3(new_n415_), .A4(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n355_), .A2(KEYINPUT32), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n361_), .A2(new_n362_), .A3(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT96), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n361_), .A2(KEYINPUT96), .A3(new_n362_), .A4(new_n435_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n435_), .ZN(new_n441_));
  AOI22_X1  g240(.A1(new_n351_), .A2(new_n441_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n440_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT98), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n440_), .A2(new_n442_), .A3(KEYINPUT98), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT94), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n447_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n361_), .A2(new_n362_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(new_n356_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n450_), .A2(KEYINPUT94), .A3(new_n364_), .ZN(new_n451_));
  OAI211_X1 g250(.A(KEYINPUT33), .B(new_n412_), .C1(new_n402_), .C2(new_n405_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n373_), .B1(new_n404_), .B2(KEYINPUT95), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT95), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n388_), .A2(new_n454_), .A3(new_n398_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n399_), .A2(new_n373_), .A3(new_n401_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(new_n410_), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT33), .B1(new_n457_), .B2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(new_n413_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n448_), .A2(new_n451_), .A3(new_n452_), .A4(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n445_), .A2(new_n446_), .A3(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n279_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n414_), .B1(new_n274_), .B2(new_n277_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(new_n372_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n432_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n434_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G1gat), .B(G8gat), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT72), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n470_), .B(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT73), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT71), .B(G15gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(G22gat), .ZN(new_n476_));
  INV_X1    g275(.A(G1gat), .ZN(new_n477_));
  INV_X1    g276(.A(G8gat), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT14), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n476_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n474_), .A2(new_n480_), .ZN(new_n481_));
  OR2_X1    g280(.A1(new_n472_), .A2(new_n473_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n472_), .A2(new_n473_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n482_), .A2(new_n479_), .A3(new_n476_), .A4(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n481_), .A2(new_n484_), .ZN(new_n485_));
  XOR2_X1   g284(.A(G29gat), .B(G36gat), .Z(new_n486_));
  XOR2_X1   g285(.A(G43gat), .B(G50gat), .Z(new_n487_));
  XOR2_X1   g286(.A(new_n486_), .B(new_n487_), .Z(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n485_), .B(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n490_), .A2(G229gat), .A3(G233gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n488_), .B(KEYINPUT15), .ZN(new_n492_));
  OR2_X1    g291(.A1(new_n485_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G229gat), .A2(G233gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n485_), .A2(new_n489_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n493_), .A2(new_n494_), .A3(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n491_), .A2(new_n496_), .ZN(new_n497_));
  XOR2_X1   g296(.A(G113gat), .B(G141gat), .Z(new_n498_));
  XNOR2_X1  g297(.A(G169gat), .B(G197gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n497_), .B(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G85gat), .B(G92gat), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT64), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n502_), .B1(new_n503_), .B2(KEYINPUT8), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G99gat), .A2(G106gat), .ZN(new_n505_));
  XOR2_X1   g304(.A(new_n505_), .B(KEYINPUT6), .Z(new_n506_));
  NOR2_X1   g305(.A1(G99gat), .A2(G106gat), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT7), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n504_), .B1(new_n506_), .B2(new_n509_), .ZN(new_n510_));
  OR2_X1    g309(.A1(new_n503_), .A2(KEYINPUT8), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(G85gat), .ZN(new_n513_));
  INV_X1    g312(.A(G92gat), .ZN(new_n514_));
  NOR3_X1   g313(.A1(new_n513_), .A2(new_n514_), .A3(KEYINPUT9), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n506_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT9), .ZN(new_n517_));
  XOR2_X1   g316(.A(KEYINPUT10), .B(G99gat), .Z(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  OAI221_X1 g318(.A(new_n516_), .B1(new_n517_), .B2(new_n502_), .C1(G106gat), .C2(new_n519_), .ZN(new_n520_));
  AND2_X1   g319(.A1(new_n512_), .A2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G57gat), .B(G64gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT11), .ZN(new_n523_));
  XOR2_X1   g322(.A(G71gat), .B(G78gat), .Z(new_n524_));
  OR2_X1    g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n522_), .A2(KEYINPUT11), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n523_), .A2(new_n524_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n525_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n521_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  OAI21_X1  g329(.A(KEYINPUT65), .B1(new_n521_), .B2(new_n528_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n530_), .B1(new_n531_), .B2(KEYINPUT12), .ZN(new_n532_));
  OR2_X1    g331(.A1(new_n531_), .A2(KEYINPUT12), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G230gat), .A2(G233gat), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n532_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n521_), .A2(new_n528_), .ZN(new_n536_));
  OAI211_X1 g335(.A(G230gat), .B(G233gat), .C1(new_n530_), .C2(new_n536_), .ZN(new_n537_));
  XOR2_X1   g336(.A(G120gat), .B(G148gat), .Z(new_n538_));
  XNOR2_X1  g337(.A(G176gat), .B(G204gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n535_), .A2(new_n537_), .A3(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n535_), .A2(new_n537_), .ZN(new_n546_));
  OR2_X1    g345(.A1(new_n546_), .A2(KEYINPUT66), .ZN(new_n547_));
  XOR2_X1   g346(.A(new_n542_), .B(KEYINPUT68), .Z(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n549_), .B1(new_n546_), .B2(KEYINPUT66), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n545_), .B1(new_n547_), .B2(new_n550_), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n551_), .A2(KEYINPUT13), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(KEYINPUT13), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NOR3_X1   g353(.A1(new_n469_), .A2(new_n501_), .A3(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n521_), .A2(new_n488_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n512_), .A2(new_n520_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(new_n492_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n556_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G232gat), .A2(G233gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT34), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n561_), .A2(KEYINPUT35), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(KEYINPUT35), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n559_), .A2(KEYINPUT70), .A3(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n556_), .A2(new_n558_), .A3(new_n562_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(KEYINPUT70), .B1(new_n559_), .B2(new_n564_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT36), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G190gat), .B(G218gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT69), .ZN(new_n572_));
  XOR2_X1   g371(.A(G134gat), .B(G162gat), .Z(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n569_), .A2(new_n570_), .A3(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n570_), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n574_), .A2(new_n570_), .ZN(new_n577_));
  OAI211_X1 g376(.A(new_n576_), .B(new_n577_), .C1(new_n567_), .C2(new_n568_), .ZN(new_n578_));
  AOI21_X1  g377(.A(KEYINPUT37), .B1(new_n575_), .B2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n575_), .A2(new_n578_), .A3(KEYINPUT37), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G231gat), .A2(G233gat), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n528_), .B(new_n583_), .Z(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(new_n485_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  XOR2_X1   g385(.A(G127gat), .B(G155gat), .Z(new_n587_));
  XNOR2_X1  g386(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G183gat), .B(G211gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n591_), .A2(KEYINPUT17), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n591_), .A2(KEYINPUT17), .ZN(new_n593_));
  NOR3_X1   g392(.A1(new_n586_), .A2(new_n592_), .A3(new_n593_), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n594_), .B(KEYINPUT76), .Z(new_n595_));
  OR2_X1    g394(.A1(new_n585_), .A2(KEYINPUT74), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n585_), .A2(KEYINPUT74), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n596_), .A2(new_n593_), .A3(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n595_), .A2(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n582_), .A2(new_n599_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n555_), .A2(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n601_), .A2(new_n477_), .A3(new_n414_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT38), .ZN(new_n603_));
  INV_X1    g402(.A(new_n501_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n599_), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n552_), .A2(new_n604_), .A3(new_n553_), .A4(new_n605_), .ZN(new_n606_));
  OR2_X1    g405(.A1(new_n606_), .A2(KEYINPUT100), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n575_), .A2(new_n578_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT101), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n469_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n606_), .A2(KEYINPUT100), .ZN(new_n612_));
  AND3_X1   g411(.A1(new_n607_), .A2(new_n611_), .A3(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT102), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n614_), .A2(new_n414_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n603_), .B1(new_n615_), .B2(new_n477_), .ZN(G1324gat));
  XNOR2_X1  g415(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n617_));
  INV_X1    g416(.A(new_n372_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n613_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT103), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(G8gat), .B1(new_n619_), .B2(KEYINPUT103), .ZN(new_n623_));
  OR3_X1    g422(.A1(new_n622_), .A2(KEYINPUT39), .A3(new_n623_), .ZN(new_n624_));
  OAI21_X1  g423(.A(KEYINPUT39), .B1(new_n622_), .B2(new_n623_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n372_), .A2(G8gat), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n601_), .A2(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n617_), .B1(new_n626_), .B2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n628_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n617_), .ZN(new_n631_));
  AOI211_X1 g430(.A(new_n630_), .B(new_n631_), .C1(new_n624_), .C2(new_n625_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n629_), .A2(new_n632_), .ZN(G1325gat));
  AOI21_X1  g432(.A(new_n421_), .B1(new_n614_), .B2(new_n432_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT41), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n601_), .A2(new_n421_), .A3(new_n432_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(G1326gat));
  INV_X1    g436(.A(G22gat), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n638_), .B1(new_n614_), .B2(new_n278_), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n639_), .B(KEYINPUT42), .Z(new_n640_));
  NAND3_X1  g439(.A1(new_n601_), .A2(new_n638_), .A3(new_n278_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(G1327gat));
  NOR2_X1   g441(.A1(new_n605_), .A2(new_n608_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n555_), .A2(new_n643_), .ZN(new_n644_));
  OR3_X1    g443(.A1(new_n644_), .A2(G29gat), .A3(new_n415_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT44), .ZN(new_n646_));
  AOI22_X1  g445(.A1(new_n463_), .A2(new_n279_), .B1(new_n465_), .B2(new_n372_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n433_), .B1(new_n647_), .B2(new_n432_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT43), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n648_), .A2(new_n649_), .A3(new_n582_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT106), .ZN(new_n652_));
  INV_X1    g451(.A(new_n581_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n652_), .B1(new_n653_), .B2(new_n579_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n580_), .A2(KEYINPUT106), .A3(new_n581_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(KEYINPUT94), .B1(new_n450_), .B2(new_n364_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT33), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n458_), .A2(new_n410_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n658_), .B1(new_n659_), .B2(new_n456_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n413_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n452_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n657_), .A2(new_n662_), .ZN(new_n663_));
  AOI22_X1  g462(.A1(new_n663_), .A2(new_n451_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n278_), .B1(new_n664_), .B2(new_n446_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n465_), .A2(new_n372_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n468_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n656_), .B1(new_n667_), .B2(new_n433_), .ZN(new_n668_));
  OAI21_X1  g467(.A(KEYINPUT107), .B1(new_n668_), .B2(new_n649_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n654_), .A2(new_n655_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n648_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT107), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n671_), .A2(new_n672_), .A3(KEYINPUT43), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n651_), .B1(new_n669_), .B2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT13), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n551_), .B(new_n675_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n676_), .A2(new_n604_), .A3(new_n599_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT105), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n646_), .B1(new_n674_), .B2(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n672_), .B1(new_n671_), .B2(KEYINPUT43), .ZN(new_n680_));
  AOI211_X1 g479(.A(KEYINPUT107), .B(new_n649_), .C1(new_n648_), .C2(new_n670_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n650_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  XOR2_X1   g481(.A(new_n677_), .B(KEYINPUT105), .Z(new_n683_));
  NAND3_X1  g482(.A1(new_n682_), .A2(KEYINPUT44), .A3(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n679_), .A2(new_n414_), .A3(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT108), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  OAI21_X1  g486(.A(G29gat), .B1(new_n685_), .B2(new_n686_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n645_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(KEYINPUT109), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT109), .ZN(new_n691_));
  OAI211_X1 g490(.A(new_n691_), .B(new_n645_), .C1(new_n687_), .C2(new_n688_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n690_), .A2(new_n692_), .ZN(G1328gat));
  INV_X1    g492(.A(KEYINPUT46), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT45), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n554_), .A2(new_n501_), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n372_), .A2(KEYINPUT110), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n372_), .A2(KEYINPUT110), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n699_), .A2(G36gat), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n696_), .A2(new_n700_), .A3(new_n648_), .A4(new_n643_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(KEYINPUT111), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n701_), .A2(KEYINPUT111), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n695_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n704_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n706_), .A2(KEYINPUT45), .A3(new_n702_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n679_), .A2(new_n618_), .A3(new_n684_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n708_), .B1(new_n709_), .B2(G36gat), .ZN(new_n710_));
  OAI211_X1 g509(.A(KEYINPUT113), .B(new_n694_), .C1(new_n710_), .C2(KEYINPUT112), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT113), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n709_), .A2(G36gat), .ZN(new_n713_));
  INV_X1    g512(.A(new_n708_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT112), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n712_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(KEYINPUT46), .B1(new_n710_), .B2(KEYINPUT113), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n711_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(G1329gat));
  AND2_X1   g519(.A1(new_n679_), .A2(new_n684_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n721_), .A2(G43gat), .A3(new_n432_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n417_), .B1(new_n644_), .B2(new_n468_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g524(.A1(new_n721_), .A2(G50gat), .A3(new_n278_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n644_), .A2(new_n279_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n726_), .B1(G50gat), .B2(new_n727_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT114), .ZN(G1331gat));
  NOR3_X1   g528(.A1(new_n469_), .A2(new_n604_), .A3(new_n676_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n730_), .A2(new_n600_), .ZN(new_n731_));
  INV_X1    g530(.A(G57gat), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n731_), .A2(new_n732_), .A3(new_n414_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n599_), .A2(new_n604_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n611_), .A2(new_n554_), .A3(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT115), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n736_), .A2(new_n414_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n733_), .B1(new_n737_), .B2(new_n732_), .ZN(G1332gat));
  INV_X1    g537(.A(G64gat), .ZN(new_n739_));
  INV_X1    g538(.A(new_n699_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n736_), .B2(new_n740_), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n741_), .B(KEYINPUT48), .Z(new_n742_));
  NAND3_X1  g541(.A1(new_n731_), .A2(new_n739_), .A3(new_n740_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(G1333gat));
  INV_X1    g543(.A(G71gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n736_), .B2(new_n432_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT49), .Z(new_n747_));
  NAND3_X1  g546(.A1(new_n731_), .A2(new_n745_), .A3(new_n432_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(G1334gat));
  INV_X1    g548(.A(G78gat), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n750_), .B1(new_n736_), .B2(new_n278_), .ZN(new_n751_));
  XOR2_X1   g550(.A(new_n751_), .B(KEYINPUT50), .Z(new_n752_));
  NAND3_X1  g551(.A1(new_n731_), .A2(new_n750_), .A3(new_n278_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(G1335gat));
  NAND2_X1  g553(.A1(new_n730_), .A2(new_n643_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n513_), .B1(new_n755_), .B2(new_n415_), .ZN(new_n756_));
  XOR2_X1   g555(.A(new_n756_), .B(KEYINPUT116), .Z(new_n757_));
  NAND3_X1  g556(.A1(new_n554_), .A2(new_n501_), .A3(new_n599_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n674_), .A2(new_n758_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n415_), .A2(new_n513_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n757_), .B1(new_n759_), .B2(new_n760_), .ZN(G1336gat));
  NOR3_X1   g560(.A1(new_n674_), .A2(new_n699_), .A3(new_n758_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n618_), .A2(new_n514_), .ZN(new_n763_));
  OAI22_X1  g562(.A1(new_n762_), .A2(new_n514_), .B1(new_n755_), .B2(new_n763_), .ZN(G1337gat));
  NOR3_X1   g563(.A1(new_n755_), .A2(new_n468_), .A3(new_n519_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n759_), .A2(new_n432_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n765_), .B1(new_n766_), .B2(G99gat), .ZN(new_n767_));
  XOR2_X1   g566(.A(new_n767_), .B(KEYINPUT51), .Z(G1338gat));
  OR3_X1    g567(.A1(new_n755_), .A2(G106gat), .A3(new_n279_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n759_), .A2(new_n278_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT52), .ZN(new_n771_));
  AND3_X1   g570(.A1(new_n770_), .A2(new_n771_), .A3(G106gat), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n771_), .B1(new_n770_), .B2(G106gat), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n769_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g574(.A(KEYINPUT120), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n493_), .A2(new_n495_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n494_), .B1(new_n777_), .B2(KEYINPUT119), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n778_), .B1(KEYINPUT119), .B2(new_n777_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n500_), .B1(new_n490_), .B2(new_n494_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n491_), .A2(new_n496_), .A3(new_n500_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  OR3_X1    g582(.A1(new_n551_), .A2(new_n776_), .A3(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n534_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT55), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n535_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n532_), .A2(new_n533_), .A3(KEYINPUT55), .A4(new_n534_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n789_), .A2(KEYINPUT56), .A3(new_n548_), .ZN(new_n790_));
  AOI21_X1  g589(.A(KEYINPUT56), .B1(new_n789_), .B2(new_n548_), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n604_), .B(new_n544_), .C1(new_n790_), .C2(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n776_), .B1(new_n551_), .B2(new_n783_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n784_), .A2(new_n792_), .A3(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(new_n608_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT121), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n796_), .A2(KEYINPUT57), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT122), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n798_), .B1(new_n783_), .B2(new_n545_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n781_), .A2(KEYINPUT122), .A3(new_n544_), .A4(new_n782_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n801_), .B(KEYINPUT58), .C1(new_n791_), .C2(new_n790_), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n802_), .A2(new_n582_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n801_), .B1(new_n791_), .B2(new_n790_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT58), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  AOI22_X1  g605(.A1(new_n795_), .A2(new_n797_), .B1(new_n803_), .B2(new_n806_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n794_), .B(new_n608_), .C1(new_n796_), .C2(KEYINPUT57), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n605_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n552_), .A2(new_n734_), .A3(new_n553_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT117), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n582_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n676_), .A2(KEYINPUT117), .A3(new_n734_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT118), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT54), .ZN(new_n815_));
  AND3_X1   g614(.A1(new_n812_), .A2(new_n813_), .A3(new_n815_), .ZN(new_n816_));
  OR2_X1    g615(.A1(new_n814_), .A2(KEYINPUT54), .ZN(new_n817_));
  AOI22_X1  g616(.A1(new_n812_), .A2(new_n813_), .B1(new_n817_), .B2(new_n815_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n816_), .A2(new_n818_), .ZN(new_n819_));
  OR2_X1    g618(.A1(new_n809_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT59), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n279_), .A2(new_n372_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n432_), .A2(new_n414_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n820_), .A2(new_n821_), .A3(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n824_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n807_), .A2(new_n808_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT123), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n605_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n829_), .B1(new_n828_), .B2(new_n827_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n819_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n826_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n825_), .B1(new_n832_), .B2(new_n821_), .ZN(new_n833_));
  OAI21_X1  g632(.A(G113gat), .B1(new_n833_), .B2(new_n501_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n832_), .ZN(new_n835_));
  OR3_X1    g634(.A1(new_n835_), .A2(G113gat), .A3(new_n501_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n836_), .ZN(G1340gat));
  OAI21_X1  g636(.A(G120gat), .B1(new_n833_), .B2(new_n676_), .ZN(new_n838_));
  INV_X1    g637(.A(G120gat), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n839_), .B1(new_n676_), .B2(KEYINPUT60), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n832_), .B(new_n840_), .C1(KEYINPUT60), .C2(new_n839_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n838_), .A2(new_n841_), .ZN(G1341gat));
  OAI21_X1  g641(.A(new_n383_), .B1(new_n835_), .B2(new_n599_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n599_), .A2(new_n383_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(KEYINPUT124), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n825_), .B(new_n845_), .C1(new_n832_), .C2(new_n821_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n843_), .A2(new_n846_), .ZN(G1342gat));
  INV_X1    g646(.A(new_n582_), .ZN(new_n848_));
  OAI21_X1  g647(.A(G134gat), .B1(new_n833_), .B2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n832_), .A2(new_n381_), .A3(new_n610_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(G1343gat));
  NAND2_X1  g650(.A1(new_n830_), .A2(new_n831_), .ZN(new_n852_));
  NOR4_X1   g651(.A1(new_n740_), .A2(new_n415_), .A3(new_n279_), .A4(new_n432_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n852_), .A2(new_n604_), .A3(new_n853_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g654(.A1(new_n852_), .A2(new_n554_), .A3(new_n853_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g656(.A1(new_n852_), .A2(new_n605_), .A3(new_n853_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(KEYINPUT61), .B(G155gat), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n858_), .B(new_n859_), .ZN(G1346gat));
  AND2_X1   g659(.A1(new_n852_), .A2(new_n853_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n610_), .ZN(new_n862_));
  INV_X1    g661(.A(G162gat), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n656_), .A2(new_n863_), .ZN(new_n864_));
  AOI22_X1  g663(.A1(new_n862_), .A2(new_n863_), .B1(new_n861_), .B2(new_n864_), .ZN(G1347gat));
  NAND2_X1  g664(.A1(new_n432_), .A2(new_n415_), .ZN(new_n866_));
  OR2_X1    g665(.A1(new_n699_), .A2(new_n866_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n867_), .A2(new_n278_), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n604_), .B(new_n868_), .C1(new_n809_), .C2(new_n819_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT125), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n869_), .A2(new_n870_), .A3(G169gat), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n870_), .B1(new_n869_), .B2(G169gat), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT62), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n872_), .A2(new_n873_), .A3(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n874_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n286_), .A2(G169gat), .ZN(new_n877_));
  OR3_X1    g676(.A1(new_n869_), .A2(new_n287_), .A3(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n878_), .ZN(new_n879_));
  OAI21_X1  g678(.A(KEYINPUT126), .B1(new_n875_), .B2(new_n879_), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n869_), .A2(new_n287_), .A3(new_n877_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n881_), .B1(new_n874_), .B2(new_n873_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT126), .ZN(new_n883_));
  OR2_X1    g682(.A1(new_n873_), .A2(new_n874_), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n882_), .B(new_n883_), .C1(new_n884_), .C2(new_n872_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n880_), .A2(new_n885_), .ZN(G1348gat));
  NAND2_X1  g685(.A1(new_n820_), .A2(new_n868_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n285_), .B1(new_n888_), .B2(new_n554_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n278_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n867_), .ZN(new_n891_));
  AND3_X1   g690(.A1(new_n891_), .A2(G176gat), .A3(new_n554_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n889_), .B1(new_n890_), .B2(new_n892_), .ZN(G1349gat));
  NAND3_X1  g692(.A1(new_n890_), .A2(new_n605_), .A3(new_n891_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n599_), .B1(new_n324_), .B2(new_n326_), .ZN(new_n895_));
  AOI22_X1  g694(.A1(new_n894_), .A2(new_n292_), .B1(new_n888_), .B2(new_n895_), .ZN(G1350gat));
  NAND3_X1  g695(.A1(new_n888_), .A2(new_n327_), .A3(new_n610_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT127), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n888_), .A2(new_n582_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n898_), .B1(new_n899_), .B2(G190gat), .ZN(new_n900_));
  AOI211_X1 g699(.A(KEYINPUT127), .B(new_n293_), .C1(new_n888_), .C2(new_n582_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n897_), .B1(new_n900_), .B2(new_n901_), .ZN(G1351gat));
  NOR4_X1   g701(.A1(new_n699_), .A2(new_n414_), .A3(new_n279_), .A4(new_n432_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n852_), .A2(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(G197gat), .B1(new_n905_), .B2(new_n604_), .ZN(new_n906_));
  NOR3_X1   g705(.A1(new_n904_), .A2(new_n238_), .A3(new_n501_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n906_), .A2(new_n907_), .ZN(G1352gat));
  NAND3_X1  g707(.A1(new_n852_), .A2(new_n554_), .A3(new_n903_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(G204gat), .ZN(G1353gat));
  XNOR2_X1  g709(.A(KEYINPUT63), .B(G211gat), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n904_), .A2(new_n599_), .A3(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n905_), .A2(new_n605_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n912_), .B1(new_n913_), .B2(new_n914_), .ZN(G1354gat));
  OR3_X1    g714(.A1(new_n904_), .A2(G218gat), .A3(new_n609_), .ZN(new_n916_));
  OAI21_X1  g715(.A(G218gat), .B1(new_n904_), .B2(new_n848_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(G1355gat));
endmodule


