//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 1 0 1 1 0 0 0 0 0 1 0 1 1 1 1 1 0 1 0 0 0 0 0 0 0 0 0 1 1 0 0 0 1 1 1 1 0 0 1 1 0 1 1 0 1 0 0 1 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n747_, new_n748_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n788_, new_n789_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n905_, new_n906_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n915_, new_n916_, new_n917_,
    new_n919_, new_n921_, new_n922_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n960_,
    new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n967_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n983_, new_n984_, new_n985_;
  INV_X1    g000(.A(KEYINPUT98), .ZN(new_n202_));
  NOR2_X1   g001(.A1(G141gat), .A2(G148gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT3), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n204_), .A2(KEYINPUT86), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT86), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n206_), .A2(KEYINPUT3), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n203_), .B1(new_n205_), .B2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT87), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT2), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n209_), .A2(KEYINPUT2), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G141gat), .A2(G148gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n210_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n203_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n204_), .A2(KEYINPUT86), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n209_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n208_), .A2(new_n213_), .A3(new_n216_), .A4(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT88), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(G141gat), .ZN(new_n221_));
  INV_X1    g020(.A(G148gat), .ZN(new_n222_));
  AOI22_X1  g021(.A1(new_n221_), .A2(new_n222_), .B1(new_n204_), .B2(KEYINPUT86), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n206_), .A2(KEYINPUT3), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(new_n215_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n223_), .B1(new_n203_), .B2(new_n225_), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n226_), .A2(KEYINPUT88), .A3(new_n213_), .A4(new_n217_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G155gat), .A2(G162gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT85), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT85), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n230_), .A2(G155gat), .A3(G162gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(G155gat), .A2(G162gat), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(KEYINPUT89), .B1(new_n232_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT89), .ZN(new_n236_));
  AOI211_X1 g035(.A(new_n236_), .B(new_n233_), .C1(new_n229_), .C2(new_n231_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n235_), .A2(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n220_), .A2(new_n227_), .A3(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n233_), .B1(new_n232_), .B2(KEYINPUT1), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n240_), .B1(KEYINPUT1), .B2(new_n232_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n241_), .A2(new_n214_), .A3(new_n212_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n239_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(G127gat), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n244_), .A2(G134gat), .ZN(new_n245_));
  INV_X1    g044(.A(G134gat), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n246_), .A2(G127gat), .ZN(new_n247_));
  INV_X1    g046(.A(G113gat), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n248_), .A2(G120gat), .ZN(new_n249_));
  INV_X1    g048(.A(G120gat), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n250_), .A2(G113gat), .ZN(new_n251_));
  OAI22_X1  g050(.A1(new_n245_), .A2(new_n247_), .B1(new_n249_), .B2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G127gat), .B(G134gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G113gat), .B(G120gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  AND3_X1   g054(.A1(new_n252_), .A2(new_n255_), .A3(KEYINPUT84), .ZN(new_n256_));
  AOI21_X1  g055(.A(KEYINPUT84), .B1(new_n252_), .B2(new_n255_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n243_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n252_), .A2(new_n255_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n239_), .A2(new_n261_), .A3(new_n242_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G225gat), .A2(G233gat), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n260_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  AND3_X1   g063(.A1(new_n239_), .A2(new_n261_), .A3(new_n242_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n258_), .B1(new_n239_), .B2(new_n242_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n267_));
  NOR3_X1   g066(.A1(new_n265_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n243_), .A2(new_n267_), .A3(new_n259_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n263_), .B(KEYINPUT94), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n264_), .B1(new_n268_), .B2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G1gat), .B(G29gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(G85gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT0), .B(G57gat), .ZN(new_n275_));
  XOR2_X1   g074(.A(new_n274_), .B(new_n275_), .Z(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n272_), .A2(new_n277_), .ZN(new_n278_));
  OAI211_X1 g077(.A(new_n276_), .B(new_n264_), .C1(new_n268_), .C2(new_n271_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT27), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G8gat), .B(G36gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT18), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G64gat), .B(G92gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G211gat), .B(G218gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G197gat), .A2(G204gat), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(G197gat), .A2(G204gat), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT21), .ZN(new_n292_));
  NOR3_X1   g091(.A1(new_n290_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  OR2_X1    g092(.A1(G197gat), .A2(G204gat), .ZN(new_n294_));
  AOI21_X1  g093(.A(KEYINPUT21), .B1(new_n294_), .B2(new_n289_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n288_), .B1(new_n293_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n288_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n294_), .A2(KEYINPUT21), .A3(new_n289_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n296_), .A2(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(G169gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G183gat), .A2(G190gat), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT23), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n306_));
  OAI211_X1 g105(.A(new_n305_), .B(new_n306_), .C1(G183gat), .C2(G190gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n302_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n305_), .A2(new_n306_), .ZN(new_n309_));
  OR2_X1    g108(.A1(G169gat), .A2(G176gat), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n310_), .A2(KEYINPUT24), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n309_), .A2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT25), .B(G183gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT26), .B(G190gat), .ZN(new_n314_));
  OAI21_X1  g113(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G169gat), .A2(G176gat), .ZN(new_n317_));
  AOI22_X1  g116(.A1(new_n313_), .A2(new_n314_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT82), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n312_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(G183gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT25), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT25), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(G183gat), .ZN(new_n324_));
  INV_X1    g123(.A(G190gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(KEYINPUT26), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT26), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(G190gat), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n322_), .A2(new_n324_), .A3(new_n326_), .A4(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n310_), .A2(KEYINPUT24), .A3(new_n317_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n331_), .A2(KEYINPUT82), .ZN(new_n332_));
  OAI211_X1 g131(.A(new_n300_), .B(new_n308_), .C1(new_n320_), .C2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT20), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT93), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G226gat), .A2(G233gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT19), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT92), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n333_), .A2(KEYINPUT93), .A3(KEYINPUT20), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n318_), .A2(new_n312_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(new_n308_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n292_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n297_), .B1(new_n343_), .B2(new_n298_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n293_), .A2(new_n288_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n342_), .A2(new_n346_), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n336_), .A2(new_n339_), .A3(new_n340_), .A4(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n331_), .A2(KEYINPUT82), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n318_), .A2(new_n319_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n349_), .A2(new_n350_), .A3(new_n312_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n300_), .B1(new_n351_), .B2(new_n308_), .ZN(new_n352_));
  OAI21_X1  g151(.A(KEYINPUT20), .B1(new_n342_), .B2(new_n346_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n338_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n287_), .B1(new_n348_), .B2(new_n354_), .ZN(new_n355_));
  NOR3_X1   g154(.A1(new_n352_), .A2(new_n353_), .A3(new_n338_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  AND3_X1   g156(.A1(new_n333_), .A2(KEYINPUT93), .A3(KEYINPUT20), .ZN(new_n358_));
  AOI21_X1  g157(.A(KEYINPUT93), .B1(new_n333_), .B2(KEYINPUT20), .ZN(new_n359_));
  INV_X1    g158(.A(new_n347_), .ZN(new_n360_));
  NOR3_X1   g159(.A1(new_n358_), .A2(new_n359_), .A3(new_n360_), .ZN(new_n361_));
  OAI211_X1 g160(.A(new_n357_), .B(new_n287_), .C1(new_n361_), .C2(new_n339_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n355_), .B1(new_n362_), .B2(KEYINPUT97), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n336_), .A2(new_n340_), .A3(new_n347_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n339_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT97), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n366_), .A2(new_n367_), .A3(new_n357_), .A4(new_n287_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n282_), .B1(new_n363_), .B2(new_n368_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n359_), .A2(new_n360_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n339_), .B1(new_n370_), .B2(new_n340_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n286_), .B1(new_n371_), .B2(new_n356_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(new_n362_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n373_), .A2(KEYINPUT27), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n281_), .B1(new_n369_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(G78gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n243_), .A2(KEYINPUT29), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n376_), .B1(new_n377_), .B2(new_n346_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT29), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n379_), .B1(new_n239_), .B2(new_n242_), .ZN(new_n380_));
  NOR3_X1   g179(.A1(new_n380_), .A2(G78gat), .A3(new_n300_), .ZN(new_n381_));
  INV_X1    g180(.A(G106gat), .ZN(new_n382_));
  NOR3_X1   g181(.A1(new_n378_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n377_), .A2(new_n376_), .A3(new_n346_), .ZN(new_n384_));
  OAI21_X1  g183(.A(G78gat), .B1(new_n380_), .B2(new_n300_), .ZN(new_n385_));
  AOI21_X1  g184(.A(G106gat), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n239_), .A2(new_n379_), .A3(new_n242_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  NOR3_X1   g188(.A1(new_n383_), .A2(new_n386_), .A3(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n389_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n382_), .B1(new_n378_), .B2(new_n381_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n384_), .A2(G106gat), .A3(new_n385_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n391_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G228gat), .A2(G233gat), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT91), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n395_), .B1(new_n300_), .B2(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G22gat), .B(G50gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NOR3_X1   g199(.A1(new_n390_), .A2(new_n394_), .A3(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n389_), .B1(new_n383_), .B2(new_n386_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n392_), .A2(new_n393_), .A3(new_n391_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n399_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n401_), .A2(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n202_), .B1(new_n375_), .B2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n362_), .A2(KEYINPUT97), .ZN(new_n407_));
  INV_X1    g206(.A(new_n355_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n407_), .A2(new_n368_), .A3(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT27), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n287_), .B1(new_n366_), .B2(new_n357_), .ZN(new_n411_));
  AOI211_X1 g210(.A(new_n356_), .B(new_n286_), .C1(new_n364_), .C2(new_n365_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(new_n282_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n410_), .A2(new_n414_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n400_), .B1(new_n390_), .B2(new_n394_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n402_), .A2(new_n399_), .A3(new_n403_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n415_), .A2(KEYINPUT98), .A3(new_n281_), .A4(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT33), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n279_), .A2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n260_), .A2(KEYINPUT4), .A3(new_n262_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n422_), .A2(new_n269_), .A3(new_n270_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n423_), .A2(KEYINPUT33), .A3(new_n276_), .A4(new_n264_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n265_), .A2(new_n266_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n276_), .B1(new_n425_), .B2(new_n270_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n422_), .A2(new_n263_), .A3(new_n269_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n421_), .A2(new_n424_), .A3(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT95), .B1(new_n429_), .B2(new_n373_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT95), .ZN(new_n431_));
  AOI22_X1  g230(.A1(new_n279_), .A2(new_n420_), .B1(new_n427_), .B2(new_n426_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n413_), .A2(new_n431_), .A3(new_n432_), .A4(new_n424_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n348_), .A2(new_n354_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n287_), .A2(KEYINPUT32), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(KEYINPUT96), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT96), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n434_), .A2(new_n439_), .A3(new_n436_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n366_), .A2(new_n357_), .A3(new_n435_), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n280_), .A2(new_n438_), .A3(new_n440_), .A4(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n430_), .A2(new_n433_), .A3(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(new_n405_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n406_), .A2(new_n419_), .A3(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n351_), .A2(new_n308_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G15gat), .B(G43gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(KEYINPUT83), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(KEYINPUT30), .ZN(new_n449_));
  XOR2_X1   g248(.A(new_n446_), .B(new_n449_), .Z(new_n450_));
  NAND2_X1  g249(.A1(G227gat), .A2(G233gat), .ZN(new_n451_));
  INV_X1    g250(.A(G71gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n451_), .B(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n450_), .B(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n258_), .B(KEYINPUT31), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(G99gat), .ZN(new_n456_));
  OR2_X1    g255(.A1(new_n454_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n454_), .A2(new_n456_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n445_), .A2(new_n459_), .ZN(new_n460_));
  NOR3_X1   g259(.A1(new_n375_), .A2(new_n459_), .A3(new_n418_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(KEYINPUT66), .B(G71gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(G78gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G57gat), .B(G64gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT11), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n466_), .A2(KEYINPUT11), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n465_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n464_), .B(new_n376_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(new_n467_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT76), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G127gat), .B(G155gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT16), .ZN(new_n476_));
  XOR2_X1   g275(.A(G183gat), .B(G211gat), .Z(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT17), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n474_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G15gat), .B(G22gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT74), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT14), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n483_), .B1(G1gat), .B2(G8gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(KEYINPUT75), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n482_), .A2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G1gat), .B(G8gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n487_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n482_), .A2(new_n489_), .A3(new_n485_), .ZN(new_n490_));
  AND2_X1   g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n480_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n488_), .A2(new_n490_), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n493_), .B(new_n474_), .C1(new_n479_), .C2(new_n478_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G231gat), .A2(G233gat), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  AND3_X1   g295(.A1(new_n492_), .A2(new_n494_), .A3(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n496_), .B1(new_n492_), .B2(new_n494_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n473_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n492_), .A2(new_n494_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(new_n495_), .ZN(new_n501_));
  AND2_X1   g300(.A1(new_n470_), .A2(new_n472_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n492_), .A2(new_n496_), .A3(new_n494_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n501_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n478_), .A2(new_n479_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n499_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(KEYINPUT77), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT77), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n499_), .A2(new_n504_), .A3(new_n508_), .A4(new_n505_), .ZN(new_n509_));
  AND3_X1   g308(.A1(new_n507_), .A2(KEYINPUT78), .A3(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(KEYINPUT78), .B1(new_n507_), .B2(new_n509_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  XOR2_X1   g312(.A(G29gat), .B(G36gat), .Z(new_n514_));
  XOR2_X1   g313(.A(G43gat), .B(G50gat), .Z(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT15), .ZN(new_n517_));
  XOR2_X1   g316(.A(KEYINPUT10), .B(G99gat), .Z(new_n518_));
  XOR2_X1   g317(.A(KEYINPUT64), .B(G106gat), .Z(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  XOR2_X1   g319(.A(G85gat), .B(G92gat), .Z(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(KEYINPUT9), .ZN(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT65), .B(G85gat), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT9), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n523_), .A2(new_n524_), .A3(G92gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G99gat), .A2(G106gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT6), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n520_), .A2(new_n522_), .A3(new_n525_), .A4(new_n527_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(G99gat), .A2(G106gat), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT7), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT6), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n526_), .B(new_n532_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n521_), .B1(new_n531_), .B2(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n534_), .A2(KEYINPUT8), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G85gat), .B(G92gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n529_), .B(KEYINPUT7), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n536_), .B1(new_n537_), .B2(new_n527_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT8), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n528_), .B1(new_n535_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n517_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n528_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n534_), .A2(KEYINPUT8), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n538_), .A2(new_n539_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n543_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(new_n516_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G232gat), .A2(G233gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT35), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n542_), .A2(new_n547_), .A3(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n550_), .A2(new_n551_), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n554_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n555_), .A2(KEYINPUT73), .A3(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G190gat), .B(G218gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT71), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT72), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G134gat), .B(G162gat), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n560_), .B(new_n561_), .Z(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n557_), .A2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n555_), .A2(new_n556_), .A3(new_n562_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT36), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n564_), .A2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n557_), .A2(new_n566_), .A3(new_n563_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(KEYINPUT37), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT37), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n568_), .A2(new_n572_), .A3(new_n569_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n571_), .A2(new_n573_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n513_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT68), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n576_), .B1(new_n546_), .B2(new_n502_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(KEYINPUT12), .ZN(new_n578_));
  AOI21_X1  g377(.A(KEYINPUT68), .B1(new_n541_), .B2(new_n473_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT12), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G230gat), .A2(G233gat), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n546_), .A2(new_n502_), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n578_), .A2(new_n581_), .A3(new_n582_), .A4(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n582_), .ZN(new_n585_));
  OAI21_X1  g384(.A(KEYINPUT67), .B1(new_n546_), .B2(new_n502_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(new_n583_), .ZN(new_n587_));
  NOR3_X1   g386(.A1(new_n546_), .A2(new_n502_), .A3(KEYINPUT67), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n585_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n584_), .A2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G120gat), .B(G148gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT5), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G176gat), .B(G204gat), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n592_), .B(new_n593_), .Z(new_n594_));
  NAND2_X1  g393(.A1(new_n590_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n594_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n584_), .A2(new_n589_), .A3(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n598_), .B1(KEYINPUT69), .B2(KEYINPUT13), .ZN(new_n599_));
  AND2_X1   g398(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n600_));
  NOR2_X1   g399(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n601_));
  OAI211_X1 g400(.A(new_n595_), .B(new_n597_), .C1(new_n600_), .C2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n599_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G113gat), .B(G141gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G169gat), .B(G197gat), .ZN(new_n606_));
  XOR2_X1   g405(.A(new_n605_), .B(new_n606_), .Z(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(KEYINPUT80), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n491_), .A2(KEYINPUT79), .A3(new_n516_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT79), .ZN(new_n612_));
  INV_X1    g411(.A(new_n516_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n612_), .B1(new_n493_), .B2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n611_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(G229gat), .A2(G233gat), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n517_), .A2(new_n493_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n615_), .A2(new_n616_), .A3(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n516_), .B1(new_n488_), .B2(new_n490_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n620_), .B1(new_n611_), .B2(new_n614_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n621_), .A2(new_n616_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n610_), .B1(new_n619_), .B2(new_n622_), .ZN(new_n623_));
  OAI211_X1 g422(.A(new_n618_), .B(new_n609_), .C1(new_n616_), .C2(new_n621_), .ZN(new_n624_));
  AND3_X1   g423(.A1(new_n623_), .A2(KEYINPUT81), .A3(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(KEYINPUT81), .B1(new_n623_), .B2(new_n624_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n604_), .A2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n463_), .A2(new_n575_), .A3(new_n628_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n629_), .A2(G1gat), .A3(new_n281_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT99), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n631_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT38), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n623_), .A2(new_n624_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n603_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n507_), .A2(new_n509_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT100), .ZN(new_n642_));
  INV_X1    g441(.A(new_n570_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n463_), .A2(new_n642_), .A3(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n461_), .B1(new_n445_), .B2(new_n459_), .ZN(new_n645_));
  OAI21_X1  g444(.A(KEYINPUT100), .B1(new_n645_), .B2(new_n570_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n641_), .B1(new_n644_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  OAI21_X1  g447(.A(G1gat), .B1(new_n648_), .B2(new_n281_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n632_), .A2(KEYINPUT38), .A3(new_n633_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n636_), .A2(new_n649_), .A3(new_n650_), .ZN(G1324gat));
  INV_X1    g450(.A(G8gat), .ZN(new_n652_));
  INV_X1    g451(.A(new_n415_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n652_), .B1(new_n647_), .B2(new_n653_), .ZN(new_n654_));
  OR2_X1    g453(.A1(new_n654_), .A2(KEYINPUT39), .ZN(new_n655_));
  INV_X1    g454(.A(new_n629_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n415_), .A2(G8gat), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n656_), .A2(KEYINPUT101), .A3(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT101), .ZN(new_n659_));
  INV_X1    g458(.A(new_n657_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n659_), .B1(new_n629_), .B2(new_n660_), .ZN(new_n661_));
  AOI22_X1  g460(.A1(new_n654_), .A2(KEYINPUT39), .B1(new_n658_), .B2(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n655_), .A2(new_n662_), .A3(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n663_), .B1(new_n655_), .B2(new_n662_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1325gat));
  OR3_X1    g465(.A1(new_n629_), .A2(G15gat), .A3(new_n459_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n459_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n647_), .A2(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(KEYINPUT103), .B(KEYINPUT41), .ZN(new_n670_));
  AND3_X1   g469(.A1(new_n669_), .A2(G15gat), .A3(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n670_), .B1(new_n669_), .B2(G15gat), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n667_), .B1(new_n671_), .B2(new_n672_), .ZN(G1326gat));
  INV_X1    g472(.A(G22gat), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n656_), .A2(new_n674_), .A3(new_n418_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT42), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n647_), .A2(new_n418_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n676_), .B1(new_n677_), .B2(G22gat), .ZN(new_n678_));
  AOI211_X1 g477(.A(KEYINPUT42), .B(new_n674_), .C1(new_n647_), .C2(new_n418_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n675_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(KEYINPUT104), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT104), .ZN(new_n682_));
  OAI211_X1 g481(.A(new_n682_), .B(new_n675_), .C1(new_n678_), .C2(new_n679_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n681_), .A2(new_n683_), .ZN(G1327gat));
  NOR2_X1   g483(.A1(new_n512_), .A2(new_n643_), .ZN(new_n685_));
  AND3_X1   g484(.A1(new_n463_), .A2(new_n628_), .A3(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(G29gat), .B1(new_n686_), .B2(new_n280_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n638_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n513_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT43), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n691_), .B1(new_n463_), .B2(new_n574_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n573_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n572_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  NOR3_X1   g494(.A1(new_n645_), .A2(KEYINPUT43), .A3(new_n695_), .ZN(new_n696_));
  OAI211_X1 g495(.A(KEYINPUT44), .B(new_n690_), .C1(new_n692_), .C2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(KEYINPUT105), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n415_), .A2(new_n281_), .A3(new_n418_), .ZN(new_n699_));
  AOI22_X1  g498(.A1(new_n699_), .A2(new_n202_), .B1(new_n405_), .B2(new_n443_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n668_), .B1(new_n700_), .B2(new_n419_), .ZN(new_n701_));
  OAI211_X1 g500(.A(new_n691_), .B(new_n574_), .C1(new_n701_), .C2(new_n461_), .ZN(new_n702_));
  OAI21_X1  g501(.A(KEYINPUT43), .B1(new_n645_), .B2(new_n695_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n689_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT105), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n704_), .A2(new_n705_), .A3(KEYINPUT44), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n698_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n704_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n707_), .A2(new_n710_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n280_), .A2(G29gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n687_), .B1(new_n711_), .B2(new_n712_), .ZN(G1328gat));
  INV_X1    g512(.A(KEYINPUT46), .ZN(new_n714_));
  INV_X1    g513(.A(G36gat), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n653_), .B1(new_n704_), .B2(KEYINPUT44), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n715_), .B1(new_n707_), .B2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT45), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT106), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n415_), .A2(G36gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n686_), .B2(new_n721_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n463_), .A2(new_n628_), .A3(new_n685_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n721_), .ZN(new_n724_));
  NOR3_X1   g523(.A1(new_n723_), .A2(KEYINPUT106), .A3(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n719_), .B1(new_n722_), .B2(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n686_), .A2(new_n720_), .A3(new_n721_), .ZN(new_n727_));
  OAI21_X1  g526(.A(KEYINPUT106), .B1(new_n723_), .B2(new_n724_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n727_), .A2(KEYINPUT45), .A3(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n726_), .A2(new_n729_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n714_), .B1(new_n718_), .B2(new_n730_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n726_), .A2(new_n729_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n716_), .B1(new_n698_), .B2(new_n706_), .ZN(new_n733_));
  OAI211_X1 g532(.A(new_n732_), .B(KEYINPUT46), .C1(new_n733_), .C2(new_n715_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n731_), .A2(new_n734_), .ZN(G1329gat));
  INV_X1    g534(.A(G43gat), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n459_), .A2(new_n736_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n697_), .A2(KEYINPUT105), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n705_), .B1(new_n704_), .B2(KEYINPUT44), .ZN(new_n739_));
  OAI211_X1 g538(.A(new_n710_), .B(new_n737_), .C1(new_n738_), .C2(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n736_), .B1(new_n723_), .B2(new_n459_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT47), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT47), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n740_), .A2(new_n744_), .A3(new_n741_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1330gat));
  AOI21_X1  g545(.A(G50gat), .B1(new_n686_), .B2(new_n418_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n418_), .A2(G50gat), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n711_), .B2(new_n748_), .ZN(G1331gat));
  NOR3_X1   g548(.A1(new_n645_), .A2(new_n603_), .A3(new_n637_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n750_), .A2(new_n575_), .ZN(new_n751_));
  INV_X1    g550(.A(G57gat), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n751_), .A2(new_n752_), .A3(new_n280_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT78), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n639_), .A2(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n507_), .A2(KEYINPUT78), .A3(new_n509_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n755_), .A2(new_n756_), .A3(new_n627_), .ZN(new_n757_));
  AOI211_X1 g556(.A(new_n603_), .B(new_n757_), .C1(new_n644_), .C2(new_n646_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n758_), .A2(new_n280_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n753_), .B1(new_n759_), .B2(new_n752_), .ZN(G1332gat));
  NOR2_X1   g559(.A1(new_n415_), .A2(G64gat), .ZN(new_n761_));
  XOR2_X1   g560(.A(new_n761_), .B(KEYINPUT107), .Z(new_n762_));
  NAND2_X1  g561(.A1(new_n751_), .A2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n758_), .A2(new_n653_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT48), .ZN(new_n765_));
  AND3_X1   g564(.A1(new_n764_), .A2(new_n765_), .A3(G64gat), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n765_), .B1(new_n764_), .B2(G64gat), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n763_), .B1(new_n766_), .B2(new_n767_), .ZN(G1333gat));
  NAND3_X1  g567(.A1(new_n751_), .A2(new_n452_), .A3(new_n668_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT49), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n758_), .A2(new_n668_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n771_), .B2(G71gat), .ZN(new_n772_));
  AOI211_X1 g571(.A(KEYINPUT49), .B(new_n452_), .C1(new_n758_), .C2(new_n668_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n769_), .B1(new_n772_), .B2(new_n773_), .ZN(G1334gat));
  NAND3_X1  g573(.A1(new_n751_), .A2(new_n376_), .A3(new_n418_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT50), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n758_), .A2(new_n418_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n776_), .B1(new_n777_), .B2(G78gat), .ZN(new_n778_));
  AOI211_X1 g577(.A(KEYINPUT50), .B(new_n376_), .C1(new_n758_), .C2(new_n418_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n775_), .B1(new_n778_), .B2(new_n779_), .ZN(G1335gat));
  NOR2_X1   g579(.A1(new_n603_), .A2(new_n637_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n513_), .A2(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n782_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n280_), .A2(new_n523_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n750_), .A2(new_n280_), .A3(new_n685_), .ZN(new_n785_));
  INV_X1    g584(.A(G85gat), .ZN(new_n786_));
  AOI22_X1  g585(.A1(new_n783_), .A2(new_n784_), .B1(new_n785_), .B2(new_n786_), .ZN(G1336gat));
  NAND3_X1  g586(.A1(new_n750_), .A2(new_n653_), .A3(new_n685_), .ZN(new_n788_));
  INV_X1    g587(.A(G92gat), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n790_), .A2(KEYINPUT108), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n790_), .A2(KEYINPUT108), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n415_), .A2(new_n789_), .ZN(new_n793_));
  AOI211_X1 g592(.A(new_n791_), .B(new_n792_), .C1(new_n783_), .C2(new_n793_), .ZN(G1337gat));
  NAND4_X1  g593(.A1(new_n750_), .A2(new_n518_), .A3(new_n668_), .A4(new_n685_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n783_), .A2(new_n668_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n796_), .B1(new_n797_), .B2(G99gat), .ZN(new_n798_));
  NAND2_X1  g597(.A1(KEYINPUT109), .A2(KEYINPUT51), .ZN(new_n799_));
  MUX2_X1   g598(.A(KEYINPUT51), .B(new_n799_), .S(KEYINPUT110), .Z(new_n800_));
  NAND2_X1  g599(.A1(new_n798_), .A2(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n801_), .B1(new_n798_), .B2(new_n799_), .ZN(G1338gat));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n803_));
  OAI21_X1  g602(.A(G106gat), .B1(new_n803_), .B2(KEYINPUT112), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(new_n783_), .B2(new_n418_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(KEYINPUT112), .ZN(new_n806_));
  OR2_X1    g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n805_), .A2(new_n806_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n750_), .A2(new_n519_), .A3(new_n418_), .A4(new_n685_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT111), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n809_), .B(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n807_), .A2(new_n808_), .A3(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(KEYINPUT53), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT53), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n807_), .A2(new_n814_), .A3(new_n808_), .A4(new_n811_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n813_), .A2(new_n815_), .ZN(G1339gat));
  OAI21_X1  g615(.A(new_n583_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n577_), .A2(KEYINPUT12), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n585_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT114), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT114), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n821_), .B(new_n585_), .C1(new_n817_), .C2(new_n818_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n584_), .A2(new_n823_), .ZN(new_n824_));
  AOI22_X1  g623(.A1(new_n577_), .A2(KEYINPUT12), .B1(new_n546_), .B2(new_n502_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n825_), .A2(KEYINPUT55), .A3(new_n582_), .A4(new_n581_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n820_), .A2(new_n822_), .A3(new_n824_), .A4(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n594_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT56), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n827_), .A2(KEYINPUT56), .A3(new_n594_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n616_), .B1(new_n615_), .B2(new_n617_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n616_), .ZN(new_n833_));
  AOI211_X1 g632(.A(new_n833_), .B(new_n620_), .C1(new_n611_), .C2(new_n614_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n608_), .B1(new_n832_), .B2(new_n834_), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n618_), .B(new_n607_), .C1(new_n616_), .C2(new_n621_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n835_), .A2(new_n836_), .A3(new_n597_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT115), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n835_), .A2(new_n836_), .A3(new_n597_), .A4(KEYINPUT115), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n830_), .A2(new_n831_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(KEYINPUT116), .B(KEYINPUT58), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  OAI211_X1 g642(.A(KEYINPUT117), .B(new_n574_), .C1(new_n841_), .C2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n841_), .A2(KEYINPUT58), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n839_), .A2(new_n840_), .ZN(new_n847_));
  AND3_X1   g646(.A1(new_n827_), .A2(KEYINPUT56), .A3(new_n594_), .ZN(new_n848_));
  AOI21_X1  g647(.A(KEYINPUT56), .B1(new_n827_), .B2(new_n594_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n847_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n842_), .ZN(new_n851_));
  AOI21_X1  g650(.A(KEYINPUT117), .B1(new_n851_), .B2(new_n574_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n846_), .A2(new_n852_), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n637_), .A2(new_n597_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n854_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n598_), .A2(new_n835_), .A3(new_n836_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n570_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(KEYINPUT57), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n639_), .B1(new_n853_), .B2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT113), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n755_), .A2(new_n860_), .A3(new_n627_), .A4(new_n756_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n861_), .A2(new_n695_), .A3(new_n603_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n860_), .B1(new_n512_), .B2(new_n627_), .ZN(new_n863_));
  OAI21_X1  g662(.A(KEYINPUT54), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n757_), .A2(KEYINPUT113), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n574_), .A2(new_n604_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n865_), .A2(new_n866_), .A3(new_n867_), .A4(new_n861_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n864_), .A2(new_n868_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n859_), .A2(KEYINPUT118), .A3(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT118), .ZN(new_n871_));
  INV_X1    g670(.A(new_n639_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT117), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n830_), .A2(new_n831_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n843_), .B1(new_n874_), .B2(new_n847_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n873_), .B1(new_n875_), .B2(new_n695_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n876_), .A2(new_n844_), .A3(new_n845_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n855_), .A2(new_n856_), .ZN(new_n878_));
  AOI21_X1  g677(.A(KEYINPUT57), .B1(new_n878_), .B2(new_n643_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n880_));
  AOI211_X1 g679(.A(new_n880_), .B(new_n570_), .C1(new_n855_), .C2(new_n856_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n879_), .A2(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n872_), .B1(new_n877_), .B2(new_n882_), .ZN(new_n883_));
  AND2_X1   g682(.A1(new_n864_), .A2(new_n868_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n871_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n653_), .A2(new_n281_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n418_), .A2(new_n459_), .ZN(new_n887_));
  AND2_X1   g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n870_), .A2(new_n885_), .A3(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(KEYINPUT59), .ZN(new_n890_));
  INV_X1    g689(.A(new_n627_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n512_), .B1(new_n877_), .B2(new_n882_), .ZN(new_n892_));
  OR2_X1    g691(.A1(new_n892_), .A2(new_n884_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n894_));
  AND2_X1   g693(.A1(new_n888_), .A2(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n893_), .A2(new_n895_), .ZN(new_n896_));
  AND3_X1   g695(.A1(new_n890_), .A2(new_n891_), .A3(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n637_), .A2(new_n248_), .ZN(new_n898_));
  OAI22_X1  g697(.A1(new_n897_), .A2(new_n248_), .B1(new_n889_), .B2(new_n898_), .ZN(G1340gat));
  AND3_X1   g698(.A1(new_n890_), .A2(new_n604_), .A3(new_n896_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n250_), .B1(new_n603_), .B2(KEYINPUT60), .ZN(new_n901_));
  OR2_X1    g700(.A1(new_n250_), .A2(KEYINPUT60), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  OAI22_X1  g702(.A1(new_n900_), .A2(new_n250_), .B1(new_n889_), .B2(new_n903_), .ZN(G1341gat));
  AND3_X1   g703(.A1(new_n890_), .A2(new_n872_), .A3(new_n896_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n512_), .A2(new_n244_), .ZN(new_n906_));
  OAI22_X1  g705(.A1(new_n905_), .A2(new_n244_), .B1(new_n889_), .B2(new_n906_), .ZN(G1342gat));
  NAND4_X1  g706(.A1(new_n890_), .A2(G134gat), .A3(new_n574_), .A4(new_n896_), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n870_), .A2(new_n885_), .A3(new_n570_), .A4(new_n888_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT119), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n909_), .A2(new_n910_), .A3(new_n246_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n909_), .A2(new_n246_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(KEYINPUT119), .ZN(new_n913_));
  AND3_X1   g712(.A1(new_n908_), .A2(new_n911_), .A3(new_n913_), .ZN(G1343gat));
  NOR2_X1   g713(.A1(new_n668_), .A2(new_n405_), .ZN(new_n915_));
  AND3_X1   g714(.A1(new_n870_), .A2(new_n885_), .A3(new_n915_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n916_), .A2(new_n637_), .A3(new_n886_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g717(.A1(new_n916_), .A2(new_n604_), .A3(new_n886_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g719(.A1(new_n916_), .A2(new_n512_), .A3(new_n886_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(KEYINPUT61), .B(G155gat), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n921_), .B(new_n922_), .ZN(G1346gat));
  NAND3_X1  g722(.A1(new_n916_), .A2(new_n574_), .A3(new_n886_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(G162gat), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n643_), .A2(G162gat), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n916_), .A2(new_n886_), .A3(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n925_), .A2(new_n927_), .ZN(G1347gat));
  NOR2_X1   g727(.A1(new_n415_), .A2(new_n280_), .ZN(new_n929_));
  AND2_X1   g728(.A1(new_n929_), .A2(new_n887_), .ZN(new_n930_));
  OAI211_X1 g729(.A(new_n637_), .B(new_n930_), .C1(new_n892_), .C2(new_n884_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n931_), .A2(G169gat), .ZN(new_n932_));
  OR2_X1    g731(.A1(new_n932_), .A2(KEYINPUT120), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(KEYINPUT120), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n933_), .A2(KEYINPUT62), .A3(new_n934_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT62), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n932_), .A2(KEYINPUT120), .A3(new_n936_), .ZN(new_n937_));
  XOR2_X1   g736(.A(KEYINPUT22), .B(G169gat), .Z(new_n938_));
  OR2_X1    g737(.A1(new_n931_), .A2(new_n938_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n935_), .A2(new_n937_), .A3(new_n939_), .ZN(G1348gat));
  INV_X1    g739(.A(G176gat), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n893_), .A2(new_n930_), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n941_), .B1(new_n942_), .B2(new_n603_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n929_), .A2(new_n668_), .ZN(new_n944_));
  NOR3_X1   g743(.A1(new_n944_), .A2(new_n941_), .A3(new_n603_), .ZN(new_n945_));
  NAND4_X1  g744(.A1(new_n870_), .A2(new_n885_), .A3(new_n405_), .A4(new_n945_), .ZN(new_n946_));
  AND2_X1   g745(.A1(new_n943_), .A2(new_n946_), .ZN(G1349gat));
  NOR2_X1   g746(.A1(new_n513_), .A2(new_n944_), .ZN(new_n948_));
  NAND4_X1  g747(.A1(new_n870_), .A2(new_n885_), .A3(new_n405_), .A4(new_n948_), .ZN(new_n949_));
  AND2_X1   g748(.A1(new_n949_), .A2(new_n321_), .ZN(new_n950_));
  NOR2_X1   g749(.A1(new_n639_), .A2(new_n313_), .ZN(new_n951_));
  OAI211_X1 g750(.A(new_n930_), .B(new_n951_), .C1(new_n892_), .C2(new_n884_), .ZN(new_n952_));
  XNOR2_X1  g751(.A(new_n952_), .B(KEYINPUT121), .ZN(new_n953_));
  OAI21_X1  g752(.A(KEYINPUT122), .B1(new_n950_), .B2(new_n953_), .ZN(new_n954_));
  XOR2_X1   g753(.A(new_n952_), .B(KEYINPUT121), .Z(new_n955_));
  NAND2_X1  g754(.A1(new_n949_), .A2(new_n321_), .ZN(new_n956_));
  INV_X1    g755(.A(KEYINPUT122), .ZN(new_n957_));
  NAND3_X1  g756(.A1(new_n955_), .A2(new_n956_), .A3(new_n957_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n954_), .A2(new_n958_), .ZN(G1350gat));
  OAI21_X1  g758(.A(G190gat), .B1(new_n942_), .B2(new_n695_), .ZN(new_n960_));
  NAND4_X1  g759(.A1(new_n893_), .A2(new_n570_), .A3(new_n314_), .A4(new_n930_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n960_), .A2(new_n961_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n962_), .A2(KEYINPUT123), .ZN(new_n963_));
  INV_X1    g762(.A(KEYINPUT123), .ZN(new_n964_));
  NAND3_X1  g763(.A1(new_n960_), .A2(new_n964_), .A3(new_n961_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n963_), .A2(new_n965_), .ZN(G1351gat));
  NAND3_X1  g765(.A1(new_n916_), .A2(new_n637_), .A3(new_n929_), .ZN(new_n967_));
  XNOR2_X1  g766(.A(new_n967_), .B(G197gat), .ZN(G1352gat));
  NAND4_X1  g767(.A1(new_n870_), .A2(new_n885_), .A3(new_n915_), .A4(new_n929_), .ZN(new_n969_));
  NOR2_X1   g768(.A1(new_n969_), .A2(new_n603_), .ZN(new_n970_));
  AND2_X1   g769(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n971_));
  NOR2_X1   g770(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n972_));
  OAI21_X1  g771(.A(new_n970_), .B1(new_n971_), .B2(new_n972_), .ZN(new_n973_));
  OAI21_X1  g772(.A(new_n973_), .B1(new_n970_), .B2(new_n972_), .ZN(G1353gat));
  NOR2_X1   g773(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n975_));
  AND2_X1   g774(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n976_));
  NOR4_X1   g775(.A1(new_n969_), .A2(new_n639_), .A3(new_n975_), .A4(new_n976_), .ZN(new_n977_));
  OAI21_X1  g776(.A(new_n975_), .B1(new_n969_), .B2(new_n639_), .ZN(new_n978_));
  NAND2_X1  g777(.A1(new_n978_), .A2(KEYINPUT125), .ZN(new_n979_));
  INV_X1    g778(.A(KEYINPUT125), .ZN(new_n980_));
  OAI211_X1 g779(.A(new_n980_), .B(new_n975_), .C1(new_n969_), .C2(new_n639_), .ZN(new_n981_));
  AOI21_X1  g780(.A(new_n977_), .B1(new_n979_), .B2(new_n981_), .ZN(G1354gat));
  XOR2_X1   g781(.A(KEYINPUT126), .B(G218gat), .Z(new_n983_));
  NOR3_X1   g782(.A1(new_n969_), .A2(new_n695_), .A3(new_n983_), .ZN(new_n984_));
  NAND3_X1  g783(.A1(new_n916_), .A2(new_n570_), .A3(new_n929_), .ZN(new_n985_));
  AOI21_X1  g784(.A(new_n984_), .B1(new_n985_), .B2(new_n983_), .ZN(G1355gat));
endmodule


