//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 1 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 0 1 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 0 1 0 0 1 0 1 0 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n767_, new_n768_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n896_, new_n897_, new_n899_, new_n900_, new_n901_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n929_, new_n930_,
    new_n931_, new_n933_, new_n934_, new_n935_, new_n936_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n950_, new_n951_;
  INV_X1    g000(.A(KEYINPUT75), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G230gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G71gat), .B(G78gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(G57gat), .B(G64gat), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  AOI21_X1  g005(.A(new_n204_), .B1(new_n206_), .B2(KEYINPUT11), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n207_), .B1(KEYINPUT11), .B2(new_n206_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n206_), .A2(new_n204_), .A3(KEYINPUT11), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT66), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT7), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n211_), .B(new_n212_), .C1(G99gat), .C2(G106gat), .ZN(new_n213_));
  INV_X1    g012(.A(G99gat), .ZN(new_n214_));
  INV_X1    g013(.A(G106gat), .ZN(new_n215_));
  OAI211_X1 g014(.A(new_n214_), .B(new_n215_), .C1(KEYINPUT66), .C2(KEYINPUT7), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n213_), .A2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(KEYINPUT70), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G99gat), .A2(G106gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT6), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT6), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(G99gat), .A3(G106gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n223_), .B(KEYINPUT69), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n218_), .A2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G85gat), .B(G92gat), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT8), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT68), .B(KEYINPUT8), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n217_), .A2(new_n223_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT67), .ZN(new_n232_));
  AOI211_X1 g031(.A(new_n226_), .B(new_n230_), .C1(new_n231_), .C2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n217_), .A2(KEYINPUT67), .A3(new_n223_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n229_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT9), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n237_), .A2(G85gat), .A3(G92gat), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n238_), .B1(new_n226_), .B2(new_n237_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT64), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  XOR2_X1   g040(.A(KEYINPUT10), .B(G99gat), .Z(new_n242_));
  AOI22_X1  g041(.A1(new_n242_), .A2(new_n215_), .B1(new_n220_), .B2(new_n222_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT65), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT65), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n241_), .A2(new_n246_), .A3(new_n243_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n210_), .B1(new_n236_), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n236_), .A2(new_n210_), .A3(new_n248_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n203_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n203_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT72), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT72), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n251_), .A2(new_n255_), .A3(new_n203_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n254_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n210_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT71), .B(KEYINPUT12), .ZN(new_n259_));
  AND2_X1   g058(.A1(new_n245_), .A2(new_n247_), .ZN(new_n260_));
  AOI22_X1  g059(.A1(new_n228_), .A2(KEYINPUT8), .B1(new_n234_), .B2(new_n233_), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n258_), .B(new_n259_), .C1(new_n260_), .C2(new_n261_), .ZN(new_n262_));
  AND2_X1   g061(.A1(KEYINPUT71), .A2(KEYINPUT12), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n262_), .B1(new_n249_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n252_), .B1(new_n257_), .B2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G120gat), .B(G148gat), .ZN(new_n267_));
  INV_X1    g066(.A(G204gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(KEYINPUT5), .B(G176gat), .ZN(new_n270_));
  XOR2_X1   g069(.A(new_n269_), .B(new_n270_), .Z(new_n271_));
  OAI21_X1  g070(.A(KEYINPUT73), .B1(new_n266_), .B2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT73), .ZN(new_n273_));
  INV_X1    g072(.A(new_n271_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n264_), .B1(new_n254_), .B2(new_n256_), .ZN(new_n275_));
  OAI211_X1 g074(.A(new_n273_), .B(new_n274_), .C1(new_n275_), .C2(new_n252_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n272_), .A2(new_n276_), .ZN(new_n277_));
  OR2_X1    g076(.A1(new_n249_), .A2(new_n263_), .ZN(new_n278_));
  AND3_X1   g077(.A1(new_n251_), .A2(new_n255_), .A3(new_n203_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n255_), .B1(new_n251_), .B2(new_n203_), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n278_), .B(new_n262_), .C1(new_n279_), .C2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n252_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n281_), .A2(new_n282_), .A3(new_n271_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT74), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT74), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n266_), .A2(new_n285_), .A3(new_n271_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT13), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n277_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n288_), .B1(new_n277_), .B2(new_n287_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n202_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n277_), .A2(new_n287_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(KEYINPUT13), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n294_), .A2(KEYINPUT75), .A3(new_n289_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n292_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G8gat), .B(G36gat), .ZN(new_n297_));
  INV_X1    g096(.A(G92gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT18), .B(G64gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G226gat), .A2(G233gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT19), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT22), .B(G169gat), .ZN(new_n306_));
  INV_X1    g105(.A(G176gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G183gat), .A2(G190gat), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT23), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n312_));
  OAI211_X1 g111(.A(new_n311_), .B(new_n312_), .C1(G183gat), .C2(G190gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G169gat), .A2(G176gat), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n308_), .A2(new_n313_), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT24), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT85), .B1(G169gat), .B2(G176gat), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NOR3_X1   g117(.A1(KEYINPUT85), .A2(G169gat), .A3(G176gat), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n316_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n311_), .A2(new_n312_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT85), .ZN(new_n323_));
  INV_X1    g122(.A(G169gat), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n323_), .A2(new_n324_), .A3(new_n307_), .ZN(new_n325_));
  NAND4_X1  g124(.A1(new_n325_), .A2(KEYINPUT24), .A3(new_n314_), .A4(new_n317_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n320_), .A2(new_n322_), .A3(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT83), .ZN(new_n328_));
  INV_X1    g127(.A(G183gat), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n328_), .B1(new_n329_), .B2(KEYINPUT25), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT25), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n331_), .A2(KEYINPUT83), .A3(G183gat), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT84), .ZN(new_n333_));
  INV_X1    g132(.A(G190gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(KEYINPUT26), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n330_), .B(new_n332_), .C1(new_n333_), .C2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n329_), .A2(KEYINPUT25), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT26), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(G190gat), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n338_), .A2(G190gat), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n337_), .B(new_n339_), .C1(new_n340_), .C2(KEYINPUT84), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n336_), .A2(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n315_), .B1(new_n327_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT92), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n344_), .A2(new_n268_), .A3(G197gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n268_), .A2(G197gat), .ZN(new_n346_));
  INV_X1    g145(.A(G197gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(G204gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(new_n348_), .ZN(new_n349_));
  OAI211_X1 g148(.A(KEYINPUT21), .B(new_n345_), .C1(new_n349_), .C2(new_n344_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G197gat), .B(G204gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT93), .B(KEYINPUT21), .ZN(new_n352_));
  OR2_X1    g151(.A1(G211gat), .A2(G218gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G211gat), .A2(G218gat), .ZN(new_n354_));
  AOI22_X1  g153(.A1(new_n351_), .A2(new_n352_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n350_), .A2(new_n355_), .ZN(new_n356_));
  AND3_X1   g155(.A1(new_n353_), .A2(KEYINPUT21), .A3(new_n354_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(new_n349_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(KEYINPUT20), .B1(new_n343_), .B2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT96), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n320_), .A2(new_n322_), .A3(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(KEYINPUT24), .B1(new_n325_), .B2(new_n317_), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT96), .B1(new_n363_), .B2(new_n321_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT25), .B(G183gat), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n365_), .A2(new_n335_), .A3(new_n339_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n314_), .A2(KEYINPUT24), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT95), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n314_), .A2(KEYINPUT95), .A3(KEYINPUT24), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n369_), .A2(new_n325_), .A3(new_n317_), .A4(new_n370_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n362_), .A2(new_n364_), .A3(new_n366_), .A4(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(new_n315_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(new_n359_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n360_), .B1(new_n374_), .B2(KEYINPUT97), .ZN(new_n375_));
  AOI22_X1  g174(.A1(new_n350_), .A2(new_n355_), .B1(new_n349_), .B2(new_n357_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n376_), .B1(new_n372_), .B2(new_n315_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT97), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n305_), .B1(new_n375_), .B2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n372_), .A2(new_n376_), .A3(new_n315_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n343_), .A2(new_n359_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n305_), .A2(KEYINPUT20), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n302_), .B1(new_n380_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT20), .ZN(new_n387_));
  AND3_X1   g186(.A1(new_n320_), .A2(new_n322_), .A3(new_n326_), .ZN(new_n388_));
  OR2_X1    g187(.A1(new_n336_), .A2(new_n341_), .ZN(new_n389_));
  AND2_X1   g188(.A1(new_n308_), .A2(new_n314_), .ZN(new_n390_));
  AOI22_X1  g189(.A1(new_n388_), .A2(new_n389_), .B1(new_n390_), .B2(new_n313_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n387_), .B1(new_n391_), .B2(new_n376_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n392_), .B1(new_n378_), .B2(new_n377_), .ZN(new_n393_));
  AOI211_X1 g192(.A(KEYINPUT97), .B(new_n376_), .C1(new_n372_), .C2(new_n315_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n304_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n385_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n395_), .A2(new_n301_), .A3(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n386_), .A2(KEYINPUT98), .A3(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT27), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n374_), .A2(KEYINPUT97), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n400_), .A2(new_n379_), .A3(new_n392_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n385_), .B1(new_n401_), .B2(new_n304_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT98), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n402_), .A2(new_n403_), .A3(new_n301_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n398_), .A2(new_n399_), .A3(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT101), .B(KEYINPUT20), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n381_), .A2(new_n382_), .A3(new_n406_), .ZN(new_n407_));
  AND2_X1   g206(.A1(new_n407_), .A2(new_n304_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n377_), .A2(new_n378_), .ZN(new_n409_));
  NOR3_X1   g208(.A1(new_n409_), .A2(new_n394_), .A3(new_n360_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n408_), .B1(new_n410_), .B2(new_n305_), .ZN(new_n411_));
  OAI211_X1 g210(.A(new_n397_), .B(KEYINPUT27), .C1(new_n411_), .C2(new_n301_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n405_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(KEYINPUT104), .ZN(new_n414_));
  INV_X1    g213(.A(G155gat), .ZN(new_n415_));
  INV_X1    g214(.A(G162gat), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n415_), .A2(new_n416_), .A3(KEYINPUT89), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT89), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n418_), .B1(G155gat), .B2(G162gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G155gat), .A2(G162gat), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT90), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n420_), .B1(new_n423_), .B2(KEYINPUT1), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n421_), .B(KEYINPUT90), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT1), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n424_), .A2(new_n427_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(G141gat), .A2(G148gat), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT88), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G141gat), .A2(G148gat), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT88), .B1(G141gat), .B2(G148gat), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n431_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n428_), .A2(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n429_), .B(KEYINPUT3), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT2), .ZN(new_n438_));
  OR3_X1    g237(.A1(new_n432_), .A2(new_n438_), .A3(KEYINPUT91), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(KEYINPUT91), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n432_), .B1(new_n438_), .B2(KEYINPUT91), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n437_), .A2(new_n439_), .A3(new_n440_), .A4(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n420_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(new_n423_), .A3(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n436_), .A2(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n376_), .B1(new_n445_), .B2(KEYINPUT29), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G22gat), .B(G50gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(KEYINPUT28), .ZN(new_n448_));
  XOR2_X1   g247(.A(G78gat), .B(G106gat), .Z(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  XOR2_X1   g249(.A(new_n446_), .B(new_n450_), .Z(new_n451_));
  NOR2_X1   g250(.A1(new_n445_), .A2(KEYINPUT29), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G228gat), .A2(G233gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(KEYINPUT94), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n452_), .B(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n451_), .B(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT104), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n405_), .A2(new_n457_), .A3(new_n412_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G71gat), .B(G99gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(G15gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(KEYINPUT30), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(new_n391_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G113gat), .B(G120gat), .ZN(new_n463_));
  OR2_X1    g262(.A1(new_n463_), .A2(KEYINPUT87), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(KEYINPUT87), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G127gat), .B(G134gat), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n464_), .A2(new_n465_), .A3(new_n467_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT31), .ZN(new_n472_));
  XOR2_X1   g271(.A(new_n462_), .B(new_n472_), .Z(new_n473_));
  XNOR2_X1  g272(.A(KEYINPUT86), .B(G43gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G227gat), .A2(G233gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n473_), .B(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n434_), .B1(new_n424_), .B2(new_n427_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n443_), .A2(new_n423_), .ZN(new_n479_));
  AND3_X1   g278(.A1(new_n439_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n479_), .B1(new_n480_), .B2(new_n437_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n471_), .B1(new_n478_), .B2(new_n481_), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n436_), .A2(new_n470_), .A3(new_n469_), .A4(new_n444_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n482_), .A2(new_n483_), .A3(KEYINPUT4), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT4), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n445_), .A2(new_n485_), .A3(new_n471_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n484_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G225gat), .A2(G233gat), .ZN(new_n488_));
  XOR2_X1   g287(.A(new_n488_), .B(KEYINPUT99), .Z(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(G1gat), .B(G29gat), .Z(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(G85gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(KEYINPUT0), .B(G57gat), .ZN(new_n493_));
  XOR2_X1   g292(.A(new_n492_), .B(new_n493_), .Z(new_n494_));
  AOI21_X1  g293(.A(new_n489_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n490_), .A2(new_n494_), .A3(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n494_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n489_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n499_), .B1(new_n484_), .B2(new_n486_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n498_), .B1(new_n500_), .B2(new_n495_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n497_), .A2(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n477_), .A2(new_n502_), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n414_), .A2(new_n456_), .A3(new_n458_), .A4(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT105), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  AND3_X1   g305(.A1(new_n405_), .A2(new_n457_), .A3(new_n412_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n457_), .B1(new_n405_), .B2(new_n412_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n509_), .A2(KEYINPUT105), .A3(new_n456_), .A4(new_n503_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT103), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT102), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n375_), .A2(new_n305_), .A3(new_n379_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n407_), .A2(new_n304_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n301_), .A2(KEYINPUT32), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n512_), .B1(new_n515_), .B2(new_n517_), .ZN(new_n518_));
  AOI211_X1 g317(.A(KEYINPUT102), .B(new_n516_), .C1(new_n513_), .C2(new_n514_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n502_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(KEYINPUT100), .B1(new_n402_), .B2(new_n516_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT100), .ZN(new_n522_));
  NOR4_X1   g321(.A1(new_n380_), .A2(new_n522_), .A3(new_n385_), .A4(new_n517_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n511_), .B1(new_n520_), .B2(new_n524_), .ZN(new_n525_));
  OAI21_X1  g324(.A(KEYINPUT102), .B1(new_n411_), .B2(new_n516_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n515_), .A2(new_n512_), .A3(new_n517_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n395_), .A2(new_n396_), .A3(new_n516_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(new_n522_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n402_), .A2(KEYINPUT100), .A3(new_n516_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n528_), .A2(new_n532_), .A3(KEYINPUT103), .A4(new_n502_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n487_), .A2(new_n489_), .ZN(new_n534_));
  AND3_X1   g333(.A1(new_n482_), .A2(new_n489_), .A3(new_n483_), .ZN(new_n535_));
  NOR3_X1   g334(.A1(new_n534_), .A2(new_n498_), .A3(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n501_), .A2(KEYINPUT33), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT33), .ZN(new_n538_));
  OAI211_X1 g337(.A(new_n538_), .B(new_n498_), .C1(new_n500_), .C2(new_n495_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n536_), .B1(new_n537_), .B2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n398_), .A2(new_n404_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n525_), .A2(new_n533_), .A3(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(new_n456_), .ZN(new_n544_));
  NOR3_X1   g343(.A1(new_n413_), .A2(new_n502_), .A3(new_n456_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(new_n546_), .ZN(new_n547_));
  AOI22_X1  g346(.A1(new_n506_), .A2(new_n510_), .B1(new_n547_), .B2(new_n477_), .ZN(new_n548_));
  INV_X1    g347(.A(G1gat), .ZN(new_n549_));
  INV_X1    g348(.A(G8gat), .ZN(new_n550_));
  OAI21_X1  g349(.A(KEYINPUT14), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(KEYINPUT77), .B(G15gat), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(G22gat), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n551_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  XOR2_X1   g354(.A(G1gat), .B(G8gat), .Z(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n552_), .A2(G22gat), .ZN(new_n558_));
  OR3_X1    g357(.A1(new_n555_), .A2(new_n557_), .A3(new_n558_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n557_), .B1(new_n555_), .B2(new_n558_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G29gat), .B(G36gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G43gat), .B(G50gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(new_n561_), .B(new_n564_), .Z(new_n565_));
  NAND3_X1  g364(.A1(new_n565_), .A2(G229gat), .A3(G233gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n564_), .B(KEYINPUT15), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n561_), .A2(new_n567_), .ZN(new_n568_));
  OR2_X1    g367(.A1(new_n568_), .A2(KEYINPUT81), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G229gat), .A2(G233gat), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n559_), .A2(new_n560_), .A3(new_n564_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n568_), .A2(KEYINPUT81), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n569_), .A2(new_n570_), .A3(new_n571_), .A4(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G113gat), .B(G141gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G169gat), .B(G197gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  AND3_X1   g376(.A1(new_n566_), .A2(new_n573_), .A3(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n577_), .B1(new_n566_), .B2(new_n573_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n580_), .B(KEYINPUT82), .Z(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NOR3_X1   g381(.A1(new_n296_), .A2(new_n548_), .A3(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n561_), .B(new_n210_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G231gat), .A2(G233gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  XOR2_X1   g385(.A(G183gat), .B(G211gat), .Z(new_n587_));
  XNOR2_X1  g386(.A(G127gat), .B(G155gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(KEYINPUT79), .B(KEYINPUT16), .Z(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(KEYINPUT17), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n592_), .A2(KEYINPUT78), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n586_), .A2(new_n593_), .ZN(new_n594_));
  AND3_X1   g393(.A1(new_n591_), .A2(KEYINPUT78), .A3(KEYINPUT17), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n591_), .B(KEYINPUT17), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT80), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n595_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  OAI211_X1 g397(.A(new_n586_), .B(new_n598_), .C1(new_n597_), .C2(new_n596_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n594_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n236_), .A2(new_n248_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(new_n567_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n236_), .A2(new_n564_), .A3(new_n248_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G232gat), .A2(G233gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT34), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT35), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n602_), .A2(new_n603_), .A3(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n606_), .A2(new_n607_), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT36), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G190gat), .B(G218gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G134gat), .B(G162gat), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n613_), .B(new_n614_), .Z(new_n615_));
  NAND2_X1  g414(.A1(new_n609_), .A2(new_n610_), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n611_), .A2(new_n612_), .A3(new_n615_), .A4(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(KEYINPUT37), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n615_), .B(KEYINPUT36), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n620_), .B1(new_n611_), .B2(new_n616_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n618_), .A2(new_n621_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n609_), .A2(new_n610_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n609_), .A2(new_n610_), .ZN(new_n624_));
  OAI21_X1  g423(.A(KEYINPUT76), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT76), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n611_), .A2(new_n626_), .A3(new_n616_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n625_), .A2(new_n627_), .A3(new_n619_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(new_n617_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT37), .ZN(new_n630_));
  AOI211_X1 g429(.A(new_n600_), .B(new_n622_), .C1(new_n629_), .C2(new_n630_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n583_), .A2(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n632_), .A2(new_n549_), .A3(new_n502_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT38), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n296_), .A2(new_n580_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n629_), .B(KEYINPUT106), .ZN(new_n637_));
  NOR3_X1   g436(.A1(new_n548_), .A2(new_n600_), .A3(new_n637_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n636_), .A2(new_n638_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n549_), .B1(new_n639_), .B2(new_n502_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n635_), .A2(new_n640_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n641_), .B1(new_n634_), .B2(new_n633_), .ZN(G1324gat));
  INV_X1    g441(.A(new_n509_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n632_), .A2(new_n550_), .A3(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT39), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n639_), .A2(new_n643_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n645_), .B1(new_n646_), .B2(G8gat), .ZN(new_n647_));
  AOI211_X1 g446(.A(KEYINPUT39), .B(new_n550_), .C1(new_n639_), .C2(new_n643_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n644_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT40), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(G1325gat));
  INV_X1    g450(.A(G15gat), .ZN(new_n652_));
  INV_X1    g451(.A(new_n477_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n632_), .A2(new_n652_), .A3(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n652_), .B1(new_n639_), .B2(new_n653_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT108), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n656_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(KEYINPUT107), .B(KEYINPUT41), .ZN(new_n659_));
  AND3_X1   g458(.A1(new_n657_), .A2(new_n658_), .A3(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n659_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n654_), .B1(new_n660_), .B2(new_n661_), .ZN(G1326gat));
  INV_X1    g461(.A(new_n456_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n554_), .B1(new_n639_), .B2(new_n663_), .ZN(new_n664_));
  XOR2_X1   g463(.A(new_n664_), .B(KEYINPUT42), .Z(new_n665_));
  NAND2_X1  g464(.A1(new_n663_), .A2(new_n554_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT109), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n632_), .A2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n665_), .A2(new_n668_), .ZN(G1327gat));
  INV_X1    g468(.A(new_n600_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n629_), .A2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n583_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(G29gat), .B1(new_n673_), .B2(new_n502_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n580_), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n292_), .A2(new_n295_), .A3(new_n600_), .A4(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT43), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n510_), .A2(new_n506_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n528_), .A2(new_n502_), .A3(new_n532_), .ZN(new_n680_));
  AOI22_X1  g479(.A1(new_n680_), .A2(new_n511_), .B1(new_n541_), .B2(new_n540_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n663_), .B1(new_n681_), .B2(new_n533_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n477_), .B1(new_n682_), .B2(new_n545_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n679_), .A2(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n622_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n678_), .B1(new_n684_), .B2(new_n686_), .ZN(new_n687_));
  AOI211_X1 g486(.A(KEYINPUT43), .B(new_n685_), .C1(new_n679_), .C2(new_n683_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n677_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  AND3_X1   g490(.A1(new_n691_), .A2(G29gat), .A3(new_n502_), .ZN(new_n692_));
  OAI21_X1  g491(.A(KEYINPUT43), .B1(new_n548_), .B2(new_n685_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n684_), .A2(new_n678_), .A3(new_n686_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n695_), .A2(KEYINPUT44), .A3(new_n677_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n674_), .B1(new_n692_), .B2(new_n696_), .ZN(G1328gat));
  NOR2_X1   g496(.A1(new_n509_), .A2(G36gat), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n583_), .A2(new_n671_), .A3(new_n698_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT45), .Z(new_n700_));
  AOI21_X1  g499(.A(new_n676_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n643_), .B1(new_n701_), .B2(KEYINPUT44), .ZN(new_n702_));
  AOI211_X1 g501(.A(new_n690_), .B(new_n676_), .C1(new_n693_), .C2(new_n694_), .ZN(new_n703_));
  OAI211_X1 g502(.A(KEYINPUT110), .B(G36gat), .C1(new_n702_), .C2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n691_), .A2(new_n643_), .A3(new_n696_), .ZN(new_n706_));
  AOI21_X1  g505(.A(KEYINPUT110), .B1(new_n706_), .B2(G36gat), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n700_), .B1(new_n705_), .B2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT46), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  OAI211_X1 g509(.A(new_n700_), .B(KEYINPUT46), .C1(new_n705_), .C2(new_n707_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1329gat));
  NAND3_X1  g511(.A1(new_n583_), .A2(new_n653_), .A3(new_n671_), .ZN(new_n713_));
  INV_X1    g512(.A(G43gat), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT112), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n715_), .B(new_n716_), .ZN(new_n717_));
  AOI211_X1 g516(.A(new_n714_), .B(new_n477_), .C1(new_n689_), .C2(new_n690_), .ZN(new_n718_));
  AOI21_X1  g517(.A(KEYINPUT111), .B1(new_n718_), .B2(new_n696_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n477_), .A2(new_n714_), .ZN(new_n720_));
  AND4_X1   g519(.A1(KEYINPUT111), .A2(new_n691_), .A3(new_n696_), .A4(new_n720_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n717_), .B1(new_n719_), .B2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(KEYINPUT47), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT47), .ZN(new_n724_));
  OAI211_X1 g523(.A(new_n717_), .B(new_n724_), .C1(new_n719_), .C2(new_n721_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(G1330gat));
  AOI21_X1  g525(.A(G50gat), .B1(new_n673_), .B2(new_n663_), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n691_), .A2(G50gat), .A3(new_n663_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n727_), .B1(new_n728_), .B2(new_n696_), .ZN(G1331gat));
  INV_X1    g528(.A(new_n502_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n675_), .B1(new_n292_), .B2(new_n295_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n731_), .A2(new_n684_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(new_n631_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n730_), .B1(new_n733_), .B2(KEYINPUT113), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n734_), .B1(KEYINPUT113), .B2(new_n733_), .ZN(new_n735_));
  INV_X1    g534(.A(G57gat), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n638_), .A2(new_n296_), .A3(new_n582_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n730_), .A2(new_n736_), .ZN(new_n738_));
  AOI22_X1  g537(.A1(new_n735_), .A2(new_n736_), .B1(new_n737_), .B2(new_n738_), .ZN(G1332gat));
  INV_X1    g538(.A(G64gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(new_n737_), .B2(new_n643_), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n741_), .B(KEYINPUT48), .Z(new_n742_));
  INV_X1    g541(.A(new_n733_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n743_), .A2(new_n740_), .A3(new_n643_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(G1333gat));
  INV_X1    g544(.A(G71gat), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n746_), .B1(new_n737_), .B2(new_n653_), .ZN(new_n747_));
  XOR2_X1   g546(.A(new_n747_), .B(KEYINPUT49), .Z(new_n748_));
  NOR2_X1   g547(.A1(new_n477_), .A2(G71gat), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT114), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n748_), .B1(new_n733_), .B2(new_n750_), .ZN(G1334gat));
  INV_X1    g550(.A(G78gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n752_), .B1(new_n737_), .B2(new_n663_), .ZN(new_n753_));
  XOR2_X1   g552(.A(new_n753_), .B(KEYINPUT50), .Z(new_n754_));
  NAND3_X1  g553(.A1(new_n743_), .A2(new_n752_), .A3(new_n663_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(G1335gat));
  AND2_X1   g555(.A1(new_n732_), .A2(new_n671_), .ZN(new_n757_));
  AOI21_X1  g556(.A(G85gat), .B1(new_n757_), .B2(new_n502_), .ZN(new_n758_));
  OR2_X1    g557(.A1(new_n695_), .A2(KEYINPUT115), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n695_), .A2(KEYINPUT115), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n731_), .A2(new_n600_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n759_), .A2(new_n760_), .A3(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n502_), .A2(G85gat), .ZN(new_n764_));
  XOR2_X1   g563(.A(new_n764_), .B(KEYINPUT116), .Z(new_n765_));
  AOI21_X1  g564(.A(new_n758_), .B1(new_n763_), .B2(new_n765_), .ZN(G1336gat));
  AOI21_X1  g565(.A(G92gat), .B1(new_n757_), .B2(new_n643_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n509_), .A2(new_n298_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n763_), .B2(new_n768_), .ZN(G1337gat));
  OAI21_X1  g568(.A(G99gat), .B1(new_n762_), .B2(new_n477_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n757_), .A2(new_n242_), .A3(new_n653_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT51), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT51), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n770_), .A2(new_n774_), .A3(new_n771_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(G1338gat));
  NOR2_X1   g575(.A1(new_n456_), .A2(G106gat), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n757_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT117), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n757_), .A2(KEYINPUT117), .A3(new_n777_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n761_), .A2(new_n695_), .A3(new_n663_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n784_));
  AND3_X1   g583(.A1(new_n783_), .A2(new_n784_), .A3(G106gat), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n784_), .B1(new_n783_), .B2(G106gat), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n782_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(KEYINPUT53), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT53), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n782_), .B(new_n789_), .C1(new_n785_), .C2(new_n786_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n790_), .ZN(G1339gat));
  INV_X1    g590(.A(G113gat), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n581_), .B1(new_n294_), .B2(new_n289_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(new_n631_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(KEYINPUT118), .B(KEYINPUT54), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n794_), .B(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT55), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n278_), .A2(new_n251_), .A3(new_n262_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n203_), .ZN(new_n800_));
  AOI22_X1  g599(.A1(new_n281_), .A2(new_n798_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n275_), .A2(KEYINPUT55), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n271_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(KEYINPUT119), .A2(KEYINPUT56), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n287_), .B(new_n675_), .C1(new_n803_), .C2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n801_), .A2(new_n802_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n807_), .A2(new_n274_), .A3(new_n804_), .ZN(new_n808_));
  AOI21_X1  g607(.A(KEYINPUT120), .B1(new_n806_), .B2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n251_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n800_), .B1(new_n264_), .B2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n811_), .B1(new_n275_), .B2(KEYINPUT55), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n281_), .A2(new_n798_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n274_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n804_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n580_), .B1(new_n284_), .B2(new_n286_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n816_), .A2(KEYINPUT120), .A3(new_n808_), .A4(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n570_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n569_), .A2(new_n819_), .A3(new_n571_), .A4(new_n572_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n577_), .B1(new_n565_), .B2(new_n570_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n578_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n293_), .A2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n818_), .A2(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n629_), .B1(new_n809_), .B2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT57), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT120), .ZN(new_n828_));
  INV_X1    g627(.A(new_n808_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n828_), .B1(new_n805_), .B2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n830_), .A2(new_n823_), .A3(new_n818_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n831_), .A2(KEYINPUT57), .A3(new_n629_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT58), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT56), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n803_), .A2(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n835_), .A2(new_n287_), .A3(new_n822_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n814_), .A2(KEYINPUT56), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n833_), .B1(new_n836_), .B2(new_n838_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n287_), .A2(new_n822_), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n840_), .A2(KEYINPUT58), .A3(new_n837_), .A4(new_n835_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n839_), .A2(new_n686_), .A3(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n827_), .A2(new_n832_), .A3(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n797_), .B1(new_n843_), .B2(new_n600_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  NOR4_X1   g644(.A1(new_n643_), .A2(new_n730_), .A3(new_n663_), .A4(new_n477_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n792_), .B1(new_n847_), .B2(new_n580_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n846_), .ZN(new_n849_));
  OAI21_X1  g648(.A(KEYINPUT59), .B1(new_n844_), .B2(new_n849_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n582_), .A2(new_n792_), .ZN(new_n851_));
  AOI21_X1  g650(.A(KEYINPUT57), .B1(new_n831_), .B2(new_n629_), .ZN(new_n852_));
  AND3_X1   g651(.A1(new_n839_), .A2(new_n686_), .A3(new_n841_), .ZN(new_n853_));
  OAI21_X1  g652(.A(KEYINPUT122), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT122), .ZN(new_n855_));
  INV_X1    g654(.A(new_n629_), .ZN(new_n856_));
  AND2_X1   g655(.A1(new_n818_), .A2(new_n823_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n856_), .B1(new_n857_), .B2(new_n830_), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n855_), .B(new_n842_), .C1(new_n858_), .C2(KEYINPUT57), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n854_), .A2(new_n859_), .A3(new_n832_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n797_), .B1(new_n860_), .B2(new_n600_), .ZN(new_n861_));
  AOI21_X1  g660(.A(KEYINPUT59), .B1(new_n849_), .B2(KEYINPUT121), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n862_), .B1(KEYINPUT121), .B2(new_n849_), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n850_), .B(new_n851_), .C1(new_n861_), .C2(new_n863_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n848_), .A2(new_n864_), .ZN(G1340gat));
  OAI211_X1 g664(.A(new_n850_), .B(new_n296_), .C1(new_n861_), .C2(new_n863_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(G120gat), .ZN(new_n867_));
  INV_X1    g666(.A(G120gat), .ZN(new_n868_));
  INV_X1    g667(.A(new_n296_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n868_), .B1(new_n869_), .B2(KEYINPUT60), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n870_), .B1(KEYINPUT60), .B2(new_n868_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n867_), .B1(new_n847_), .B2(new_n871_), .ZN(G1341gat));
  INV_X1    g671(.A(G127gat), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n873_), .B1(new_n847_), .B2(new_n600_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n600_), .A2(new_n873_), .ZN(new_n875_));
  OAI211_X1 g674(.A(new_n850_), .B(new_n875_), .C1(new_n861_), .C2(new_n863_), .ZN(new_n876_));
  AND2_X1   g675(.A1(new_n874_), .A2(new_n876_), .ZN(G1342gat));
  INV_X1    g676(.A(G134gat), .ZN(new_n878_));
  INV_X1    g677(.A(new_n637_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n847_), .B2(new_n879_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n685_), .A2(new_n878_), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n850_), .B(new_n881_), .C1(new_n861_), .C2(new_n863_), .ZN(new_n882_));
  AND2_X1   g681(.A1(new_n880_), .A2(new_n882_), .ZN(G1343gat));
  NOR2_X1   g682(.A1(new_n653_), .A2(new_n456_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n509_), .A2(new_n502_), .A3(new_n884_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(KEYINPUT123), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(KEYINPUT124), .B1(new_n844_), .B2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT124), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n852_), .A2(new_n853_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n670_), .B1(new_n890_), .B2(new_n832_), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n889_), .B(new_n886_), .C1(new_n891_), .C2(new_n797_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n580_), .B1(new_n888_), .B2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(G141gat), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n893_), .B(new_n894_), .ZN(G1344gat));
  AOI21_X1  g694(.A(new_n869_), .B1(new_n888_), .B2(new_n892_), .ZN(new_n896_));
  INV_X1    g695(.A(G148gat), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n896_), .B(new_n897_), .ZN(G1345gat));
  AOI21_X1  g697(.A(new_n600_), .B1(new_n888_), .B2(new_n892_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(KEYINPUT61), .B(G155gat), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n899_), .B(new_n901_), .ZN(G1346gat));
  NAND2_X1  g701(.A1(new_n888_), .A2(new_n892_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n637_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n686_), .A2(G162gat), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(KEYINPUT125), .ZN(new_n906_));
  AOI22_X1  g705(.A1(new_n904_), .A2(new_n416_), .B1(new_n903_), .B2(new_n906_), .ZN(G1347gat));
  INV_X1    g706(.A(KEYINPUT62), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n643_), .A2(new_n456_), .A3(new_n503_), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n861_), .A2(new_n580_), .A3(new_n909_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n908_), .B1(new_n910_), .B2(new_n324_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n860_), .A2(new_n600_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n797_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n909_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n914_), .A2(new_n675_), .A3(new_n915_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n916_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n910_), .A2(new_n306_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n911_), .A2(new_n917_), .A3(new_n918_), .ZN(G1348gat));
  NOR2_X1   g718(.A1(new_n861_), .A2(new_n909_), .ZN(new_n920_));
  AOI21_X1  g719(.A(G176gat), .B1(new_n920_), .B2(new_n296_), .ZN(new_n921_));
  NOR3_X1   g720(.A1(new_n869_), .A2(new_n307_), .A3(new_n909_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n921_), .B1(new_n845_), .B2(new_n922_), .ZN(G1349gat));
  NAND2_X1  g722(.A1(new_n915_), .A2(new_n670_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n924_), .ZN(new_n925_));
  AOI21_X1  g724(.A(G183gat), .B1(new_n797_), .B2(new_n925_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n600_), .A2(new_n365_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n926_), .B1(new_n920_), .B2(new_n927_), .ZN(G1350gat));
  NAND2_X1  g727(.A1(new_n914_), .A2(new_n915_), .ZN(new_n929_));
  OAI21_X1  g728(.A(G190gat), .B1(new_n929_), .B2(new_n685_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n637_), .A2(new_n335_), .A3(new_n339_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n930_), .B1(new_n929_), .B2(new_n931_), .ZN(G1351gat));
  NAND2_X1  g731(.A1(new_n884_), .A2(new_n730_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(KEYINPUT126), .ZN(new_n934_));
  NOR3_X1   g733(.A1(new_n844_), .A2(new_n509_), .A3(new_n934_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(new_n675_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n936_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g736(.A1(new_n934_), .A2(new_n509_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n845_), .A2(new_n296_), .A3(new_n938_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n940_));
  AND2_X1   g739(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n941_));
  NOR3_X1   g740(.A1(new_n939_), .A2(new_n940_), .A3(new_n941_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n942_), .B1(new_n939_), .B2(new_n940_), .ZN(G1353gat));
  NOR2_X1   g742(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n944_));
  AND2_X1   g743(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n945_));
  OAI211_X1 g744(.A(new_n935_), .B(new_n670_), .C1(new_n944_), .C2(new_n945_), .ZN(new_n946_));
  INV_X1    g745(.A(new_n935_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n947_), .A2(new_n600_), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n946_), .B1(new_n948_), .B2(new_n944_), .ZN(G1354gat));
  AND3_X1   g748(.A1(new_n935_), .A2(G218gat), .A3(new_n686_), .ZN(new_n950_));
  AOI21_X1  g749(.A(G218gat), .B1(new_n935_), .B2(new_n637_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n950_), .A2(new_n951_), .ZN(G1355gat));
endmodule


