//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 1 0 0 0 0 0 0 1 1 1 0 0 0 0 1 0 1 0 0 1 1 1 0 0 0 0 1 1 1 0 0 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n671_,
    new_n672_, new_n673_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n757_, new_n758_,
    new_n759_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n770_, new_n771_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n885_, new_n886_, new_n888_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n913_, new_n914_, new_n915_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n922_, new_n923_, new_n924_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n932_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_, new_n943_;
  NOR2_X1   g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT78), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT78), .ZN(new_n204_));
  OAI21_X1  g003(.A(new_n204_), .B1(G169gat), .B2(G176gat), .ZN(new_n205_));
  AOI21_X1  g004(.A(KEYINPUT24), .B1(new_n203_), .B2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT25), .B(G183gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT77), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT26), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n208_), .B1(new_n209_), .B2(G190gat), .ZN(new_n210_));
  AND2_X1   g009(.A1(new_n207_), .A2(new_n210_), .ZN(new_n211_));
  XOR2_X1   g010(.A(KEYINPUT26), .B(G190gat), .Z(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT77), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n206_), .B1(new_n211_), .B2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(KEYINPUT79), .A2(G169gat), .A3(G176gat), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  AOI21_X1  g015(.A(KEYINPUT79), .B1(G169gat), .B2(G176gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n203_), .A2(new_n205_), .A3(KEYINPUT24), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT80), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  AND2_X1   g020(.A1(new_n203_), .A2(new_n205_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT80), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n222_), .A2(new_n223_), .A3(new_n218_), .A4(KEYINPUT24), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT23), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(KEYINPUT81), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT81), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n228_), .A2(G183gat), .A3(G190gat), .ZN(new_n229_));
  AND2_X1   g028(.A1(new_n227_), .A2(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n226_), .B1(new_n230_), .B2(KEYINPUT23), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n214_), .A2(new_n221_), .A3(new_n224_), .A4(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n227_), .A2(new_n229_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n233_), .B1(new_n234_), .B2(KEYINPUT23), .ZN(new_n235_));
  OR2_X1    g034(.A1(G183gat), .A2(G190gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(KEYINPUT22), .B(G169gat), .ZN(new_n238_));
  INV_X1    g037(.A(G176gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n237_), .A2(new_n218_), .A3(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n232_), .A2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT30), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G227gat), .A2(G233gat), .ZN(new_n244_));
  XOR2_X1   g043(.A(new_n243_), .B(new_n244_), .Z(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT31), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G15gat), .B(G43gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT82), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G71gat), .B(G99gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G127gat), .B(G134gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G113gat), .B(G120gat), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n251_), .B(new_n252_), .Z(new_n253_));
  XNOR2_X1  g052(.A(new_n250_), .B(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n246_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT31), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n245_), .B(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n254_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  AND2_X1   g058(.A1(new_n255_), .A2(new_n259_), .ZN(new_n260_));
  XOR2_X1   g059(.A(G57gat), .B(G85gat), .Z(new_n261_));
  XNOR2_X1  g060(.A(G1gat), .B(G29gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n261_), .B(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT92), .B(KEYINPUT0), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G225gat), .A2(G233gat), .ZN(new_n267_));
  NOR2_X1   g066(.A1(G155gat), .A2(G162gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G155gat), .A2(G162gat), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n268_), .B1(KEYINPUT1), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT83), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT1), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n271_), .A2(new_n272_), .A3(G155gat), .A4(G162gat), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT83), .B1(new_n269_), .B2(KEYINPUT1), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n270_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(G141gat), .A2(G148gat), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G141gat), .A2(G148gat), .ZN(new_n278_));
  AND2_X1   g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  AND2_X1   g078(.A1(new_n275_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n269_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n281_), .A2(new_n268_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n276_), .B(KEYINPUT3), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n278_), .B(KEYINPUT2), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n283_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n253_), .B1(new_n280_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n284_), .A2(new_n285_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(new_n282_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n251_), .B(new_n252_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n275_), .A2(new_n279_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n289_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n287_), .A2(new_n292_), .A3(KEYINPUT4), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT91), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT4), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n290_), .B1(new_n289_), .B2(new_n291_), .ZN(new_n296_));
  AOI22_X1  g095(.A1(new_n293_), .A2(new_n294_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n287_), .A2(new_n292_), .A3(KEYINPUT91), .A4(KEYINPUT4), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n267_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n287_), .A2(new_n292_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n267_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n266_), .B1(new_n299_), .B2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n293_), .A2(new_n294_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n296_), .A2(new_n295_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n304_), .A2(new_n298_), .A3(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(new_n301_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n302_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n307_), .A2(new_n265_), .A3(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n303_), .A2(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n260_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT99), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G8gat), .B(G36gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT18), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(G64gat), .ZN(new_n315_));
  XOR2_X1   g114(.A(new_n315_), .B(G92gat), .Z(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G211gat), .B(G218gat), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT21), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(G204gat), .ZN(new_n321_));
  OAI21_X1  g120(.A(KEYINPUT85), .B1(new_n321_), .B2(G197gat), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT85), .ZN(new_n323_));
  INV_X1    g122(.A(G197gat), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n323_), .A2(new_n324_), .A3(G204gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n321_), .A2(G197gat), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n322_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n320_), .A2(new_n327_), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n322_), .A2(new_n325_), .A3(new_n319_), .A4(new_n326_), .ZN(new_n329_));
  AND2_X1   g128(.A1(new_n329_), .A2(new_n318_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G197gat), .B(G204gat), .ZN(new_n331_));
  OAI21_X1  g130(.A(KEYINPUT84), .B1(new_n331_), .B2(new_n319_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n324_), .A2(G204gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n326_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT84), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n334_), .A2(new_n335_), .A3(KEYINPUT21), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n332_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT86), .ZN(new_n338_));
  AND3_X1   g137(.A1(new_n330_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n338_), .B1(new_n330_), .B2(new_n337_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n328_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  OR3_X1    g140(.A1(new_n216_), .A2(KEYINPUT89), .A3(new_n217_), .ZN(new_n342_));
  OAI21_X1  g141(.A(KEYINPUT89), .B1(new_n216_), .B2(new_n217_), .ZN(new_n343_));
  AND3_X1   g142(.A1(new_n342_), .A2(new_n240_), .A3(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n231_), .A2(new_n236_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT26), .B(G190gat), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT24), .ZN(new_n348_));
  AOI22_X1  g147(.A1(new_n347_), .A2(new_n207_), .B1(new_n348_), .B2(new_n202_), .ZN(new_n349_));
  AND2_X1   g148(.A1(new_n235_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G169gat), .A2(G176gat), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n222_), .A2(KEYINPUT24), .A3(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n346_), .A2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT20), .B1(new_n341_), .B2(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n335_), .B1(new_n334_), .B2(KEYINPUT21), .ZN(new_n356_));
  AOI211_X1 g155(.A(KEYINPUT84), .B(new_n319_), .C1(new_n326_), .C2(new_n333_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n329_), .A2(new_n318_), .ZN(new_n359_));
  OAI21_X1  g158(.A(KEYINPUT86), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n330_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  AOI22_X1  g161(.A1(new_n362_), .A2(new_n328_), .B1(new_n232_), .B2(new_n241_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G226gat), .A2(G233gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT19), .ZN(new_n365_));
  NOR3_X1   g164(.A1(new_n355_), .A2(new_n363_), .A3(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n365_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT20), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n368_), .B1(new_n341_), .B2(new_n354_), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n362_), .A2(new_n232_), .A3(new_n241_), .A4(new_n328_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n367_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n317_), .B1(new_n366_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n328_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n373_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n374_));
  AOI22_X1  g173(.A1(new_n345_), .A2(new_n344_), .B1(new_n350_), .B2(new_n352_), .ZN(new_n375_));
  OAI21_X1  g174(.A(KEYINPUT20), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n341_), .A2(new_n242_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n365_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n368_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n341_), .A2(new_n242_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n379_), .A2(new_n367_), .A3(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n378_), .A2(new_n316_), .A3(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n372_), .A2(KEYINPUT90), .A3(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT27), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT90), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n378_), .A2(new_n381_), .A3(new_n385_), .A4(new_n316_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n383_), .A2(new_n384_), .A3(new_n386_), .ZN(new_n387_));
  AND2_X1   g186(.A1(new_n382_), .A2(KEYINPUT27), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n365_), .B1(new_n355_), .B2(new_n363_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT95), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  OAI211_X1 g190(.A(KEYINPUT95), .B(new_n365_), .C1(new_n355_), .C2(new_n363_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n341_), .A2(new_n354_), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n370_), .A2(new_n393_), .A3(KEYINPUT20), .A4(new_n367_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(KEYINPUT96), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT96), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n369_), .A2(new_n396_), .A3(new_n367_), .A4(new_n370_), .ZN(new_n397_));
  AOI22_X1  g196(.A1(new_n391_), .A2(new_n392_), .B1(new_n395_), .B2(new_n397_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n388_), .B1(new_n398_), .B2(new_n316_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT98), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n387_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n400_), .B1(new_n387_), .B2(new_n399_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n289_), .A2(new_n291_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(KEYINPUT29), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n341_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(G228gat), .ZN(new_n407_));
  INV_X1    g206(.A(G233gat), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n406_), .A2(new_n409_), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n341_), .B(new_n405_), .C1(new_n407_), .C2(new_n408_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G78gat), .B(G106gat), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n410_), .A2(new_n411_), .A3(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT87), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n404_), .A2(KEYINPUT29), .ZN(new_n417_));
  XOR2_X1   g216(.A(G22gat), .B(G50gat), .Z(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(KEYINPUT28), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n417_), .B(new_n419_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n416_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n410_), .A2(new_n411_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(new_n412_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n423_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n421_), .A2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n423_), .A2(new_n414_), .A3(new_n420_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT88), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT88), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n423_), .A2(new_n414_), .A3(new_n428_), .A4(new_n420_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n425_), .A2(new_n427_), .A3(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n312_), .B1(new_n403_), .B2(new_n431_), .ZN(new_n432_));
  NOR4_X1   g231(.A1(new_n401_), .A2(new_n402_), .A3(KEYINPUT99), .A4(new_n430_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n311_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n310_), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n430_), .A2(new_n435_), .A3(new_n387_), .A4(new_n399_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n383_), .A2(new_n386_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n265_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT93), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n438_), .A2(new_n439_), .A3(KEYINPUT33), .ZN(new_n440_));
  OAI211_X1 g239(.A(KEYINPUT33), .B(new_n266_), .C1(new_n299_), .C2(new_n302_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT93), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n304_), .A2(new_n267_), .A3(new_n298_), .A4(new_n305_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n287_), .A2(new_n292_), .A3(new_n301_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(new_n265_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT94), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n444_), .A2(new_n265_), .A3(KEYINPUT94), .ZN(new_n448_));
  AND3_X1   g247(.A1(new_n443_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT33), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n449_), .B1(new_n303_), .B2(new_n450_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n437_), .A2(new_n440_), .A3(new_n442_), .A4(new_n451_), .ZN(new_n452_));
  AND2_X1   g251(.A1(new_n391_), .A2(new_n392_), .ZN(new_n453_));
  AND2_X1   g252(.A1(new_n395_), .A2(new_n397_), .ZN(new_n454_));
  OAI211_X1 g253(.A(KEYINPUT32), .B(new_n316_), .C1(new_n453_), .C2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n316_), .A2(KEYINPUT32), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n456_), .A2(new_n378_), .A3(new_n381_), .ZN(new_n457_));
  AND2_X1   g256(.A1(new_n310_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n455_), .A2(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n430_), .B1(new_n452_), .B2(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n436_), .B1(new_n460_), .B2(KEYINPUT97), .ZN(new_n461_));
  AND3_X1   g260(.A1(new_n451_), .A2(new_n440_), .A3(new_n442_), .ZN(new_n462_));
  AOI22_X1  g261(.A1(new_n462_), .A2(new_n437_), .B1(new_n455_), .B2(new_n458_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT97), .ZN(new_n464_));
  NOR3_X1   g263(.A1(new_n463_), .A2(new_n464_), .A3(new_n430_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n260_), .B1(new_n461_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n434_), .A2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(KEYINPUT74), .B(G8gat), .ZN(new_n468_));
  INV_X1    g267(.A(G1gat), .ZN(new_n469_));
  OAI21_X1  g268(.A(KEYINPUT14), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G15gat), .B(G22gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(G1gat), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n470_), .A2(new_n469_), .A3(new_n471_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(G8gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n473_), .A2(G8gat), .A3(new_n474_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  XOR2_X1   g278(.A(G29gat), .B(G36gat), .Z(new_n480_));
  XOR2_X1   g279(.A(G43gat), .B(G50gat), .Z(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n479_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G229gat), .A2(G233gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n482_), .B(KEYINPUT15), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n485_), .A2(new_n478_), .A3(new_n477_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n483_), .A2(new_n484_), .A3(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G113gat), .B(G141gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(G169gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(new_n324_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n482_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n477_), .A2(new_n478_), .A3(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n483_), .A2(KEYINPUT76), .A3(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(KEYINPUT76), .B1(new_n483_), .B2(new_n492_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n487_), .B(new_n490_), .C1(new_n496_), .C2(new_n484_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n490_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n483_), .A2(new_n492_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT76), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n484_), .B1(new_n501_), .B2(new_n493_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n487_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n498_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n497_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n467_), .A2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n479_), .B(KEYINPUT75), .ZN(new_n507_));
  AND2_X1   g306(.A1(G231gat), .A2(G233gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G71gat), .B(G78gat), .ZN(new_n511_));
  XOR2_X1   g310(.A(G57gat), .B(G64gat), .Z(new_n512_));
  INV_X1    g311(.A(KEYINPUT11), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n511_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G57gat), .B(G64gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT11), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n514_), .A2(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n515_), .A2(new_n511_), .A3(KEYINPUT11), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n510_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n519_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n509_), .A2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G127gat), .B(G155gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT16), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(G183gat), .ZN(new_n525_));
  XOR2_X1   g324(.A(new_n525_), .B(G211gat), .Z(new_n526_));
  INV_X1    g325(.A(KEYINPUT17), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n520_), .A2(new_n522_), .A3(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n519_), .B(KEYINPUT66), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n510_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT66), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n519_), .B(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n509_), .A2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n526_), .B(KEYINPUT17), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n531_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n529_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G190gat), .B(G218gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G134gat), .B(G162gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT36), .ZN(new_n542_));
  NOR2_X1   g341(.A1(G99gat), .A2(G106gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT7), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT8), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  XOR2_X1   g345(.A(KEYINPUT10), .B(G99gat), .Z(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(KEYINPUT64), .ZN(new_n548_));
  XNOR2_X1  g347(.A(KEYINPUT10), .B(G99gat), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT64), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(G106gat), .B1(new_n548_), .B2(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G85gat), .B(G92gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(KEYINPUT65), .B(KEYINPUT9), .ZN(new_n554_));
  OR2_X1    g353(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G85gat), .A2(G92gat), .ZN(new_n556_));
  OAI22_X1  g355(.A1(new_n553_), .A2(new_n554_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n546_), .B1(new_n552_), .B2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G99gat), .A2(G106gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT6), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n553_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n562_), .A2(KEYINPUT8), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n544_), .A2(new_n560_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n553_), .A2(new_n545_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n563_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n561_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT35), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G232gat), .A2(G233gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT71), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT34), .ZN(new_n571_));
  AOI22_X1  g370(.A1(new_n567_), .A2(new_n485_), .B1(new_n568_), .B2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n566_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n573_), .B1(new_n558_), .B2(new_n560_), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n574_), .A2(KEYINPUT72), .A3(new_n482_), .ZN(new_n575_));
  AOI21_X1  g374(.A(KEYINPUT72), .B1(new_n574_), .B2(new_n482_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n572_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n571_), .A2(new_n568_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  OAI221_X1 g378(.A(new_n572_), .B1(new_n568_), .B2(new_n571_), .C1(new_n575_), .C2(new_n576_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n542_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n579_), .A2(new_n580_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n541_), .A2(KEYINPUT36), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n582_), .A2(KEYINPUT73), .A3(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n579_), .A2(new_n580_), .A3(new_n583_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT73), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n581_), .B1(new_n584_), .B2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT37), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  AOI211_X1 g389(.A(KEYINPUT37), .B(new_n581_), .C1(new_n584_), .C2(new_n587_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n538_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G120gat), .B(G148gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(new_n321_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(KEYINPUT5), .B(G176gat), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n594_), .B(new_n595_), .Z(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n567_), .A2(KEYINPUT12), .A3(new_n521_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n533_), .A2(new_n574_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G230gat), .A2(G233gat), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT12), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n602_), .B1(new_n533_), .B2(new_n574_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n600_), .A2(new_n601_), .A3(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT67), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n605_), .B1(new_n533_), .B2(new_n574_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(new_n599_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n533_), .A2(new_n605_), .A3(new_n574_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n601_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT68), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n604_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  AOI211_X1 g410(.A(KEYINPUT68), .B(new_n601_), .C1(new_n607_), .C2(new_n608_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n597_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n601_), .ZN(new_n614_));
  AOI21_X1  g413(.A(KEYINPUT67), .B1(new_n530_), .B2(new_n567_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n530_), .A2(new_n567_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n608_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n614_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(KEYINPUT68), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n609_), .A2(new_n610_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n620_), .A2(new_n621_), .A3(new_n604_), .A4(new_n596_), .ZN(new_n622_));
  AND3_X1   g421(.A1(new_n613_), .A2(new_n622_), .A3(KEYINPUT69), .ZN(new_n623_));
  AOI21_X1  g422(.A(KEYINPUT69), .B1(new_n613_), .B2(new_n622_), .ZN(new_n624_));
  XOR2_X1   g423(.A(KEYINPUT70), .B(KEYINPUT13), .Z(new_n625_));
  OR3_X1    g424(.A1(new_n623_), .A2(new_n624_), .A3(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(KEYINPUT70), .A2(KEYINPUT13), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n627_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n592_), .B1(new_n626_), .B2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n506_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n632_), .A2(G1gat), .A3(new_n435_), .ZN(new_n633_));
  OR2_X1    g432(.A1(new_n633_), .A2(KEYINPUT38), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(KEYINPUT38), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n403_), .A2(new_n312_), .A3(new_n431_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n387_), .A2(new_n399_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(KEYINPUT98), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n387_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n638_), .A2(new_n431_), .A3(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(KEYINPUT99), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n636_), .A2(new_n641_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n464_), .B1(new_n463_), .B2(new_n430_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n452_), .A2(new_n459_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n644_), .A2(KEYINPUT97), .A3(new_n431_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n643_), .A2(new_n645_), .A3(new_n436_), .ZN(new_n646_));
  AOI22_X1  g445(.A1(new_n642_), .A2(new_n311_), .B1(new_n646_), .B2(new_n260_), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n647_), .A2(new_n537_), .A3(new_n588_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n626_), .A2(new_n628_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n505_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n648_), .A2(new_n652_), .ZN(new_n653_));
  OAI21_X1  g452(.A(G1gat), .B1(new_n653_), .B2(new_n435_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n634_), .A2(new_n635_), .A3(new_n654_), .ZN(G1324gat));
  INV_X1    g454(.A(new_n403_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n631_), .A2(new_n468_), .A3(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n648_), .A2(new_n656_), .A3(new_n652_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT39), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n658_), .A2(new_n659_), .A3(G8gat), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n659_), .B1(new_n658_), .B2(G8gat), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n657_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(KEYINPUT101), .ZN(new_n664_));
  XNOR2_X1  g463(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT101), .ZN(new_n666_));
  OAI211_X1 g465(.A(new_n666_), .B(new_n657_), .C1(new_n661_), .C2(new_n662_), .ZN(new_n667_));
  AND3_X1   g466(.A1(new_n664_), .A2(new_n665_), .A3(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n665_), .B1(new_n664_), .B2(new_n667_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n668_), .A2(new_n669_), .ZN(G1325gat));
  OAI21_X1  g469(.A(G15gat), .B1(new_n653_), .B2(new_n260_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT41), .ZN(new_n672_));
  NOR3_X1   g471(.A1(new_n632_), .A2(G15gat), .A3(new_n260_), .ZN(new_n673_));
  OR2_X1    g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1326gat));
  OR3_X1    g473(.A1(new_n632_), .A2(G22gat), .A3(new_n431_), .ZN(new_n675_));
  OAI21_X1  g474(.A(G22gat), .B1(new_n653_), .B2(new_n431_), .ZN(new_n676_));
  OR2_X1    g475(.A1(new_n676_), .A2(KEYINPUT102), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(KEYINPUT102), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n677_), .A2(KEYINPUT42), .A3(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(KEYINPUT42), .B1(new_n677_), .B2(new_n678_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n675_), .B1(new_n679_), .B2(new_n680_), .ZN(G1327gat));
  NAND2_X1  g480(.A1(new_n537_), .A2(new_n588_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT104), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n467_), .A2(new_n505_), .A3(new_n649_), .A4(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(G29gat), .B1(new_n685_), .B2(new_n310_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT103), .ZN(new_n687_));
  INV_X1    g486(.A(new_n588_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(KEYINPUT37), .ZN(new_n689_));
  INV_X1    g488(.A(new_n591_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n691_), .B1(new_n434_), .B2(new_n466_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT43), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n687_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  OAI211_X1 g493(.A(KEYINPUT103), .B(KEYINPUT43), .C1(new_n647_), .C2(new_n691_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n692_), .A2(new_n693_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n694_), .A2(new_n695_), .A3(new_n696_), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n650_), .A2(new_n651_), .A3(new_n538_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n697_), .A2(KEYINPUT44), .A3(new_n698_), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n699_), .A2(G29gat), .A3(new_n310_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n697_), .A2(new_n698_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n686_), .B1(new_n700_), .B2(new_n703_), .ZN(G1328gat));
  NAND2_X1  g503(.A1(new_n699_), .A2(new_n656_), .ZN(new_n705_));
  AOI21_X1  g504(.A(KEYINPUT44), .B1(new_n697_), .B2(new_n698_), .ZN(new_n706_));
  OAI21_X1  g505(.A(G36gat), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  NOR3_X1   g506(.A1(new_n684_), .A2(G36gat), .A3(new_n403_), .ZN(new_n708_));
  XOR2_X1   g507(.A(new_n708_), .B(KEYINPUT45), .Z(new_n709_));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n709_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(KEYINPUT105), .B(KEYINPUT46), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n710_), .B(new_n712_), .ZN(G1329gat));
  INV_X1    g512(.A(KEYINPUT47), .ZN(new_n714_));
  INV_X1    g513(.A(G43gat), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n715_), .B1(new_n684_), .B2(new_n260_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT106), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT107), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n260_), .A2(new_n715_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n699_), .A2(new_n719_), .ZN(new_n720_));
  OAI211_X1 g519(.A(new_n717_), .B(new_n718_), .C1(new_n720_), .C2(new_n706_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n703_), .A2(new_n699_), .A3(new_n719_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n718_), .B1(new_n723_), .B2(new_n717_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n714_), .B1(new_n722_), .B2(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n717_), .B1(new_n720_), .B2(new_n706_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT107), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n727_), .A2(KEYINPUT47), .A3(new_n721_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n725_), .A2(new_n728_), .ZN(G1330gat));
  NAND2_X1  g528(.A1(new_n699_), .A2(new_n430_), .ZN(new_n730_));
  OAI21_X1  g529(.A(G50gat), .B1(new_n730_), .B2(new_n706_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n431_), .A2(G50gat), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT108), .Z(new_n733_));
  OAI21_X1  g532(.A(new_n731_), .B1(new_n684_), .B2(new_n733_), .ZN(G1331gat));
  NAND3_X1  g533(.A1(new_n648_), .A2(new_n651_), .A3(new_n650_), .ZN(new_n735_));
  INV_X1    g534(.A(G57gat), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n735_), .A2(new_n736_), .A3(new_n435_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n537_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n650_), .A2(new_n738_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT109), .ZN(new_n740_));
  NOR3_X1   g539(.A1(new_n647_), .A2(KEYINPUT110), .A3(new_n505_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT110), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n742_), .B1(new_n467_), .B2(new_n651_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n740_), .B1(new_n741_), .B2(new_n743_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n736_), .B1(new_n744_), .B2(new_n435_), .ZN(new_n745_));
  OR2_X1    g544(.A1(new_n745_), .A2(KEYINPUT111), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(KEYINPUT111), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n737_), .B1(new_n746_), .B2(new_n747_), .ZN(G1332gat));
  OAI21_X1  g547(.A(G64gat), .B1(new_n735_), .B2(new_n403_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT48), .ZN(new_n750_));
  OR2_X1    g549(.A1(new_n403_), .A2(G64gat), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n750_), .B1(new_n744_), .B2(new_n751_), .ZN(G1333gat));
  OAI21_X1  g551(.A(G71gat), .B1(new_n735_), .B2(new_n260_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT49), .ZN(new_n754_));
  OR2_X1    g553(.A1(new_n260_), .A2(G71gat), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n754_), .B1(new_n744_), .B2(new_n755_), .ZN(G1334gat));
  OAI21_X1  g555(.A(G78gat), .B1(new_n735_), .B2(new_n431_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT50), .ZN(new_n758_));
  OR2_X1    g557(.A1(new_n431_), .A2(G78gat), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n758_), .B1(new_n744_), .B2(new_n759_), .ZN(G1335gat));
  NOR2_X1   g559(.A1(new_n741_), .A2(new_n743_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n683_), .A2(new_n650_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(G85gat), .B1(new_n763_), .B2(new_n310_), .ZN(new_n764_));
  NOR3_X1   g563(.A1(new_n649_), .A2(new_n505_), .A3(new_n538_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n697_), .A2(new_n765_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT112), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n310_), .A2(G85gat), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n764_), .B1(new_n767_), .B2(new_n768_), .ZN(G1336gat));
  AOI21_X1  g568(.A(G92gat), .B1(new_n763_), .B2(new_n656_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n656_), .A2(G92gat), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n767_), .B2(new_n771_), .ZN(G1337gat));
  OAI21_X1  g571(.A(G99gat), .B1(new_n766_), .B2(new_n260_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n260_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n548_), .A2(new_n551_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n763_), .A2(new_n774_), .A3(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n773_), .A2(new_n776_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g577(.A1(new_n697_), .A2(new_n430_), .A3(new_n765_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n779_), .A2(G106gat), .A3(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n780_), .B1(new_n779_), .B2(G106gat), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT114), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n782_), .A2(new_n783_), .A3(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n784_), .ZN(new_n786_));
  INV_X1    g585(.A(G106gat), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n763_), .A2(new_n787_), .A3(new_n430_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(KEYINPUT53), .B1(new_n785_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n783_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n791_), .A2(KEYINPUT114), .A3(new_n781_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n792_), .A2(new_n793_), .A3(new_n788_), .A4(new_n786_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n790_), .A2(new_n794_), .ZN(G1339gat));
  INV_X1    g594(.A(KEYINPUT54), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n629_), .A2(KEYINPUT115), .A3(new_n796_), .A4(new_n651_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n649_), .A2(new_n796_), .A3(new_n651_), .A4(new_n738_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT115), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n649_), .A2(new_n651_), .A3(new_n738_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT54), .ZN(new_n802_));
  AND3_X1   g601(.A1(new_n797_), .A2(new_n800_), .A3(new_n802_), .ZN(new_n803_));
  XNOR2_X1  g602(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT117), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n505_), .A2(new_n622_), .A3(KEYINPUT116), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n601_), .B1(new_n600_), .B2(new_n603_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT55), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n604_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n603_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n810_), .A2(new_n808_), .A3(new_n614_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n809_), .A2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT56), .B1(new_n813_), .B2(new_n597_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT56), .ZN(new_n815_));
  AOI211_X1 g614(.A(new_n815_), .B(new_n596_), .C1(new_n809_), .C2(new_n812_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n806_), .B1(new_n814_), .B2(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(KEYINPUT116), .B1(new_n505_), .B2(new_n622_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n805_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n813_), .A2(KEYINPUT56), .A3(new_n597_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n808_), .B1(new_n810_), .B2(new_n614_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n810_), .A2(new_n614_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n597_), .B1(new_n823_), .B2(new_n811_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n815_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n820_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n505_), .A2(new_n622_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT116), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n826_), .A2(new_n829_), .A3(KEYINPUT117), .A4(new_n806_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n623_), .A2(new_n624_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n484_), .B1(new_n479_), .B2(new_n482_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n490_), .B1(new_n832_), .B2(new_n486_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n484_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n833_), .B1(new_n496_), .B2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n497_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n831_), .A2(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n819_), .A2(new_n830_), .A3(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n804_), .B1(new_n839_), .B2(new_n688_), .ZN(new_n840_));
  AND2_X1   g639(.A1(new_n837_), .A2(new_n622_), .ZN(new_n841_));
  AND3_X1   g640(.A1(new_n841_), .A2(new_n826_), .A3(KEYINPUT58), .ZN(new_n842_));
  AOI21_X1  g641(.A(KEYINPUT58), .B1(new_n841_), .B2(new_n826_), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n691_), .A2(new_n842_), .A3(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(KEYINPUT119), .B1(new_n840_), .B2(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n839_), .A2(KEYINPUT57), .A3(new_n688_), .ZN(new_n846_));
  OR3_X1    g645(.A1(new_n691_), .A2(new_n842_), .A3(new_n843_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT119), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n826_), .A2(new_n829_), .A3(new_n806_), .ZN(new_n849_));
  AOI22_X1  g648(.A1(new_n849_), .A2(new_n805_), .B1(new_n831_), .B2(new_n837_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n588_), .B1(new_n850_), .B2(new_n830_), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n847_), .B(new_n848_), .C1(new_n851_), .C2(new_n804_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n845_), .A2(new_n846_), .A3(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n803_), .B1(new_n853_), .B2(new_n537_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n642_), .A2(new_n774_), .A3(new_n310_), .ZN(new_n855_));
  OR2_X1    g654(.A1(new_n855_), .A2(KEYINPUT59), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n846_), .B(new_n847_), .C1(new_n851_), .C2(new_n804_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n537_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n797_), .A2(new_n800_), .A3(new_n802_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n855_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT59), .ZN(new_n861_));
  OAI22_X1  g660(.A1(new_n854_), .A2(new_n856_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(G113gat), .B1(new_n862_), .B2(new_n651_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n860_), .ZN(new_n864_));
  OR2_X1    g663(.A1(new_n651_), .A2(G113gat), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n863_), .B1(new_n864_), .B2(new_n865_), .ZN(G1340gat));
  OAI21_X1  g665(.A(G120gat), .B1(new_n862_), .B2(new_n649_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT60), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(G120gat), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n649_), .A2(KEYINPUT60), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n869_), .B1(new_n870_), .B2(G120gat), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n867_), .B1(new_n864_), .B2(new_n871_), .ZN(G1341gat));
  OAI21_X1  g671(.A(G127gat), .B1(new_n862_), .B2(new_n537_), .ZN(new_n873_));
  OR2_X1    g672(.A1(new_n537_), .A2(G127gat), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n873_), .B1(new_n864_), .B2(new_n874_), .ZN(G1342gat));
  OAI21_X1  g674(.A(G134gat), .B1(new_n862_), .B2(new_n691_), .ZN(new_n876_));
  OR3_X1    g675(.A1(new_n864_), .A2(G134gat), .A3(new_n688_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(KEYINPUT120), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT120), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n876_), .A2(new_n880_), .A3(new_n877_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n881_), .ZN(G1343gat));
  NAND4_X1  g681(.A1(new_n260_), .A2(new_n430_), .A3(new_n403_), .A4(new_n310_), .ZN(new_n883_));
  XOR2_X1   g682(.A(new_n883_), .B(KEYINPUT121), .Z(new_n884_));
  AOI21_X1  g683(.A(new_n884_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n505_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g686(.A1(new_n885_), .A2(new_n650_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g688(.A1(new_n885_), .A2(new_n538_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(KEYINPUT61), .B(G155gat), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n890_), .B(new_n891_), .ZN(G1346gat));
  AOI21_X1  g691(.A(G162gat), .B1(new_n885_), .B2(new_n588_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n691_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(G162gat), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(KEYINPUT122), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n893_), .B1(new_n885_), .B2(new_n896_), .ZN(G1347gat));
  NAND3_X1  g696(.A1(new_n311_), .A2(new_n431_), .A3(new_n656_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n854_), .A2(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(new_n505_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(KEYINPUT123), .ZN(new_n901_));
  NOR4_X1   g700(.A1(new_n854_), .A2(KEYINPUT123), .A3(new_n651_), .A4(new_n898_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  NAND4_X1  g702(.A1(new_n901_), .A2(KEYINPUT62), .A3(new_n903_), .A4(G169gat), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT62), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n854_), .A2(new_n651_), .A3(new_n898_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT123), .ZN(new_n907_));
  OAI21_X1  g706(.A(G169gat), .B1(new_n906_), .B2(new_n907_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n905_), .B1(new_n908_), .B2(new_n902_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n906_), .A2(new_n238_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n904_), .A2(new_n909_), .A3(new_n910_), .ZN(G1348gat));
  AOI21_X1  g710(.A(new_n898_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n912_), .A2(G176gat), .A3(new_n650_), .ZN(new_n913_));
  XOR2_X1   g712(.A(new_n913_), .B(KEYINPUT124), .Z(new_n914_));
  AOI21_X1  g713(.A(G176gat), .B1(new_n899_), .B2(new_n650_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n914_), .A2(new_n915_), .ZN(G1349gat));
  NOR4_X1   g715(.A1(new_n854_), .A2(new_n207_), .A3(new_n537_), .A4(new_n898_), .ZN(new_n917_));
  AND2_X1   g716(.A1(new_n917_), .A2(KEYINPUT125), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n917_), .A2(KEYINPUT125), .ZN(new_n919_));
  AOI21_X1  g718(.A(G183gat), .B1(new_n912_), .B2(new_n538_), .ZN(new_n920_));
  NOR3_X1   g719(.A1(new_n918_), .A2(new_n919_), .A3(new_n920_), .ZN(G1350gat));
  NAND3_X1  g720(.A1(new_n899_), .A2(new_n347_), .A3(new_n588_), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n854_), .A2(new_n691_), .A3(new_n898_), .ZN(new_n923_));
  INV_X1    g722(.A(G190gat), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n922_), .B1(new_n923_), .B2(new_n924_), .ZN(G1351gat));
  NAND2_X1  g724(.A1(new_n858_), .A2(new_n859_), .ZN(new_n926_));
  NOR4_X1   g725(.A1(new_n774_), .A2(new_n431_), .A3(new_n310_), .A4(new_n403_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n926_), .A2(new_n927_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n928_), .A2(new_n651_), .ZN(new_n929_));
  XOR2_X1   g728(.A(KEYINPUT126), .B(G197gat), .Z(new_n930_));
  XNOR2_X1  g729(.A(new_n929_), .B(new_n930_), .ZN(G1352gat));
  NOR2_X1   g730(.A1(new_n928_), .A2(new_n649_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(new_n321_), .ZN(G1353gat));
  INV_X1    g732(.A(new_n928_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(new_n538_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n936_));
  AND2_X1   g735(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n937_));
  NOR3_X1   g736(.A1(new_n935_), .A2(new_n936_), .A3(new_n937_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n938_), .B1(new_n935_), .B2(new_n936_), .ZN(G1354gat));
  AND3_X1   g738(.A1(new_n934_), .A2(G218gat), .A3(new_n894_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n934_), .A2(new_n588_), .ZN(new_n941_));
  OR2_X1    g740(.A1(new_n941_), .A2(KEYINPUT127), .ZN(new_n942_));
  AOI21_X1  g741(.A(G218gat), .B1(new_n941_), .B2(KEYINPUT127), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n940_), .B1(new_n942_), .B2(new_n943_), .ZN(G1355gat));
endmodule


