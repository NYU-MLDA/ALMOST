//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 1 0 0 0 0 1 0 0 1 0 1 1 0 1 0 1 1 1 0 1 0 0 1 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 1 0 0 1 0 0 0 0 1 1 0 0 0 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n674_, new_n675_, new_n676_, new_n677_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n738_, new_n739_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n760_, new_n761_, new_n762_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n770_, new_n771_, new_n772_,
    new_n774_, new_n775_, new_n776_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n859_, new_n860_, new_n862_,
    new_n863_, new_n864_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n872_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n909_, new_n910_, new_n912_,
    new_n913_, new_n915_, new_n916_, new_n917_, new_n919_, new_n920_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(G169gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT22), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT22), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G169gat), .ZN(new_n206_));
  INV_X1    g005(.A(G176gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n204_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT82), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT82), .ZN(new_n211_));
  NAND4_X1  g010(.A1(new_n204_), .A2(new_n206_), .A3(new_n211_), .A4(new_n207_), .ZN(new_n212_));
  AND3_X1   g011(.A1(new_n209_), .A2(new_n210_), .A3(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT23), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT23), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n216_), .A2(G183gat), .A3(G190gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n215_), .A2(new_n217_), .A3(KEYINPUT83), .ZN(new_n218_));
  OR3_X1    g017(.A1(new_n214_), .A2(KEYINPUT83), .A3(KEYINPUT23), .ZN(new_n219_));
  INV_X1    g018(.A(G183gat), .ZN(new_n220_));
  INV_X1    g019(.A(G190gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n218_), .A2(new_n219_), .A3(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n220_), .A2(KEYINPUT25), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT25), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(G183gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n221_), .A2(KEYINPUT26), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT26), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(G190gat), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n224_), .A2(new_n226_), .A3(new_n227_), .A4(new_n229_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(G169gat), .A2(G176gat), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n232_), .A2(KEYINPUT24), .A3(new_n210_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT24), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n231_), .A2(new_n234_), .ZN(new_n235_));
  AND3_X1   g034(.A1(new_n230_), .A2(new_n233_), .A3(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT81), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n237_), .B1(new_n214_), .B2(KEYINPUT23), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n216_), .A2(KEYINPUT81), .A3(G183gat), .A4(G190gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n238_), .A2(new_n239_), .A3(new_n215_), .ZN(new_n240_));
  AOI22_X1  g039(.A1(new_n213_), .A2(new_n223_), .B1(new_n236_), .B2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT30), .ZN(new_n242_));
  OR2_X1    g041(.A1(new_n242_), .A2(KEYINPUT86), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G15gat), .B(G43gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT84), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(G71gat), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n246_), .A2(G99gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(G99gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G227gat), .A2(G233gat), .ZN(new_n249_));
  XOR2_X1   g048(.A(new_n249_), .B(KEYINPUT85), .Z(new_n250_));
  NAND3_X1  g049(.A1(new_n247_), .A2(new_n248_), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n247_), .A2(new_n248_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n250_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n243_), .A2(new_n251_), .A3(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT31), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT31), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n243_), .A2(new_n254_), .A3(new_n257_), .A4(new_n251_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n242_), .A2(KEYINPUT86), .ZN(new_n260_));
  OR2_X1    g059(.A1(new_n260_), .A2(KEYINPUT88), .ZN(new_n261_));
  INV_X1    g060(.A(G134gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(G127gat), .ZN(new_n263_));
  INV_X1    g062(.A(G127gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(G134gat), .ZN(new_n265_));
  INV_X1    g064(.A(G120gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(G113gat), .ZN(new_n267_));
  INV_X1    g066(.A(G113gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(G120gat), .ZN(new_n269_));
  AND4_X1   g068(.A1(new_n263_), .A2(new_n265_), .A3(new_n267_), .A4(new_n269_), .ZN(new_n270_));
  AOI22_X1  g069(.A1(new_n263_), .A2(new_n265_), .B1(new_n267_), .B2(new_n269_), .ZN(new_n271_));
  OAI21_X1  g070(.A(KEYINPUT87), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT87), .ZN(new_n273_));
  AND2_X1   g072(.A1(new_n263_), .A2(new_n265_), .ZN(new_n274_));
  AND2_X1   g073(.A1(new_n267_), .A2(new_n269_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n273_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n272_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n260_), .A2(KEYINPUT88), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n261_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n277_), .B1(new_n261_), .B2(new_n278_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n259_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n260_), .B(KEYINPUT88), .ZN(new_n283_));
  INV_X1    g082(.A(new_n277_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n285_), .A2(new_n256_), .A3(new_n258_), .A4(new_n279_), .ZN(new_n286_));
  AND2_X1   g085(.A1(new_n282_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT92), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G141gat), .A2(G148gat), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT89), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(KEYINPUT89), .A2(G141gat), .A3(G148gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  AND2_X1   g092(.A1(KEYINPUT91), .A2(KEYINPUT2), .ZN(new_n294_));
  NOR2_X1   g093(.A1(KEYINPUT91), .A2(KEYINPUT2), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n288_), .B1(new_n293_), .B2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(KEYINPUT91), .B(KEYINPUT2), .ZN(new_n298_));
  NAND4_X1  g097(.A1(new_n298_), .A2(KEYINPUT92), .A3(new_n291_), .A4(new_n292_), .ZN(new_n299_));
  INV_X1    g098(.A(G141gat), .ZN(new_n300_));
  INV_X1    g099(.A(G148gat), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n300_), .A2(new_n301_), .A3(KEYINPUT3), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT3), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n303_), .B1(G141gat), .B2(G148gat), .ZN(new_n304_));
  INV_X1    g103(.A(new_n289_), .ZN(new_n305_));
  AOI22_X1  g104(.A1(new_n302_), .A2(new_n304_), .B1(new_n305_), .B2(KEYINPUT2), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n297_), .A2(new_n299_), .A3(new_n306_), .ZN(new_n307_));
  OR2_X1    g106(.A1(G155gat), .A2(G162gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n307_), .A2(new_n310_), .ZN(new_n311_));
  AND2_X1   g110(.A1(new_n291_), .A2(new_n292_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n300_), .A2(new_n301_), .A3(KEYINPUT90), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT90), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n315_), .B1(G141gat), .B2(G148gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT1), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n308_), .A2(new_n318_), .A3(new_n309_), .ZN(new_n319_));
  AND4_X1   g118(.A1(new_n312_), .A2(new_n313_), .A3(new_n317_), .A4(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  OR2_X1    g120(.A1(new_n270_), .A2(new_n271_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n311_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G225gat), .A2(G233gat), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n320_), .B1(new_n307_), .B2(new_n310_), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n323_), .B(new_n324_), .C1(new_n325_), .C2(new_n277_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n277_), .B1(new_n311_), .B2(new_n321_), .ZN(new_n327_));
  XOR2_X1   g126(.A(KEYINPUT100), .B(KEYINPUT4), .Z(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n324_), .B1(new_n327_), .B2(new_n329_), .ZN(new_n330_));
  OAI211_X1 g129(.A(new_n323_), .B(KEYINPUT4), .C1(new_n325_), .C2(new_n277_), .ZN(new_n331_));
  AND3_X1   g130(.A1(new_n330_), .A2(new_n331_), .A3(KEYINPUT101), .ZN(new_n332_));
  AOI21_X1  g131(.A(KEYINPUT101), .B1(new_n330_), .B2(new_n331_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n326_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G1gat), .B(G29gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(G85gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT0), .B(G57gat), .ZN(new_n337_));
  XOR2_X1   g136(.A(new_n336_), .B(new_n337_), .Z(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n334_), .A2(new_n339_), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n326_), .B(new_n338_), .C1(new_n332_), .C2(new_n333_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n340_), .A2(KEYINPUT104), .A3(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT27), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G197gat), .A2(G204gat), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(G197gat), .A2(G204gat), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT21), .ZN(new_n348_));
  NOR3_X1   g147(.A1(new_n346_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G211gat), .B(G218gat), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(KEYINPUT95), .B1(new_n349_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(G197gat), .ZN(new_n353_));
  INV_X1    g152(.A(G204gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n355_), .A2(KEYINPUT21), .A3(new_n345_), .ZN(new_n356_));
  AOI21_X1  g155(.A(KEYINPUT21), .B1(new_n355_), .B2(new_n345_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT94), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n356_), .B(new_n350_), .C1(new_n357_), .C2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n355_), .A2(new_n345_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n360_), .A2(new_n358_), .A3(new_n348_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n352_), .B1(new_n359_), .B2(new_n362_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n349_), .A2(new_n351_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT95), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n365_), .B1(new_n356_), .B2(new_n350_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n348_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT94), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n364_), .A2(new_n366_), .A3(new_n361_), .A4(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n363_), .A2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n236_), .A2(new_n219_), .A3(new_n218_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n240_), .A2(new_n222_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(KEYINPUT98), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT98), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n240_), .A2(new_n374_), .A3(new_n222_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n204_), .A2(new_n206_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(KEYINPUT97), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT97), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n204_), .A2(new_n206_), .A3(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n377_), .A2(new_n379_), .A3(new_n207_), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n373_), .A2(new_n210_), .A3(new_n375_), .A4(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n370_), .A2(new_n371_), .A3(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n236_), .A2(new_n240_), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n223_), .A2(new_n210_), .A3(new_n212_), .A4(new_n209_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n385_), .A2(new_n369_), .A3(new_n363_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G226gat), .A2(G233gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(KEYINPUT19), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  AND4_X1   g188(.A1(KEYINPUT20), .A2(new_n382_), .A3(new_n386_), .A4(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n381_), .A2(new_n371_), .ZN(new_n391_));
  AND2_X1   g190(.A1(new_n363_), .A2(new_n369_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT20), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n394_), .B1(new_n370_), .B2(new_n241_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n389_), .B1(new_n393_), .B2(new_n395_), .ZN(new_n396_));
  XOR2_X1   g195(.A(G8gat), .B(G36gat), .Z(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(KEYINPUT18), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G64gat), .B(G92gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NOR3_X1   g200(.A1(new_n390_), .A2(new_n396_), .A3(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(KEYINPUT20), .B1(new_n392_), .B2(new_n385_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n370_), .B1(new_n371_), .B2(new_n381_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n388_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n394_), .B1(new_n392_), .B2(new_n385_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n406_), .A2(new_n389_), .A3(new_n382_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n400_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n344_), .B1(new_n402_), .B2(new_n408_), .ZN(new_n409_));
  NOR3_X1   g208(.A1(new_n403_), .A2(new_n404_), .A3(new_n388_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n389_), .B1(new_n406_), .B2(new_n382_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n401_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n405_), .A2(new_n407_), .A3(new_n400_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n412_), .A2(KEYINPUT27), .A3(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n311_), .A2(new_n321_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n370_), .B1(new_n415_), .B2(KEYINPUT29), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G228gat), .A2(G233gat), .ZN(new_n417_));
  INV_X1    g216(.A(G78gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n417_), .B(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(G106gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n416_), .B(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT96), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT29), .ZN(new_n423_));
  XOR2_X1   g222(.A(KEYINPUT93), .B(KEYINPUT28), .Z(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n325_), .A2(new_n423_), .A3(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  XOR2_X1   g226(.A(G22gat), .B(G50gat), .Z(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n425_), .B1(new_n325_), .B2(new_n423_), .ZN(new_n430_));
  NOR3_X1   g229(.A1(new_n427_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n424_), .B1(new_n415_), .B2(KEYINPUT29), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n428_), .B1(new_n432_), .B2(new_n426_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n421_), .B(new_n422_), .C1(new_n431_), .C2(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n422_), .B1(new_n431_), .B2(new_n433_), .ZN(new_n435_));
  XOR2_X1   g234(.A(new_n416_), .B(new_n420_), .Z(new_n436_));
  OAI21_X1  g235(.A(new_n429_), .B1(new_n427_), .B2(new_n430_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n432_), .A2(new_n428_), .A3(new_n426_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n437_), .A2(KEYINPUT96), .A3(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n435_), .A2(new_n436_), .A3(new_n439_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n409_), .A2(new_n414_), .A3(new_n434_), .A4(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(KEYINPUT104), .B1(new_n340_), .B2(new_n341_), .ZN(new_n442_));
  NOR3_X1   g241(.A1(new_n343_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  AND2_X1   g242(.A1(new_n440_), .A2(new_n434_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n330_), .A2(new_n331_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT101), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n330_), .A2(new_n331_), .A3(KEYINPUT101), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  AND3_X1   g248(.A1(new_n326_), .A2(KEYINPUT33), .A3(new_n338_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n324_), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n323_), .B(new_n451_), .C1(new_n325_), .C2(new_n277_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(new_n339_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n327_), .A2(new_n329_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n331_), .A2(new_n324_), .A3(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT103), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n453_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n331_), .A2(KEYINPUT103), .A3(new_n454_), .A4(new_n324_), .ZN(new_n458_));
  AOI22_X1  g257(.A1(new_n449_), .A2(new_n450_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  XOR2_X1   g258(.A(KEYINPUT102), .B(KEYINPUT33), .Z(new_n460_));
  NAND2_X1  g259(.A1(new_n341_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT99), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n462_), .B1(new_n402_), .B2(new_n408_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n401_), .B1(new_n390_), .B2(new_n396_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n464_), .A2(new_n413_), .A3(KEYINPUT99), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n459_), .A2(new_n461_), .A3(new_n463_), .A4(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n326_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n467_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n341_), .B1(new_n468_), .B2(new_n338_), .ZN(new_n469_));
  OAI211_X1 g268(.A(KEYINPUT32), .B(new_n400_), .C1(new_n410_), .C2(new_n411_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n400_), .A2(KEYINPUT32), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n405_), .A2(new_n407_), .A3(new_n471_), .ZN(new_n472_));
  AND2_X1   g271(.A1(new_n470_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n469_), .A2(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n444_), .B1(new_n466_), .B2(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n287_), .B1(new_n443_), .B2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT105), .ZN(new_n477_));
  INV_X1    g276(.A(new_n287_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n343_), .A2(new_n442_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n409_), .A2(new_n414_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n444_), .A2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n478_), .A2(new_n479_), .A3(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT105), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n287_), .B(new_n483_), .C1(new_n443_), .C2(new_n475_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n477_), .A2(new_n482_), .A3(new_n484_), .ZN(new_n485_));
  XOR2_X1   g284(.A(KEYINPUT10), .B(G99gat), .Z(new_n486_));
  INV_X1    g285(.A(G106gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  XOR2_X1   g287(.A(G85gat), .B(G92gat), .Z(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(KEYINPUT9), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G99gat), .A2(G106gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT6), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT6), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n493_), .A2(G99gat), .A3(G106gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(G85gat), .ZN(new_n496_));
  INV_X1    g295(.A(G92gat), .ZN(new_n497_));
  OR3_X1    g296(.A1(new_n496_), .A2(new_n497_), .A3(KEYINPUT9), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n488_), .A2(new_n490_), .A3(new_n495_), .A4(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT8), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n495_), .A2(KEYINPUT64), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT64), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n492_), .A2(new_n494_), .A3(new_n502_), .ZN(new_n503_));
  OAI21_X1  g302(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NOR3_X1   g304(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n501_), .A2(new_n503_), .A3(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n500_), .B1(new_n508_), .B2(new_n489_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n489_), .A2(new_n500_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n510_), .B1(new_n495_), .B2(new_n507_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n499_), .B1(new_n509_), .B2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(KEYINPUT65), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G29gat), .B(G36gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G43gat), .B(G50gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT65), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n517_), .B(new_n499_), .C1(new_n509_), .C2(new_n511_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n513_), .A2(new_n516_), .A3(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n516_), .B(KEYINPUT15), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT35), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G232gat), .A2(G233gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(KEYINPUT34), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  AOI22_X1  g323(.A1(new_n512_), .A2(new_n520_), .B1(new_n521_), .B2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n519_), .A2(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n524_), .A2(new_n521_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n527_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n519_), .A2(new_n529_), .A3(new_n525_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G190gat), .B(G218gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G134gat), .B(G162gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n534_), .A2(KEYINPUT36), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(KEYINPUT36), .ZN(new_n537_));
  AND2_X1   g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n531_), .A2(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n528_), .A2(new_n530_), .A3(new_n535_), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(KEYINPUT106), .B1(new_n485_), .B2(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G1gat), .B(G8gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT75), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G15gat), .B(G22gat), .ZN(new_n546_));
  INV_X1    g345(.A(G8gat), .ZN(new_n547_));
  OAI21_X1  g346(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n546_), .A2(new_n548_), .ZN(new_n549_));
  OR2_X1    g348(.A1(new_n545_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n545_), .A2(new_n549_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G231gat), .A2(G233gat), .ZN(new_n553_));
  XOR2_X1   g352(.A(new_n552_), .B(new_n553_), .Z(new_n554_));
  XNOR2_X1  g353(.A(G57gat), .B(G64gat), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(KEYINPUT11), .ZN(new_n556_));
  XOR2_X1   g355(.A(G71gat), .B(G78gat), .Z(new_n557_));
  OR2_X1    g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n556_), .A2(new_n557_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n555_), .A2(KEYINPUT11), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n558_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n561_), .B(KEYINPUT66), .Z(new_n562_));
  OR2_X1    g361(.A1(new_n554_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n554_), .A2(new_n562_), .ZN(new_n564_));
  XOR2_X1   g363(.A(G127gat), .B(G155gat), .Z(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT16), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G183gat), .B(G211gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT17), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n563_), .A2(new_n564_), .A3(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n561_), .B(KEYINPUT68), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n554_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT17), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n568_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n554_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n575_), .B1(new_n576_), .B2(new_n571_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n570_), .B1(new_n573_), .B2(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT76), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n543_), .A2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n485_), .A2(KEYINPUT106), .A3(new_n542_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n520_), .A2(new_n552_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT78), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n520_), .A2(new_n552_), .A3(KEYINPUT78), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n550_), .A2(new_n551_), .A3(new_n516_), .ZN(new_n588_));
  AND3_X1   g387(.A1(new_n586_), .A2(new_n587_), .A3(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(G229gat), .A2(G233gat), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n591_), .A2(KEYINPUT79), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(KEYINPUT79), .ZN(new_n593_));
  INV_X1    g392(.A(new_n516_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n552_), .A2(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n590_), .B1(new_n595_), .B2(new_n588_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT77), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n592_), .A2(new_n593_), .A3(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G113gat), .B(G141gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT80), .ZN(new_n600_));
  XOR2_X1   g399(.A(G169gat), .B(G197gat), .Z(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n598_), .B(new_n602_), .Z(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n572_), .A2(KEYINPUT12), .A3(new_n512_), .ZN(new_n605_));
  OR2_X1    g404(.A1(new_n605_), .A2(KEYINPUT69), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(KEYINPUT69), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n562_), .B1(new_n513_), .B2(new_n518_), .ZN(new_n608_));
  OAI211_X1 g407(.A(new_n606_), .B(new_n607_), .C1(KEYINPUT12), .C2(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n562_), .A2(new_n513_), .A3(new_n518_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(G230gat), .A2(G233gat), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT70), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n609_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n611_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n610_), .B(KEYINPUT67), .ZN(new_n616_));
  OR2_X1    g415(.A1(new_n616_), .A2(new_n608_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n614_), .B1(new_n615_), .B2(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G120gat), .B(G148gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT5), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G176gat), .B(G204gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n618_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n622_), .B(KEYINPUT71), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n618_), .A2(new_n626_), .ZN(new_n627_));
  OAI21_X1  g426(.A(KEYINPUT13), .B1(new_n624_), .B2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT13), .ZN(new_n629_));
  OAI211_X1 g428(.A(new_n623_), .B(new_n629_), .C1(new_n618_), .C2(new_n626_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n583_), .A2(new_n604_), .A3(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n479_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n202_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT107), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT74), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n540_), .A2(KEYINPUT72), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT72), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n528_), .A2(new_n639_), .A3(new_n530_), .A4(new_n535_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n638_), .A2(new_n539_), .A3(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT73), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n641_), .A2(new_n642_), .A3(KEYINPUT37), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT37), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n541_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n643_), .A2(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n642_), .B1(new_n641_), .B2(KEYINPUT37), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n637_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n641_), .A2(KEYINPUT37), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(KEYINPUT73), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n650_), .A2(KEYINPUT74), .A3(new_n645_), .A4(new_n643_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n648_), .A2(new_n651_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n652_), .A2(new_n580_), .ZN(new_n653_));
  AND4_X1   g452(.A1(new_n603_), .A2(new_n653_), .A3(new_n631_), .A4(new_n485_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n654_), .A2(new_n202_), .A3(new_n634_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT38), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n636_), .A2(new_n656_), .ZN(G1324gat));
  INV_X1    g456(.A(KEYINPUT108), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n633_), .A2(new_n480_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n658_), .B1(new_n659_), .B2(G8gat), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT39), .ZN(new_n661_));
  AOI21_X1  g460(.A(G8gat), .B1(new_n409_), .B2(new_n414_), .ZN(new_n662_));
  AOI22_X1  g461(.A1(new_n660_), .A2(new_n661_), .B1(new_n654_), .B2(new_n662_), .ZN(new_n663_));
  OR2_X1    g462(.A1(new_n660_), .A2(new_n661_), .ZN(new_n664_));
  AOI211_X1 g463(.A(KEYINPUT108), .B(new_n547_), .C1(new_n633_), .C2(new_n480_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n663_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(KEYINPUT109), .B(KEYINPUT40), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n666_), .B(new_n667_), .ZN(G1325gat));
  INV_X1    g467(.A(G15gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n669_), .B1(new_n633_), .B2(new_n478_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT41), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n654_), .A2(new_n669_), .A3(new_n478_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1326gat));
  INV_X1    g472(.A(G22gat), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n674_), .B1(new_n633_), .B2(new_n444_), .ZN(new_n675_));
  XOR2_X1   g474(.A(new_n675_), .B(KEYINPUT42), .Z(new_n676_));
  NAND3_X1  g475(.A1(new_n654_), .A2(new_n674_), .A3(new_n444_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(G1327gat));
  NOR2_X1   g477(.A1(new_n579_), .A2(new_n542_), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n631_), .A2(new_n603_), .A3(new_n485_), .A4(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(G29gat), .B1(new_n681_), .B2(new_n634_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT112), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n631_), .A2(new_n603_), .A3(new_n580_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT43), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n686_), .B1(new_n485_), .B2(new_n652_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n485_), .A2(new_n686_), .A3(new_n652_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(KEYINPUT110), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT110), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n485_), .A2(new_n652_), .A3(new_n690_), .A4(new_n686_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n685_), .B1(new_n689_), .B2(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n684_), .B1(new_n692_), .B2(KEYINPUT111), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n688_), .A2(KEYINPUT110), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n485_), .A2(new_n652_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(KEYINPUT43), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n694_), .A2(new_n691_), .A3(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n685_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n697_), .A2(KEYINPUT111), .A3(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n683_), .B1(new_n693_), .B2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n697_), .A2(new_n698_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT111), .ZN(new_n703_));
  AOI21_X1  g502(.A(KEYINPUT44), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n704_), .A2(KEYINPUT112), .A3(new_n699_), .ZN(new_n705_));
  AOI22_X1  g504(.A1(new_n701_), .A2(new_n705_), .B1(KEYINPUT44), .B2(new_n692_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n634_), .A2(G29gat), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n682_), .B1(new_n706_), .B2(new_n707_), .ZN(G1328gat));
  INV_X1    g507(.A(G36gat), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n681_), .A2(new_n709_), .A3(new_n480_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(KEYINPUT114), .B(KEYINPUT45), .ZN(new_n711_));
  XOR2_X1   g510(.A(new_n710_), .B(new_n711_), .Z(new_n712_));
  NAND2_X1  g511(.A1(new_n692_), .A2(KEYINPUT44), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(new_n480_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n714_), .B1(new_n701_), .B2(new_n705_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT113), .ZN(new_n716_));
  NOR3_X1   g515(.A1(new_n715_), .A2(new_n716_), .A3(new_n709_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n714_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n702_), .A2(new_n703_), .ZN(new_n719_));
  AND4_X1   g518(.A1(KEYINPUT112), .A2(new_n719_), .A3(new_n684_), .A4(new_n699_), .ZN(new_n720_));
  AOI21_X1  g519(.A(KEYINPUT112), .B1(new_n704_), .B2(new_n699_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n718_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(KEYINPUT113), .B1(new_n722_), .B2(G36gat), .ZN(new_n723_));
  OAI211_X1 g522(.A(KEYINPUT46), .B(new_n712_), .C1(new_n717_), .C2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n712_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n716_), .B1(new_n715_), .B2(new_n709_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n722_), .A2(KEYINPUT113), .A3(G36gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n725_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  XOR2_X1   g527(.A(KEYINPUT115), .B(KEYINPUT46), .Z(new_n729_));
  OAI21_X1  g528(.A(new_n724_), .B1(new_n728_), .B2(new_n729_), .ZN(G1329gat));
  INV_X1    g529(.A(G43gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n731_), .B1(new_n706_), .B2(new_n478_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT47), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n680_), .A2(G43gat), .A3(new_n287_), .ZN(new_n734_));
  OR3_X1    g533(.A1(new_n732_), .A2(new_n733_), .A3(new_n734_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n733_), .B1(new_n732_), .B2(new_n734_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(G1330gat));
  AOI21_X1  g536(.A(G50gat), .B1(new_n681_), .B2(new_n444_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n444_), .A2(G50gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n706_), .B2(new_n739_), .ZN(G1331gat));
  NOR3_X1   g539(.A1(new_n583_), .A2(new_n603_), .A3(new_n631_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(G57gat), .B1(new_n742_), .B2(new_n479_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n631_), .A2(new_n603_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n744_), .A2(new_n485_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n745_), .A2(new_n653_), .ZN(new_n746_));
  INV_X1    g545(.A(G57gat), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n746_), .A2(new_n747_), .A3(new_n634_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n743_), .A2(new_n748_), .ZN(G1332gat));
  INV_X1    g548(.A(G64gat), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n750_), .B1(new_n741_), .B2(new_n480_), .ZN(new_n751_));
  XOR2_X1   g550(.A(new_n751_), .B(KEYINPUT48), .Z(new_n752_));
  NAND3_X1  g551(.A1(new_n746_), .A2(new_n750_), .A3(new_n480_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(G1333gat));
  INV_X1    g553(.A(G71gat), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n755_), .B1(new_n741_), .B2(new_n478_), .ZN(new_n756_));
  XOR2_X1   g555(.A(new_n756_), .B(KEYINPUT49), .Z(new_n757_));
  NAND3_X1  g556(.A1(new_n746_), .A2(new_n755_), .A3(new_n478_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(G1334gat));
  AOI21_X1  g558(.A(new_n418_), .B1(new_n741_), .B2(new_n444_), .ZN(new_n760_));
  XOR2_X1   g559(.A(new_n760_), .B(KEYINPUT50), .Z(new_n761_));
  NAND3_X1  g560(.A1(new_n746_), .A2(new_n418_), .A3(new_n444_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(G1335gat));
  NAND2_X1  g562(.A1(new_n745_), .A2(new_n679_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n765_), .A2(new_n496_), .A3(new_n634_), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n697_), .A2(new_n580_), .A3(new_n744_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n767_), .A2(new_n634_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n766_), .B1(new_n768_), .B2(new_n496_), .ZN(G1336gat));
  AOI21_X1  g568(.A(new_n497_), .B1(new_n767_), .B2(new_n480_), .ZN(new_n770_));
  AOI21_X1  g569(.A(G92gat), .B1(new_n409_), .B2(new_n414_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n765_), .B2(new_n771_), .ZN(new_n772_));
  XOR2_X1   g571(.A(new_n772_), .B(KEYINPUT116), .Z(G1337gat));
  NAND2_X1  g572(.A1(new_n767_), .A2(new_n478_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n478_), .A2(new_n486_), .ZN(new_n775_));
  AOI22_X1  g574(.A1(new_n774_), .A2(G99gat), .B1(new_n765_), .B2(new_n775_), .ZN(new_n776_));
  XOR2_X1   g575(.A(new_n776_), .B(KEYINPUT51), .Z(G1338gat));
  NAND2_X1  g576(.A1(new_n767_), .A2(new_n444_), .ZN(new_n778_));
  AND3_X1   g577(.A1(new_n778_), .A2(KEYINPUT118), .A3(G106gat), .ZN(new_n779_));
  AOI21_X1  g578(.A(KEYINPUT118), .B1(new_n778_), .B2(G106gat), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT52), .ZN(new_n781_));
  OR3_X1    g580(.A1(new_n779_), .A2(new_n780_), .A3(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n765_), .A2(new_n487_), .A3(new_n444_), .ZN(new_n783_));
  OR2_X1    g582(.A1(new_n783_), .A2(KEYINPUT117), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(KEYINPUT117), .ZN(new_n785_));
  AOI22_X1  g584(.A1(new_n784_), .A2(new_n785_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n782_), .A2(new_n786_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n787_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g587(.A1(new_n653_), .A2(new_n604_), .A3(new_n631_), .ZN(new_n789_));
  XOR2_X1   g588(.A(new_n789_), .B(KEYINPUT54), .Z(new_n790_));
  NAND4_X1  g589(.A1(new_n592_), .A2(new_n593_), .A3(new_n597_), .A4(new_n602_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n595_), .A2(new_n588_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n602_), .B1(new_n792_), .B2(new_n590_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n589_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n793_), .B1(new_n794_), .B2(new_n590_), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n791_), .B(new_n795_), .C1(new_n624_), .C2(new_n627_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n603_), .A2(new_n623_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n614_), .A2(KEYINPUT55), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n615_), .B1(new_n609_), .B2(new_n616_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n801_), .B1(new_n609_), .B2(new_n613_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n799_), .A2(new_n800_), .A3(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n625_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT56), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n803_), .A2(KEYINPUT56), .A3(new_n625_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n798_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n542_), .B1(new_n797_), .B2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT119), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT57), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n809_), .A2(KEYINPUT119), .ZN(new_n813_));
  OAI21_X1  g612(.A(KEYINPUT120), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n808_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n541_), .B1(new_n815_), .B2(new_n796_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT57), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n806_), .A2(new_n807_), .ZN(new_n818_));
  AND3_X1   g617(.A1(new_n623_), .A2(new_n791_), .A3(new_n795_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n652_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT122), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n818_), .A2(KEYINPUT58), .A3(new_n819_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n822_), .A2(KEYINPUT122), .A3(new_n652_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n825_), .A2(new_n826_), .A3(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT119), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n816_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT120), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n830_), .A2(new_n831_), .A3(new_n811_), .A4(new_n810_), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n814_), .A2(new_n817_), .A3(new_n828_), .A4(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n790_), .B1(new_n833_), .B2(new_n580_), .ZN(new_n834_));
  NOR3_X1   g633(.A1(new_n287_), .A2(new_n444_), .A3(new_n480_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n634_), .ZN(new_n836_));
  NOR3_X1   g635(.A1(new_n834_), .A2(new_n604_), .A3(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(KEYINPUT123), .B1(new_n837_), .B2(G113gat), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT123), .ZN(new_n839_));
  OR2_X1    g638(.A1(new_n834_), .A2(new_n836_), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n839_), .B(new_n268_), .C1(new_n840_), .C2(new_n604_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n830_), .A2(new_n811_), .A3(new_n810_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n828_), .A2(new_n842_), .A3(new_n817_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n580_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n790_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n836_), .A2(KEYINPUT59), .ZN(new_n847_));
  AOI22_X1  g646(.A1(new_n840_), .A2(KEYINPUT59), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n604_), .A2(new_n268_), .ZN(new_n849_));
  AOI22_X1  g648(.A1(new_n838_), .A2(new_n841_), .B1(new_n848_), .B2(new_n849_), .ZN(G1340gat));
  NAND2_X1  g649(.A1(new_n846_), .A2(new_n847_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n834_), .A2(new_n836_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT59), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n851_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(G120gat), .B1(new_n854_), .B2(new_n631_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n266_), .B1(new_n631_), .B2(KEYINPUT60), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n852_), .B(new_n856_), .C1(KEYINPUT60), .C2(new_n266_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n857_), .ZN(G1341gat));
  OAI21_X1  g657(.A(G127gat), .B1(new_n854_), .B2(new_n580_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n852_), .A2(new_n264_), .A3(new_n579_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(G1342gat));
  INV_X1    g660(.A(new_n652_), .ZN(new_n862_));
  OAI21_X1  g661(.A(G134gat), .B1(new_n854_), .B2(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n852_), .A2(new_n262_), .A3(new_n541_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(G1343gat));
  NAND2_X1  g664(.A1(new_n833_), .A2(new_n580_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n845_), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n478_), .A2(new_n479_), .A3(new_n441_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n869_), .A2(new_n604_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(new_n300_), .ZN(G1344gat));
  NOR2_X1   g670(.A1(new_n869_), .A2(new_n631_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(new_n301_), .ZN(G1345gat));
  NOR2_X1   g672(.A1(new_n869_), .A2(new_n580_), .ZN(new_n874_));
  XOR2_X1   g673(.A(KEYINPUT61), .B(G155gat), .Z(new_n875_));
  XNOR2_X1  g674(.A(new_n874_), .B(new_n875_), .ZN(G1346gat));
  OAI21_X1  g675(.A(G162gat), .B1(new_n869_), .B2(new_n862_), .ZN(new_n877_));
  OR2_X1    g676(.A1(new_n542_), .A2(G162gat), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n869_), .B2(new_n878_), .ZN(G1347gat));
  INV_X1    g678(.A(KEYINPUT62), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n790_), .B1(new_n843_), .B2(new_n580_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n634_), .A2(new_n287_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(new_n480_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n883_), .A2(new_n444_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n881_), .A2(new_n604_), .A3(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT124), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(G169gat), .B1(new_n886_), .B2(new_n887_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n880_), .B1(new_n889_), .B2(new_n890_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n886_), .A2(new_n377_), .A3(new_n379_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n846_), .A2(new_n884_), .ZN(new_n893_));
  OAI21_X1  g692(.A(KEYINPUT124), .B1(new_n893_), .B2(new_n604_), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n894_), .A2(KEYINPUT62), .A3(new_n888_), .A4(G169gat), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n891_), .A2(new_n892_), .A3(new_n895_), .ZN(G1348gat));
  INV_X1    g695(.A(new_n444_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n867_), .A2(KEYINPUT126), .A3(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n883_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT126), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n900_), .B1(new_n834_), .B2(new_n444_), .ZN(new_n901_));
  AND3_X1   g700(.A1(new_n898_), .A2(new_n899_), .A3(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n631_), .A2(new_n207_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n207_), .B1(new_n893_), .B2(new_n631_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT125), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  OAI211_X1 g705(.A(KEYINPUT125), .B(new_n207_), .C1(new_n893_), .C2(new_n631_), .ZN(new_n907_));
  AOI22_X1  g706(.A1(new_n902_), .A2(new_n903_), .B1(new_n906_), .B2(new_n907_), .ZN(G1349gat));
  AOI211_X1 g707(.A(new_n580_), .B(new_n893_), .C1(new_n224_), .C2(new_n226_), .ZN(new_n909_));
  NAND4_X1  g708(.A1(new_n898_), .A2(new_n901_), .A3(new_n579_), .A4(new_n899_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n909_), .B1(new_n910_), .B2(new_n220_), .ZN(G1350gat));
  OAI21_X1  g710(.A(G190gat), .B1(new_n893_), .B2(new_n862_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n541_), .A2(new_n227_), .A3(new_n229_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n893_), .B2(new_n913_), .ZN(G1351gat));
  AND4_X1   g713(.A1(new_n479_), .A2(new_n287_), .A3(new_n444_), .A4(new_n480_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n867_), .A2(new_n915_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n916_), .A2(new_n604_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(new_n353_), .ZN(G1352gat));
  NOR2_X1   g717(.A1(new_n916_), .A2(new_n631_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n919_), .B(new_n920_), .ZN(G1353gat));
  NOR2_X1   g720(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n922_));
  AND2_X1   g721(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n923_));
  NOR4_X1   g722(.A1(new_n916_), .A2(new_n580_), .A3(new_n922_), .A4(new_n923_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n916_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(new_n579_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n924_), .B1(new_n926_), .B2(new_n922_), .ZN(G1354gat));
  OR3_X1    g726(.A1(new_n916_), .A2(G218gat), .A3(new_n542_), .ZN(new_n928_));
  OAI21_X1  g727(.A(G218gat), .B1(new_n916_), .B2(new_n862_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(G1355gat));
endmodule


