//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 1 0 1 1 0 1 0 0 1 0 1 1 0 0 1 0 1 1 1 1 0 1 0 0 1 0 0 0 0 1 0 0 1 1 1 0 0 1 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n614_, new_n615_, new_n616_, new_n617_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n685_, new_n686_, new_n687_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n711_, new_n712_, new_n713_, new_n715_, new_n716_,
    new_n717_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n812_, new_n813_,
    new_n814_, new_n816_, new_n817_, new_n818_, new_n820_, new_n821_,
    new_n822_, new_n824_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n855_, new_n856_, new_n858_,
    new_n859_, new_n861_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n879_, new_n880_;
  XOR2_X1   g000(.A(G85gat), .B(G92gat), .Z(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT9), .ZN(new_n203_));
  INV_X1    g002(.A(G85gat), .ZN(new_n204_));
  INV_X1    g003(.A(G92gat), .ZN(new_n205_));
  OR3_X1    g004(.A1(new_n204_), .A2(new_n205_), .A3(KEYINPUT9), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT6), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n203_), .A2(new_n206_), .A3(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT10), .B(G99gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT64), .ZN(new_n211_));
  INV_X1    g010(.A(G106gat), .ZN(new_n212_));
  AOI21_X1  g011(.A(KEYINPUT65), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n211_), .A2(KEYINPUT65), .A3(new_n212_), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n209_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT8), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT6), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n207_), .B(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT66), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT66), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n208_), .A2(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(G99gat), .A2(G106gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n223_), .B(KEYINPUT7), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n220_), .A2(new_n222_), .A3(new_n224_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n217_), .B1(new_n225_), .B2(new_n202_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(new_n208_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n227_), .A2(new_n217_), .A3(new_n202_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n226_), .A2(new_n229_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n216_), .A2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G57gat), .B(G64gat), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n232_), .A2(KEYINPUT11), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(KEYINPUT11), .ZN(new_n234_));
  XOR2_X1   g033(.A(G71gat), .B(G78gat), .Z(new_n235_));
  NAND3_X1  g034(.A1(new_n233_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  OR2_X1    g035(.A1(new_n234_), .A2(new_n235_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n231_), .A2(new_n238_), .ZN(new_n239_));
  OAI211_X1 g038(.A(new_n237_), .B(new_n236_), .C1(new_n216_), .C2(new_n230_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(KEYINPUT12), .A3(new_n240_), .ZN(new_n241_));
  OR3_X1    g040(.A1(new_n231_), .A2(KEYINPUT12), .A3(new_n238_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G230gat), .A2(G233gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT67), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n240_), .A2(new_n246_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n247_), .A2(new_n244_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n239_), .A2(new_n246_), .A3(new_n240_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n245_), .A2(new_n250_), .ZN(new_n251_));
  XOR2_X1   g050(.A(G120gat), .B(G148gat), .Z(new_n252_));
  XNOR2_X1  g051(.A(G176gat), .B(G204gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n252_), .B(new_n253_), .ZN(new_n254_));
  XOR2_X1   g053(.A(KEYINPUT68), .B(KEYINPUT5), .Z(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n251_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n256_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n245_), .A2(new_n250_), .A3(new_n258_), .ZN(new_n259_));
  AND2_X1   g058(.A1(new_n259_), .A2(KEYINPUT69), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n259_), .A2(KEYINPUT69), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n257_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT13), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n259_), .B(KEYINPUT69), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n265_), .A2(KEYINPUT13), .A3(new_n257_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G190gat), .B(G218gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G134gat), .B(G162gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n270_), .A2(KEYINPUT36), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G232gat), .A2(G233gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT34), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT35), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n230_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n209_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n215_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n279_), .B1(new_n280_), .B2(new_n213_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G29gat), .B(G36gat), .ZN(new_n282_));
  AND2_X1   g081(.A1(new_n282_), .A2(KEYINPUT70), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n282_), .A2(KEYINPUT70), .ZN(new_n284_));
  XOR2_X1   g083(.A(G43gat), .B(G50gat), .Z(new_n285_));
  OR3_X1    g084(.A1(new_n283_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n285_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n278_), .A2(new_n281_), .A3(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n275_), .A2(new_n276_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n289_), .A2(KEYINPUT15), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT15), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n288_), .A2(new_n294_), .ZN(new_n295_));
  AOI22_X1  g094(.A1(new_n278_), .A2(new_n281_), .B1(new_n293_), .B2(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n277_), .B1(new_n292_), .B2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n293_), .A2(new_n295_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n298_), .B1(new_n216_), .B2(new_n230_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n277_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n299_), .A2(new_n300_), .A3(new_n290_), .A4(new_n291_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n297_), .A2(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n272_), .B1(new_n302_), .B2(KEYINPUT71), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT71), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n297_), .A2(new_n301_), .A3(new_n304_), .A4(new_n271_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n302_), .A2(KEYINPUT36), .A3(new_n270_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(KEYINPUT72), .A2(KEYINPUT37), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n306_), .A2(new_n307_), .A3(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(KEYINPUT72), .A2(KEYINPUT37), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n311_), .B(KEYINPUT73), .Z(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n310_), .A2(new_n313_), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n306_), .A2(new_n307_), .A3(new_n309_), .A4(new_n312_), .ZN(new_n315_));
  AND2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  XOR2_X1   g115(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT75), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G127gat), .B(G155gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  XOR2_X1   g119(.A(G183gat), .B(G211gat), .Z(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT17), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G15gat), .B(G22gat), .ZN(new_n324_));
  INV_X1    g123(.A(G1gat), .ZN(new_n325_));
  INV_X1    g124(.A(G8gat), .ZN(new_n326_));
  OAI21_X1  g125(.A(KEYINPUT14), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n324_), .A2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G1gat), .B(G8gat), .ZN(new_n329_));
  XOR2_X1   g128(.A(new_n328_), .B(new_n329_), .Z(new_n330_));
  NAND2_X1  g129(.A1(G231gat), .A2(G233gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(new_n238_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n323_), .B1(KEYINPUT77), .B2(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n334_), .B1(KEYINPUT77), .B2(new_n333_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n322_), .A2(KEYINPUT17), .ZN(new_n336_));
  XOR2_X1   g135(.A(new_n336_), .B(KEYINPUT76), .Z(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(new_n333_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n335_), .A2(new_n338_), .ZN(new_n339_));
  NOR3_X1   g138(.A1(new_n267_), .A2(new_n316_), .A3(new_n339_), .ZN(new_n340_));
  OR2_X1    g139(.A1(KEYINPUT78), .A2(G183gat), .ZN(new_n341_));
  INV_X1    g140(.A(G190gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(KEYINPUT78), .A2(G183gat), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n341_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G183gat), .A2(G190gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT23), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT23), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n347_), .A2(G183gat), .A3(G190gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(KEYINPUT81), .B1(new_n344_), .B2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT22), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n351_), .A2(KEYINPUT80), .A3(G169gat), .ZN(new_n352_));
  INV_X1    g151(.A(G176gat), .ZN(new_n353_));
  AND2_X1   g152(.A1(KEYINPUT80), .A2(G169gat), .ZN(new_n354_));
  OAI211_X1 g153(.A(new_n352_), .B(new_n353_), .C1(new_n351_), .C2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G169gat), .A2(G176gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n350_), .A2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n344_), .A2(new_n349_), .A3(KEYINPUT81), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n356_), .A2(KEYINPUT24), .ZN(new_n360_));
  NOR2_X1   g159(.A1(G169gat), .A2(G176gat), .ZN(new_n361_));
  OR2_X1    g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT24), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n361_), .A2(new_n363_), .ZN(new_n364_));
  AND3_X1   g163(.A1(new_n362_), .A2(new_n349_), .A3(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT79), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(G190gat), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT26), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT25), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n371_), .B1(new_n341_), .B2(new_n343_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n369_), .B1(new_n370_), .B2(new_n372_), .ZN(new_n373_));
  AOI22_X1  g172(.A1(new_n358_), .A2(new_n359_), .B1(new_n365_), .B2(new_n373_), .ZN(new_n374_));
  XOR2_X1   g173(.A(G71gat), .B(G99gat), .Z(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(G43gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n374_), .B(new_n376_), .ZN(new_n377_));
  XOR2_X1   g176(.A(G127gat), .B(G134gat), .Z(new_n378_));
  XOR2_X1   g177(.A(G113gat), .B(G120gat), .Z(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n377_), .B(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G227gat), .A2(G233gat), .ZN(new_n383_));
  INV_X1    g182(.A(G15gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(KEYINPUT30), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT31), .ZN(new_n387_));
  AND2_X1   g186(.A1(new_n382_), .A2(new_n387_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n382_), .A2(new_n387_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT87), .ZN(new_n391_));
  NOR2_X1   g190(.A1(G197gat), .A2(G204gat), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT84), .B(G197gat), .ZN(new_n394_));
  INV_X1    g193(.A(G204gat), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n393_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT21), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G211gat), .B(G218gat), .ZN(new_n398_));
  NOR3_X1   g197(.A1(new_n396_), .A2(new_n397_), .A3(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT85), .ZN(new_n400_));
  INV_X1    g199(.A(G197gat), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n400_), .B1(new_n401_), .B2(G204gat), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n402_), .B1(new_n394_), .B2(G204gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(KEYINPUT84), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT84), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(G197gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n404_), .A2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n407_), .A2(new_n400_), .A3(new_n395_), .ZN(new_n408_));
  AND3_X1   g207(.A1(new_n403_), .A2(new_n408_), .A3(KEYINPUT21), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n392_), .B1(new_n407_), .B2(G204gat), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n398_), .B1(new_n410_), .B2(KEYINPUT21), .ZN(new_n411_));
  OAI21_X1  g210(.A(KEYINPUT86), .B1(new_n409_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n398_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n413_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT86), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n403_), .A2(new_n408_), .A3(KEYINPUT21), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n414_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n399_), .B1(new_n412_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G228gat), .A2(G233gat), .ZN(new_n419_));
  AOI21_X1  g218(.A(KEYINPUT82), .B1(G155gat), .B2(G162gat), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT1), .ZN(new_n422_));
  NAND3_X1  g221(.A1(KEYINPUT82), .A2(G155gat), .A3(G162gat), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n421_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n423_), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT1), .B1(new_n425_), .B2(new_n420_), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n424_), .B(new_n426_), .C1(G155gat), .C2(G162gat), .ZN(new_n427_));
  INV_X1    g226(.A(G141gat), .ZN(new_n428_));
  INV_X1    g227(.A(G148gat), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(G141gat), .A2(G148gat), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT83), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT2), .B1(new_n430_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT2), .ZN(new_n435_));
  OAI211_X1 g234(.A(KEYINPUT83), .B(new_n435_), .C1(new_n428_), .C2(new_n429_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT3), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n431_), .A2(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n434_), .A2(new_n436_), .A3(new_n438_), .A4(new_n439_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(G155gat), .A2(G162gat), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n441_), .B1(new_n421_), .B2(new_n423_), .ZN(new_n442_));
  AOI22_X1  g241(.A1(new_n427_), .A2(new_n432_), .B1(new_n440_), .B2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT29), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n419_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n391_), .B1(new_n418_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n399_), .ZN(new_n447_));
  AND3_X1   g246(.A1(new_n414_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n415_), .B1(new_n414_), .B2(new_n416_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n447_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n427_), .A2(new_n432_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n440_), .A2(new_n442_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT29), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n450_), .A2(KEYINPUT87), .A3(new_n419_), .A4(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n446_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n454_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n450_), .A2(KEYINPUT88), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT88), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n459_), .B(new_n447_), .C1(new_n448_), .C2(new_n449_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n457_), .B1(new_n458_), .B2(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n456_), .B1(new_n461_), .B2(new_n419_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G78gat), .B(G106gat), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G22gat), .B(G50gat), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n443_), .A2(new_n444_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(KEYINPUT28), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n468_), .A2(KEYINPUT28), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n467_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n471_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n473_), .A2(new_n469_), .A3(new_n466_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  OAI211_X1 g274(.A(new_n456_), .B(new_n463_), .C1(new_n461_), .C2(new_n419_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n465_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n464_), .A2(KEYINPUT89), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n462_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n475_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n478_), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n456_), .B(new_n481_), .C1(new_n461_), .C2(new_n419_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n479_), .A2(new_n480_), .A3(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT90), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n477_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n475_), .B1(new_n462_), .B2(new_n478_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n486_), .A2(KEYINPUT90), .A3(new_n482_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n485_), .A2(new_n487_), .ZN(new_n488_));
  XOR2_X1   g287(.A(G1gat), .B(G29gat), .Z(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT94), .B(G85gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(KEYINPUT0), .B(G57gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n453_), .A2(new_n381_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n443_), .A2(new_n380_), .ZN(new_n495_));
  AND2_X1   g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G225gat), .A2(G233gat), .ZN(new_n497_));
  XOR2_X1   g296(.A(new_n497_), .B(KEYINPUT93), .Z(new_n498_));
  NOR2_X1   g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n498_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n494_), .A2(KEYINPUT4), .A3(new_n495_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT4), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n453_), .A2(new_n502_), .A3(new_n381_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n500_), .B1(new_n501_), .B2(new_n503_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n493_), .B1(new_n499_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT33), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  OAI211_X1 g306(.A(KEYINPUT33), .B(new_n493_), .C1(new_n499_), .C2(new_n504_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n493_), .B1(new_n496_), .B2(new_n498_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n501_), .A2(new_n500_), .A3(new_n503_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  AND3_X1   g310(.A1(new_n507_), .A2(new_n508_), .A3(new_n511_), .ZN(new_n512_));
  OAI211_X1 g311(.A(new_n374_), .B(new_n447_), .C1(new_n448_), .C2(new_n449_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n349_), .B1(G183gat), .B2(G190gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(KEYINPUT22), .B(G169gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(new_n353_), .ZN(new_n516_));
  AND3_X1   g315(.A1(new_n514_), .A2(new_n356_), .A3(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(KEYINPUT25), .B(G183gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(KEYINPUT26), .B(G190gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n520_), .A2(new_n362_), .A3(new_n349_), .A4(new_n364_), .ZN(new_n521_));
  OR2_X1    g320(.A1(new_n521_), .A2(KEYINPUT91), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(KEYINPUT91), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n517_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  OAI211_X1 g323(.A(new_n513_), .B(KEYINPUT20), .C1(new_n418_), .C2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G226gat), .A2(G233gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT19), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n525_), .A2(new_n527_), .ZN(new_n528_));
  XOR2_X1   g327(.A(G8gat), .B(G36gat), .Z(new_n529_));
  XNOR2_X1  g328(.A(G64gat), .B(G92gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT20), .ZN(new_n535_));
  INV_X1    g334(.A(new_n374_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n535_), .B1(new_n450_), .B2(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n527_), .B1(new_n418_), .B2(new_n524_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  AND3_X1   g338(.A1(new_n528_), .A2(new_n534_), .A3(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n534_), .B1(new_n528_), .B2(new_n539_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  OR3_X1    g341(.A1(new_n499_), .A2(new_n504_), .A3(new_n493_), .ZN(new_n543_));
  AOI22_X1  g342(.A1(new_n525_), .A2(new_n527_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n534_), .A2(KEYINPUT32), .ZN(new_n545_));
  AOI22_X1  g344(.A1(new_n543_), .A2(new_n505_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n527_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n521_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n517_), .A2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n458_), .A2(new_n460_), .A3(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n547_), .B1(new_n550_), .B2(new_n537_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n525_), .A2(new_n527_), .ZN(new_n552_));
  OAI211_X1 g351(.A(KEYINPUT32), .B(new_n534_), .C1(new_n551_), .C2(new_n552_), .ZN(new_n553_));
  AOI22_X1  g352(.A1(new_n512_), .A2(new_n542_), .B1(new_n546_), .B2(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n390_), .B1(new_n488_), .B2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT27), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n556_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n543_), .A2(new_n505_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n533_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n556_), .B1(new_n544_), .B2(new_n534_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n557_), .A2(new_n559_), .A3(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n563_), .A2(new_n485_), .A3(new_n487_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n557_), .A2(new_n562_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n565_), .B1(new_n485_), .B2(new_n487_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n390_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n567_), .A2(new_n558_), .ZN(new_n568_));
  AOI22_X1  g367(.A1(new_n555_), .A2(new_n564_), .B1(new_n566_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n330_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(new_n288_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G229gat), .A2(G233gat), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n571_), .A2(new_n573_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n570_), .A2(new_n288_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n575_), .B1(new_n298_), .B2(new_n570_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n574_), .B1(new_n572_), .B2(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(G113gat), .B(G141gat), .Z(new_n578_));
  XNOR2_X1  g377(.A(G169gat), .B(G197gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n577_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n577_), .A2(new_n580_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n569_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n340_), .A2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT95), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n558_), .B(KEYINPUT96), .Z(new_n588_));
  NAND3_X1  g387(.A1(new_n587_), .A2(new_n325_), .A3(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT38), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n306_), .A2(new_n307_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n569_), .A2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT97), .ZN(new_n594_));
  NOR3_X1   g393(.A1(new_n267_), .A2(new_n584_), .A3(new_n339_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  OAI21_X1  g395(.A(G1gat), .B1(new_n596_), .B2(new_n559_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n589_), .A2(new_n590_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n591_), .A2(new_n597_), .A3(new_n598_), .ZN(G1324gat));
  NAND3_X1  g398(.A1(new_n587_), .A2(new_n326_), .A3(new_n565_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT98), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n565_), .ZN(new_n603_));
  OAI21_X1  g402(.A(G8gat), .B1(new_n596_), .B2(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT39), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n602_), .A2(new_n605_), .ZN(new_n606_));
  XOR2_X1   g405(.A(new_n606_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g406(.A(G15gat), .B1(new_n596_), .B2(new_n567_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(KEYINPUT99), .B(KEYINPUT41), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n609_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n390_), .A2(new_n384_), .ZN(new_n612_));
  OAI211_X1 g411(.A(new_n610_), .B(new_n611_), .C1(new_n586_), .C2(new_n612_), .ZN(G1326gat));
  OAI21_X1  g412(.A(G22gat), .B1(new_n596_), .B2(new_n488_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT42), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n488_), .A2(G22gat), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n616_), .B(KEYINPUT100), .Z(new_n617_));
  OAI21_X1  g416(.A(new_n615_), .B1(new_n586_), .B2(new_n617_), .ZN(G1327gat));
  INV_X1    g417(.A(G29gat), .ZN(new_n619_));
  XOR2_X1   g418(.A(KEYINPUT102), .B(KEYINPUT44), .Z(new_n620_));
  INV_X1    g419(.A(KEYINPUT101), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n314_), .A2(new_n315_), .ZN(new_n622_));
  OAI21_X1  g421(.A(KEYINPUT43), .B1(new_n569_), .B2(new_n622_), .ZN(new_n623_));
  AND4_X1   g422(.A1(KEYINPUT90), .A2(new_n479_), .A3(new_n480_), .A4(new_n482_), .ZN(new_n624_));
  AOI21_X1  g423(.A(KEYINPUT90), .B1(new_n486_), .B2(new_n482_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n624_), .B1(new_n477_), .B2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n512_), .A2(new_n542_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n546_), .A2(new_n553_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  OAI211_X1 g428(.A(new_n564_), .B(new_n567_), .C1(new_n626_), .C2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n566_), .A2(new_n568_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT43), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n632_), .A2(new_n316_), .A3(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n623_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n584_), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n264_), .A2(new_n266_), .A3(new_n636_), .A4(new_n339_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n621_), .B1(new_n635_), .B2(new_n638_), .ZN(new_n639_));
  AOI211_X1 g438(.A(KEYINPUT101), .B(new_n637_), .C1(new_n623_), .C2(new_n634_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n620_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n637_), .B1(new_n623_), .B2(new_n634_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(KEYINPUT44), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n641_), .A2(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n619_), .B1(new_n644_), .B2(new_n588_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT103), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n592_), .A2(new_n339_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n267_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(new_n585_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n558_), .A2(new_n619_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n646_), .B1(new_n649_), .B2(new_n650_), .ZN(G1328gat));
  INV_X1    g450(.A(KEYINPUT104), .ZN(new_n652_));
  INV_X1    g451(.A(new_n620_), .ZN(new_n653_));
  NOR3_X1   g452(.A1(new_n569_), .A2(KEYINPUT43), .A3(new_n622_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n633_), .B1(new_n632_), .B2(new_n316_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n638_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(KEYINPUT101), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n642_), .A2(new_n621_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n653_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n603_), .B1(new_n642_), .B2(KEYINPUT44), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(G36gat), .B1(new_n659_), .B2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(G36gat), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n648_), .A2(new_n585_), .A3(new_n663_), .A4(new_n565_), .ZN(new_n664_));
  XOR2_X1   g463(.A(new_n664_), .B(KEYINPUT45), .Z(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n662_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT46), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n652_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  AOI211_X1 g468(.A(KEYINPUT104), .B(KEYINPUT46), .C1(new_n662_), .C2(new_n666_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n641_), .A2(new_n660_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n665_), .B1(new_n671_), .B2(G36gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(KEYINPUT105), .B1(new_n672_), .B2(KEYINPUT46), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n663_), .B1(new_n641_), .B2(new_n660_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT105), .ZN(new_n675_));
  NOR4_X1   g474(.A1(new_n674_), .A2(new_n675_), .A3(new_n668_), .A4(new_n665_), .ZN(new_n676_));
  OAI22_X1  g475(.A1(new_n669_), .A2(new_n670_), .B1(new_n673_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT106), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  OAI21_X1  g478(.A(KEYINPUT104), .B1(new_n672_), .B2(KEYINPUT46), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n667_), .A2(new_n652_), .A3(new_n668_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  OAI211_X1 g481(.A(new_n682_), .B(KEYINPUT106), .C1(new_n673_), .C2(new_n676_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n679_), .A2(new_n683_), .ZN(G1329gat));
  NOR3_X1   g483(.A1(new_n649_), .A2(G43gat), .A3(new_n567_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n644_), .A2(new_n390_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n685_), .B1(new_n686_), .B2(G43gat), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g487(.A1(new_n649_), .A2(G50gat), .A3(new_n488_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n644_), .A2(KEYINPUT107), .A3(new_n626_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(G50gat), .ZN(new_n691_));
  AOI21_X1  g490(.A(KEYINPUT107), .B1(new_n644_), .B2(new_n626_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n689_), .B1(new_n691_), .B2(new_n692_), .ZN(G1331gat));
  INV_X1    g492(.A(new_n339_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n267_), .A2(new_n694_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n695_), .A2(new_n636_), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n594_), .A2(G57gat), .A3(new_n558_), .A4(new_n696_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n697_), .A2(KEYINPUT108), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n697_), .A2(KEYINPUT108), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n695_), .A2(new_n316_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n569_), .A2(new_n636_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(G57gat), .B1(new_n703_), .B2(new_n588_), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n698_), .A2(new_n699_), .A3(new_n704_), .ZN(G1332gat));
  NAND2_X1  g504(.A1(new_n594_), .A2(new_n696_), .ZN(new_n706_));
  OAI21_X1  g505(.A(G64gat), .B1(new_n706_), .B2(new_n603_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT48), .ZN(new_n708_));
  OR2_X1    g507(.A1(new_n603_), .A2(G64gat), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n708_), .B1(new_n702_), .B2(new_n709_), .ZN(G1333gat));
  OAI21_X1  g509(.A(G71gat), .B1(new_n706_), .B2(new_n567_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT49), .ZN(new_n712_));
  OR2_X1    g511(.A1(new_n567_), .A2(G71gat), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n712_), .B1(new_n702_), .B2(new_n713_), .ZN(G1334gat));
  OAI21_X1  g513(.A(G78gat), .B1(new_n706_), .B2(new_n488_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT50), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n488_), .A2(G78gat), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n716_), .B1(new_n702_), .B2(new_n717_), .ZN(G1335gat));
  NAND4_X1  g517(.A1(new_n635_), .A2(new_n584_), .A3(new_n267_), .A4(new_n339_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n719_), .A2(KEYINPUT110), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n719_), .A2(KEYINPUT110), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  NOR3_X1   g521(.A1(new_n722_), .A2(new_n204_), .A3(new_n559_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n267_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n724_), .A2(new_n647_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(new_n701_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n588_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n204_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT109), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n723_), .A2(new_n729_), .ZN(G1336gat));
  OAI21_X1  g529(.A(G92gat), .B1(new_n722_), .B2(new_n603_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n726_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n732_), .A2(new_n205_), .A3(new_n565_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT111), .Z(G1337gat));
  AND3_X1   g534(.A1(new_n732_), .A2(new_n390_), .A3(new_n211_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n390_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n737_), .B2(G99gat), .ZN(new_n738_));
  XNOR2_X1  g537(.A(KEYINPUT112), .B(KEYINPUT51), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n738_), .B(new_n739_), .Z(G1338gat));
  OAI21_X1  g539(.A(G106gat), .B1(new_n719_), .B2(new_n488_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT52), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n732_), .A2(new_n212_), .A3(new_n626_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n744_), .B(new_n745_), .Z(G1339gat));
  NAND2_X1  g545(.A1(new_n340_), .A2(new_n584_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(KEYINPUT114), .A2(KEYINPUT54), .ZN(new_n748_));
  AND2_X1   g547(.A1(KEYINPUT114), .A2(KEYINPUT54), .ZN(new_n749_));
  OR3_X1    g548(.A1(new_n747_), .A2(new_n748_), .A3(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n747_), .A2(new_n748_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n244_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT55), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n258_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n245_), .A2(KEYINPUT55), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n243_), .A2(new_n244_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n756_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT56), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  OR2_X1    g560(.A1(new_n761_), .A2(KEYINPUT116), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(KEYINPUT116), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n759_), .A2(new_n760_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n762_), .A2(new_n763_), .A3(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT115), .ZN(new_n766_));
  OR2_X1    g565(.A1(new_n576_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n576_), .A2(new_n766_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n767_), .A2(new_n573_), .A3(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n580_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n582_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n265_), .A2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n765_), .A2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT58), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n622_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n775_), .B1(new_n774_), .B2(new_n773_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n262_), .A2(new_n771_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n759_), .B(KEYINPUT56), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n265_), .A2(new_n636_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n777_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n592_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT57), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n694_), .B1(new_n776_), .B2(new_n783_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n752_), .A2(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n566_), .A2(new_n390_), .A3(new_n588_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n636_), .ZN(new_n788_));
  INV_X1    g587(.A(G113gat), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n788_), .A2(KEYINPUT117), .A3(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n636_), .A2(G113gat), .ZN(new_n791_));
  NAND2_X1  g590(.A1(KEYINPUT118), .A2(KEYINPUT59), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT118), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT59), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n787_), .A2(new_n792_), .A3(new_n795_), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n793_), .B(new_n794_), .C1(new_n785_), .C2(new_n786_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n791_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(KEYINPUT117), .B1(new_n788_), .B2(new_n789_), .ZN(new_n799_));
  NOR3_X1   g598(.A1(new_n790_), .A2(new_n798_), .A3(new_n799_), .ZN(G1340gat));
  AND2_X1   g599(.A1(new_n776_), .A2(new_n783_), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n751_), .B(new_n750_), .C1(new_n801_), .C2(new_n694_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n786_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT60), .ZN(new_n804_));
  AOI21_X1  g603(.A(G120gat), .B1(new_n267_), .B2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n805_), .B1(new_n804_), .B2(G120gat), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n802_), .A2(new_n803_), .A3(new_n806_), .ZN(new_n807_));
  XOR2_X1   g606(.A(new_n807_), .B(KEYINPUT119), .Z(new_n808_));
  INV_X1    g607(.A(G120gat), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n724_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n808_), .B1(new_n809_), .B2(new_n810_), .ZN(G1341gat));
  INV_X1    g610(.A(G127gat), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n787_), .A2(new_n812_), .A3(new_n694_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n339_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n813_), .B1(new_n814_), .B2(new_n812_), .ZN(G1342gat));
  INV_X1    g614(.A(G134gat), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n787_), .A2(new_n816_), .A3(new_n592_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n622_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n817_), .B1(new_n818_), .B2(new_n816_), .ZN(G1343gat));
  NOR3_X1   g618(.A1(new_n727_), .A2(new_n390_), .A3(new_n565_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n802_), .A2(new_n626_), .A3(new_n820_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n821_), .A2(new_n584_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n822_), .B(new_n428_), .ZN(G1344gat));
  NOR2_X1   g622(.A1(new_n821_), .A2(new_n724_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n824_), .B(new_n429_), .ZN(G1345gat));
  OAI21_X1  g624(.A(KEYINPUT120), .B1(new_n821_), .B2(new_n339_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n785_), .A2(new_n488_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT120), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n827_), .A2(new_n828_), .A3(new_n694_), .A4(new_n820_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(KEYINPUT61), .B(G155gat), .ZN(new_n830_));
  AND3_X1   g629(.A1(new_n826_), .A2(new_n829_), .A3(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n830_), .B1(new_n826_), .B2(new_n829_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n831_), .A2(new_n832_), .ZN(G1346gat));
  INV_X1    g632(.A(new_n821_), .ZN(new_n834_));
  AOI21_X1  g633(.A(G162gat), .B1(new_n834_), .B2(new_n592_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n316_), .A2(G162gat), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n836_), .B(KEYINPUT121), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n835_), .B1(new_n834_), .B2(new_n837_), .ZN(G1347gat));
  NOR4_X1   g637(.A1(new_n626_), .A2(new_n588_), .A3(new_n603_), .A4(new_n567_), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n636_), .B(new_n839_), .C1(new_n752_), .C2(new_n784_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT62), .ZN(new_n841_));
  AND3_X1   g640(.A1(new_n840_), .A2(new_n841_), .A3(G169gat), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n841_), .B1(new_n840_), .B2(G169gat), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n802_), .A2(new_n839_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n636_), .A2(new_n515_), .ZN(new_n845_));
  XOR2_X1   g644(.A(new_n845_), .B(KEYINPUT122), .Z(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  OAI22_X1  g646(.A1(new_n842_), .A2(new_n843_), .B1(new_n844_), .B2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT123), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  OAI221_X1 g649(.A(KEYINPUT123), .B1(new_n844_), .B2(new_n847_), .C1(new_n842_), .C2(new_n843_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(G1348gat));
  NOR2_X1   g651(.A1(new_n844_), .A2(new_n724_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(new_n353_), .ZN(G1349gat));
  NAND2_X1  g653(.A1(new_n341_), .A2(new_n343_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n844_), .A2(new_n339_), .ZN(new_n856_));
  MUX2_X1   g655(.A(new_n855_), .B(new_n518_), .S(new_n856_), .Z(G1350gat));
  OAI21_X1  g656(.A(G190gat), .B1(new_n844_), .B2(new_n622_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n592_), .A2(new_n519_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n844_), .B2(new_n859_), .ZN(G1351gat));
  NOR3_X1   g659(.A1(new_n603_), .A2(new_n390_), .A3(new_n558_), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n626_), .B(new_n861_), .C1(new_n752_), .C2(new_n784_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n862_), .A2(new_n584_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(KEYINPUT124), .B(G197gat), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n863_), .B(new_n864_), .ZN(G1352gat));
  INV_X1    g664(.A(new_n862_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n267_), .ZN(new_n867_));
  AND2_X1   g666(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n868_));
  NOR2_X1   g667(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n867_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n870_), .B1(new_n867_), .B2(new_n868_), .ZN(G1353gat));
  XNOR2_X1  g670(.A(KEYINPUT63), .B(G211gat), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n866_), .A2(new_n694_), .A3(new_n872_), .ZN(new_n873_));
  OAI22_X1  g672(.A1(new_n862_), .A2(new_n339_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT126), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n875_), .B(new_n876_), .ZN(G1354gat));
  XNOR2_X1  g676(.A(KEYINPUT127), .B(G218gat), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n862_), .A2(new_n622_), .A3(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n866_), .A2(new_n592_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n879_), .B1(new_n880_), .B2(new_n878_), .ZN(G1355gat));
endmodule


