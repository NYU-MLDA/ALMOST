//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 0 1 1 0 0 0 1 1 1 1 0 1 1 1 1 1 1 0 1 0 1 1 0 0 1 0 0 0 1 1 0 0 0 0 1 0 1 1 1 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n790_,
    new_n791_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n825_, new_n826_,
    new_n828_, new_n829_, new_n830_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n928_, new_n929_, new_n930_,
    new_n931_, new_n933_, new_n934_, new_n935_, new_n936_, new_n938_,
    new_n939_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n953_, new_n954_, new_n956_, new_n957_, new_n959_, new_n960_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n967_, new_n968_,
    new_n969_, new_n970_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n977_, new_n978_;
  INV_X1    g000(.A(KEYINPUT37), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT70), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT64), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT10), .B(G99gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(new_n204_), .B1(new_n205_), .B2(G106gat), .ZN(new_n206_));
  OR2_X1    g005(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n207_));
  INV_X1    g006(.A(G106gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n209_));
  NAND4_X1  g008(.A1(new_n207_), .A2(KEYINPUT64), .A3(new_n208_), .A4(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n206_), .A2(new_n210_), .ZN(new_n211_));
  AND2_X1   g010(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n212_));
  NOR2_X1   g011(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n213_));
  INV_X1    g012(.A(G85gat), .ZN(new_n214_));
  INV_X1    g013(.A(G92gat), .ZN(new_n215_));
  OAI22_X1  g014(.A1(new_n212_), .A2(new_n213_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n217_));
  OR2_X1    g016(.A1(new_n217_), .A2(KEYINPUT66), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n214_), .A2(new_n215_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(KEYINPUT66), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n216_), .A2(new_n218_), .A3(new_n219_), .A4(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G99gat), .A2(G106gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT6), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT6), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n224_), .A2(G99gat), .A3(G106gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n223_), .A2(new_n225_), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n211_), .A2(KEYINPUT67), .A3(new_n221_), .A4(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT7), .ZN(new_n228_));
  INV_X1    g027(.A(G99gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n228_), .A2(new_n229_), .A3(new_n208_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT68), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n228_), .A2(new_n229_), .A3(new_n208_), .A4(KEYINPUT68), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n232_), .A2(new_n226_), .A3(new_n233_), .A4(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT8), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT69), .B1(new_n214_), .B2(new_n215_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n237_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n238_));
  AND3_X1   g037(.A1(new_n235_), .A2(new_n236_), .A3(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n236_), .B1(new_n235_), .B2(new_n238_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n227_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  AOI22_X1  g040(.A1(new_n206_), .A2(new_n210_), .B1(new_n223_), .B2(new_n225_), .ZN(new_n242_));
  AOI21_X1  g041(.A(KEYINPUT67), .B1(new_n242_), .B2(new_n221_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n203_), .B1(new_n241_), .B2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G29gat), .B(G36gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G43gat), .B(G50gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT15), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n235_), .A2(new_n238_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT8), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n235_), .A2(new_n236_), .A3(new_n238_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n211_), .A2(new_n221_), .A3(new_n226_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT67), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n252_), .A2(new_n255_), .A3(KEYINPUT70), .A4(new_n227_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n244_), .A2(new_n248_), .A3(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G232gat), .A2(G233gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT34), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n259_), .A2(KEYINPUT35), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n241_), .A2(new_n243_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n260_), .B1(new_n261_), .B2(new_n247_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n259_), .A2(KEYINPUT35), .ZN(new_n263_));
  AND3_X1   g062(.A1(new_n257_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n263_), .B1(new_n257_), .B2(new_n262_), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT74), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  XOR2_X1   g065(.A(G190gat), .B(G218gat), .Z(new_n267_));
  XNOR2_X1  g066(.A(G134gat), .B(G162gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  XOR2_X1   g068(.A(KEYINPUT72), .B(KEYINPUT73), .Z(new_n270_));
  XOR2_X1   g069(.A(new_n269_), .B(new_n270_), .Z(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(KEYINPUT36), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT36), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n257_), .A2(new_n262_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n263_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n257_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n274_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  OAI211_X1 g078(.A(new_n266_), .B(new_n273_), .C1(new_n279_), .C2(new_n272_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  OAI21_X1  g080(.A(KEYINPUT36), .B1(new_n264_), .B2(new_n265_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(new_n271_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n266_), .B1(new_n283_), .B2(new_n273_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n202_), .B1(new_n281_), .B2(new_n284_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n273_), .B1(new_n279_), .B2(new_n272_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n266_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n288_), .A2(KEYINPUT37), .A3(new_n280_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n285_), .A2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT75), .B(G1gat), .ZN(new_n291_));
  INV_X1    g090(.A(G8gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT14), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G15gat), .B(G22gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G1gat), .B(G8gat), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n295_), .A2(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n293_), .A2(new_n294_), .A3(new_n296_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G231gat), .A2(G233gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT76), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n300_), .B(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G57gat), .B(G64gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT11), .ZN(new_n305_));
  XOR2_X1   g104(.A(G71gat), .B(G78gat), .Z(new_n306_));
  NOR2_X1   g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  AND2_X1   g106(.A1(new_n305_), .A2(new_n306_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n304_), .A2(KEYINPUT11), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n307_), .B1(new_n308_), .B2(new_n310_), .ZN(new_n311_));
  AND2_X1   g110(.A1(new_n303_), .A2(new_n311_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n303_), .A2(new_n311_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n314_), .A2(KEYINPUT77), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(KEYINPUT77), .ZN(new_n316_));
  XOR2_X1   g115(.A(G127gat), .B(G155gat), .Z(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT16), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G183gat), .B(G211gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT17), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n315_), .A2(new_n316_), .A3(new_n322_), .ZN(new_n323_));
  OR2_X1    g122(.A1(new_n314_), .A2(KEYINPUT78), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n314_), .A2(KEYINPUT78), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n320_), .B(KEYINPUT17), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n324_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n323_), .A2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT79), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n290_), .A2(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n252_), .A2(new_n255_), .A3(new_n227_), .ZN(new_n331_));
  OAI21_X1  g130(.A(KEYINPUT12), .B1(new_n331_), .B2(new_n311_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n311_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G230gat), .A2(G233gat), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n244_), .A2(KEYINPUT12), .A3(new_n256_), .A4(new_n311_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n334_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  OR2_X1    g136(.A1(new_n331_), .A2(new_n311_), .ZN(new_n338_));
  AND2_X1   g137(.A1(new_n338_), .A2(new_n333_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n337_), .B1(new_n335_), .B2(new_n339_), .ZN(new_n340_));
  XOR2_X1   g139(.A(G120gat), .B(G148gat), .Z(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT5), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G176gat), .B(G204gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  XOR2_X1   g143(.A(new_n340_), .B(new_n344_), .Z(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT71), .B(KEYINPUT13), .ZN(new_n346_));
  OR2_X1    g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT13), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n345_), .B1(KEYINPUT71), .B2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n347_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n330_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n300_), .A2(new_n247_), .ZN(new_n352_));
  XOR2_X1   g151(.A(new_n352_), .B(KEYINPUT80), .Z(new_n353_));
  INV_X1    g152(.A(new_n300_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n247_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n353_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G229gat), .A2(G233gat), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n357_), .A2(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n352_), .B(KEYINPUT80), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n248_), .A2(new_n354_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(new_n358_), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT81), .B1(new_n361_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT81), .ZN(new_n365_));
  INV_X1    g164(.A(new_n363_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n353_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G113gat), .B(G141gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G169gat), .B(G197gat), .ZN(new_n369_));
  XOR2_X1   g168(.A(new_n368_), .B(new_n369_), .Z(new_n370_));
  NAND4_X1  g169(.A1(new_n360_), .A2(new_n364_), .A3(new_n367_), .A4(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(KEYINPUT83), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n361_), .A2(new_n363_), .ZN(new_n373_));
  AOI22_X1  g172(.A1(new_n357_), .A2(new_n359_), .B1(new_n373_), .B2(new_n365_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT83), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n374_), .A2(new_n375_), .A3(new_n364_), .A4(new_n370_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n372_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT82), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n361_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n367_), .B1(new_n379_), .B2(new_n358_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n364_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n378_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n370_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n374_), .A2(KEYINPUT82), .A3(new_n364_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n382_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n377_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT27), .ZN(new_n388_));
  XOR2_X1   g187(.A(G8gat), .B(G36gat), .Z(new_n389_));
  XNOR2_X1  g188(.A(G64gat), .B(G92gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT101), .B(KEYINPUT18), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT96), .ZN(new_n394_));
  NOR2_X1   g193(.A1(G197gat), .A2(G204gat), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G197gat), .A2(G204gat), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n396_), .A2(KEYINPUT21), .A3(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT21), .ZN(new_n399_));
  INV_X1    g198(.A(new_n397_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n399_), .B1(new_n400_), .B2(new_n395_), .ZN(new_n401_));
  INV_X1    g200(.A(G218gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(G211gat), .ZN(new_n403_));
  INV_X1    g202(.A(G211gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(G218gat), .ZN(new_n405_));
  AND3_X1   g204(.A1(new_n403_), .A2(new_n405_), .A3(KEYINPUT95), .ZN(new_n406_));
  AOI21_X1  g205(.A(KEYINPUT95), .B1(new_n403_), .B2(new_n405_), .ZN(new_n407_));
  OAI211_X1 g206(.A(new_n398_), .B(new_n401_), .C1(new_n406_), .C2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n403_), .A2(new_n405_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT95), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n403_), .A2(new_n405_), .A3(KEYINPUT95), .ZN(new_n412_));
  NOR3_X1   g211(.A1(new_n400_), .A2(new_n395_), .A3(new_n399_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n411_), .A2(new_n412_), .A3(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n394_), .B1(new_n408_), .B2(new_n414_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n398_), .A2(new_n401_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n411_), .A2(new_n412_), .ZN(new_n417_));
  AOI21_X1  g216(.A(KEYINPUT96), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n415_), .A2(new_n418_), .ZN(new_n419_));
  OR3_X1    g218(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G183gat), .A2(G190gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT23), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(KEYINPUT84), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT84), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n424_), .A2(G183gat), .A3(G190gat), .ZN(new_n425_));
  AOI21_X1  g224(.A(KEYINPUT23), .B1(new_n423_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT85), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n422_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  AOI211_X1 g227(.A(KEYINPUT85), .B(KEYINPUT23), .C1(new_n423_), .C2(new_n425_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n420_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT86), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  OAI211_X1 g231(.A(KEYINPUT86), .B(new_n420_), .C1(new_n428_), .C2(new_n429_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(KEYINPUT25), .B(G183gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(KEYINPUT26), .B(G190gat), .ZN(new_n435_));
  OAI21_X1  g234(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G169gat), .A2(G176gat), .ZN(new_n438_));
  AOI22_X1  g237(.A1(new_n434_), .A2(new_n435_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n432_), .A2(new_n433_), .A3(new_n439_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(G169gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n423_), .A2(new_n425_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(KEYINPUT23), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT23), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n421_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n444_), .A2(new_n446_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(G183gat), .A2(G190gat), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n442_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n419_), .B1(new_n440_), .B2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G226gat), .A2(G233gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(KEYINPUT19), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT20), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT99), .ZN(new_n455_));
  INV_X1    g254(.A(G183gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT25), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT25), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(G183gat), .ZN(new_n459_));
  INV_X1    g258(.A(G190gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT26), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT26), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(G190gat), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n457_), .A2(new_n459_), .A3(new_n461_), .A4(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n437_), .A2(new_n438_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n464_), .A2(new_n465_), .A3(new_n420_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n455_), .B1(new_n447_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n446_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n468_), .B1(new_n443_), .B2(KEYINPUT23), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n469_), .A2(new_n439_), .A3(KEYINPUT99), .A4(new_n420_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n422_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n424_), .B1(G183gat), .B2(G190gat), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n421_), .A2(KEYINPUT84), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n445_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n471_), .B1(new_n474_), .B2(KEYINPUT85), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n426_), .A2(new_n427_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n448_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n442_), .ZN(new_n478_));
  OAI211_X1 g277(.A(new_n467_), .B(new_n470_), .C1(new_n477_), .C2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n408_), .A2(new_n394_), .ZN(new_n480_));
  AND2_X1   g279(.A1(new_n408_), .A2(new_n414_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n480_), .B1(new_n481_), .B2(new_n394_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n454_), .B1(new_n479_), .B2(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n450_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT100), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n453_), .B1(new_n479_), .B2(new_n482_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n440_), .A2(new_n419_), .A3(new_n449_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  AOI22_X1  g287(.A1(new_n484_), .A2(new_n485_), .B1(new_n488_), .B2(new_n452_), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT100), .B1(new_n450_), .B2(new_n483_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n393_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n488_), .A2(new_n452_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n440_), .A2(new_n449_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(new_n482_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n454_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n474_), .A2(KEYINPUT85), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n496_), .A2(new_n476_), .A3(new_n422_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n448_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n478_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n467_), .A2(new_n470_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n495_), .B1(new_n501_), .B2(new_n419_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n494_), .A2(new_n485_), .A3(new_n502_), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n492_), .A2(new_n503_), .A3(new_n490_), .A4(new_n393_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n388_), .B1(new_n491_), .B2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT104), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n489_), .A2(new_n507_), .A3(new_n393_), .A4(new_n490_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n504_), .A2(KEYINPUT104), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n498_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(new_n442_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n469_), .A2(new_n439_), .A3(new_n420_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n419_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n513_));
  XOR2_X1   g312(.A(KEYINPUT103), .B(KEYINPUT20), .Z(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n452_), .B1(new_n450_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n452_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n486_), .A2(new_n487_), .A3(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n393_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n388_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n508_), .A2(new_n509_), .A3(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G78gat), .B(G106gat), .ZN(new_n523_));
  XOR2_X1   g322(.A(new_n523_), .B(KEYINPUT97), .Z(new_n524_));
  INV_X1    g323(.A(KEYINPUT29), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT90), .ZN(new_n526_));
  INV_X1    g325(.A(G155gat), .ZN(new_n527_));
  INV_X1    g326(.A(G162gat), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n526_), .A2(new_n527_), .A3(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT90), .B1(G155gat), .B2(G162gat), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G155gat), .A2(G162gat), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(KEYINPUT1), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT1), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n534_), .A2(G155gat), .A3(G162gat), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n531_), .A2(new_n533_), .A3(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G141gat), .B(G148gat), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT3), .ZN(new_n539_));
  INV_X1    g338(.A(G141gat), .ZN(new_n540_));
  INV_X1    g339(.A(G148gat), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n539_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G141gat), .A2(G148gat), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT2), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n546_));
  OAI21_X1  g345(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n542_), .A2(new_n545_), .A3(new_n546_), .A4(new_n547_), .ZN(new_n548_));
  AOI22_X1  g347(.A1(new_n529_), .A2(new_n530_), .B1(G155gat), .B2(G162gat), .ZN(new_n549_));
  AOI22_X1  g348(.A1(new_n536_), .A2(new_n538_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  OAI22_X1  g349(.A1(new_n415_), .A2(new_n418_), .B1(new_n525_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT94), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n552_), .A2(G233gat), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(G233gat), .ZN(new_n554_));
  AND2_X1   g353(.A1(KEYINPUT93), .A2(G228gat), .ZN(new_n555_));
  NOR2_X1   g354(.A1(KEYINPUT93), .A2(G228gat), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n553_), .B(new_n554_), .C1(new_n555_), .C2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n551_), .A2(new_n558_), .ZN(new_n559_));
  OAI221_X1 g358(.A(new_n557_), .B1(new_n525_), .B2(new_n550_), .C1(new_n415_), .C2(new_n418_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n524_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n559_), .A2(new_n560_), .A3(new_n524_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(G22gat), .B(G50gat), .Z(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n536_), .A2(new_n538_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n549_), .A2(new_n548_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n567_), .A2(new_n568_), .A3(new_n525_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(KEYINPUT91), .B(KEYINPUT28), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n570_), .B1(new_n550_), .B2(new_n525_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n566_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n569_), .A2(new_n571_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n550_), .A2(new_n525_), .A3(new_n570_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n575_), .A2(new_n565_), .A3(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(KEYINPUT92), .B1(new_n574_), .B2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n574_), .A2(KEYINPUT92), .A3(new_n577_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n559_), .A2(new_n560_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(KEYINPUT98), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT98), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n559_), .A2(new_n584_), .A3(new_n560_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n583_), .A2(new_n523_), .A3(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n574_), .A2(new_n577_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n563_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  AOI22_X1  g388(.A1(new_n564_), .A2(new_n581_), .B1(new_n586_), .B2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G1gat), .B(G29gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(G85gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(KEYINPUT0), .B(G57gat), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n592_), .B(new_n593_), .Z(new_n594_));
  NAND2_X1  g393(.A1(G225gat), .A2(G233gat), .ZN(new_n595_));
  INV_X1    g394(.A(G134gat), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(G127gat), .ZN(new_n597_));
  INV_X1    g396(.A(G127gat), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(G134gat), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(G120gat), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(G113gat), .ZN(new_n602_));
  INV_X1    g401(.A(G113gat), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(G120gat), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n600_), .A2(new_n605_), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n597_), .A2(new_n599_), .A3(new_n602_), .A4(new_n604_), .ZN(new_n607_));
  AND3_X1   g406(.A1(new_n606_), .A2(KEYINPUT89), .A3(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(KEYINPUT89), .B1(new_n606_), .B2(new_n607_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n549_), .A2(new_n548_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n533_), .A2(new_n535_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n537_), .B1(new_n611_), .B2(new_n531_), .ZN(new_n612_));
  OAI22_X1  g411(.A1(new_n608_), .A2(new_n609_), .B1(new_n610_), .B2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n606_), .A2(new_n607_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n550_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n613_), .A2(KEYINPUT4), .A3(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT102), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT4), .ZN(new_n618_));
  INV_X1    g417(.A(new_n608_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n609_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n550_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  AOI22_X1  g420(.A1(new_n616_), .A2(new_n617_), .B1(new_n618_), .B2(new_n621_), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n613_), .A2(new_n615_), .A3(KEYINPUT102), .A4(KEYINPUT4), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n595_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n613_), .A2(new_n615_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n595_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n594_), .B1(new_n624_), .B2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n616_), .A2(new_n617_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n621_), .A2(new_n618_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n629_), .A2(new_n623_), .A3(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(new_n626_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n594_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n627_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n632_), .A2(new_n633_), .A3(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n628_), .A2(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n590_), .A2(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n506_), .A2(new_n522_), .A3(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n492_), .A2(new_n503_), .A3(new_n490_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(new_n520_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n629_), .A2(new_n595_), .A3(new_n630_), .A4(new_n623_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n594_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(KEYINPUT33), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n628_), .A2(new_n644_), .ZN(new_n645_));
  OAI211_X1 g444(.A(KEYINPUT33), .B(new_n594_), .C1(new_n624_), .C2(new_n627_), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n640_), .A2(new_n645_), .A3(new_n504_), .A4(new_n646_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n393_), .A2(KEYINPUT32), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n519_), .A2(new_n648_), .ZN(new_n649_));
  OAI211_X1 g448(.A(new_n636_), .B(new_n649_), .C1(new_n639_), .C2(new_n648_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n647_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n563_), .ZN(new_n652_));
  AND3_X1   g451(.A1(new_n574_), .A2(KEYINPUT92), .A3(new_n577_), .ZN(new_n653_));
  OAI22_X1  g452(.A1(new_n652_), .A2(new_n561_), .B1(new_n653_), .B2(new_n578_), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n559_), .A2(new_n584_), .A3(new_n560_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n584_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n523_), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n655_), .A2(new_n656_), .A3(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n654_), .B1(new_n658_), .B2(new_n588_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n638_), .B1(new_n651_), .B2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT88), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n440_), .A2(KEYINPUT30), .A3(new_n449_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(KEYINPUT30), .B1(new_n440_), .B2(new_n449_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n661_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT30), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n493_), .A2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n667_), .A2(KEYINPUT88), .A3(new_n662_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(G227gat), .A2(G233gat), .ZN(new_n669_));
  INV_X1    g468(.A(G15gat), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n669_), .B(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(G71gat), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(new_n229_), .ZN(new_n673_));
  XOR2_X1   g472(.A(KEYINPUT87), .B(G43gat), .Z(new_n674_));
  XNOR2_X1  g473(.A(new_n673_), .B(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n665_), .A2(new_n668_), .A3(new_n675_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n673_), .B(new_n674_), .Z(new_n677_));
  NAND4_X1  g476(.A1(new_n677_), .A2(KEYINPUT88), .A3(new_n667_), .A4(new_n662_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n619_), .A2(new_n620_), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n679_), .B(KEYINPUT31), .Z(new_n680_));
  AND3_X1   g479(.A1(new_n676_), .A2(new_n678_), .A3(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n680_), .B1(new_n676_), .B2(new_n678_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n506_), .A2(new_n522_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n659_), .A2(new_n636_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n685_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n686_));
  OAI21_X1  g485(.A(KEYINPUT105), .B1(new_n684_), .B2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n586_), .A2(new_n589_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n688_), .A2(new_n628_), .A3(new_n635_), .A4(new_n654_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n676_), .A2(new_n678_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n680_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n676_), .A2(new_n678_), .A3(new_n680_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n689_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT105), .ZN(new_n695_));
  NAND4_X1  g494(.A1(new_n694_), .A2(new_n695_), .A3(new_n506_), .A4(new_n522_), .ZN(new_n696_));
  AOI22_X1  g495(.A1(new_n660_), .A2(new_n683_), .B1(new_n687_), .B2(new_n696_), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n351_), .A2(new_n387_), .A3(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n698_), .A2(new_n636_), .A3(new_n291_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT38), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n687_), .A2(new_n696_), .ZN(new_n701_));
  AND3_X1   g500(.A1(new_n506_), .A2(new_n522_), .A3(new_n637_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n659_), .B1(new_n647_), .B2(new_n650_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n683_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n701_), .A2(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n387_), .B1(new_n347_), .B2(new_n349_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n281_), .A2(new_n284_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n329_), .A2(new_n707_), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n705_), .A2(new_n706_), .A3(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n636_), .ZN(new_n711_));
  OAI21_X1  g510(.A(G1gat), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n700_), .A2(new_n712_), .ZN(G1324gat));
  NAND3_X1  g512(.A1(new_n698_), .A2(new_n292_), .A3(new_n684_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n684_), .ZN(new_n715_));
  OAI21_X1  g514(.A(G8gat), .B1(new_n710_), .B2(new_n715_), .ZN(new_n716_));
  XOR2_X1   g515(.A(KEYINPUT106), .B(KEYINPUT39), .Z(new_n717_));
  AND2_X1   g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n716_), .A2(new_n717_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n714_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT40), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n720_), .B(new_n721_), .ZN(G1325gat));
  INV_X1    g521(.A(new_n683_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n670_), .B1(new_n709_), .B2(new_n723_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT41), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n698_), .A2(new_n670_), .A3(new_n723_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1326gat));
  INV_X1    g526(.A(G22gat), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n698_), .A2(new_n728_), .A3(new_n659_), .ZN(new_n729_));
  OAI21_X1  g528(.A(G22gat), .B1(new_n710_), .B2(new_n590_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n730_), .A2(KEYINPUT42), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n730_), .A2(KEYINPUT42), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n729_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT107), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n733_), .B(new_n734_), .ZN(G1327gat));
  INV_X1    g534(.A(KEYINPUT79), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n328_), .B(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n707_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n705_), .A2(new_n706_), .A3(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT109), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT109), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n705_), .A2(new_n739_), .A3(new_n706_), .A4(new_n742_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n741_), .A2(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(G29gat), .B1(new_n744_), .B2(new_n636_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT43), .ZN(new_n746_));
  OAI211_X1 g545(.A(new_n705_), .B(new_n290_), .C1(KEYINPUT108), .C2(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n290_), .B2(KEYINPUT108), .ZN(new_n748_));
  INV_X1    g547(.A(new_n290_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n748_), .B1(new_n697_), .B2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n747_), .A2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n706_), .A2(new_n329_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(KEYINPUT44), .B1(new_n751_), .B2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT44), .ZN(new_n755_));
  AOI211_X1 g554(.A(new_n755_), .B(new_n752_), .C1(new_n747_), .C2(new_n750_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n754_), .A2(new_n756_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n636_), .A2(G29gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n745_), .B1(new_n757_), .B2(new_n758_), .ZN(G1328gat));
  NAND2_X1  g558(.A1(KEYINPUT110), .A2(KEYINPUT46), .ZN(new_n760_));
  NOR2_X1   g559(.A1(KEYINPUT110), .A2(KEYINPUT46), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n715_), .A2(G36gat), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n741_), .A2(new_n743_), .A3(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT45), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT45), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n741_), .A2(new_n765_), .A3(new_n743_), .A4(new_n762_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n761_), .B1(new_n764_), .B2(new_n766_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n754_), .A2(new_n756_), .A3(new_n715_), .ZN(new_n768_));
  INV_X1    g567(.A(G36gat), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n760_), .B(new_n767_), .C1(new_n768_), .C2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n751_), .A2(new_n753_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(new_n755_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n751_), .A2(KEYINPUT44), .A3(new_n753_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n773_), .A2(new_n684_), .A3(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(G36gat), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n760_), .B1(new_n776_), .B2(new_n767_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n771_), .A2(new_n777_), .ZN(G1329gat));
  AND3_X1   g577(.A1(new_n757_), .A2(G43gat), .A3(new_n723_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n741_), .A2(new_n723_), .A3(new_n743_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(KEYINPUT111), .B(G43gat), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n780_), .A2(KEYINPUT112), .A3(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT112), .B1(new_n780_), .B2(new_n781_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  OAI21_X1  g583(.A(KEYINPUT47), .B1(new_n779_), .B2(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n757_), .A2(G43gat), .A3(new_n723_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT47), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n786_), .B(new_n787_), .C1(new_n783_), .C2(new_n782_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n785_), .A2(new_n788_), .ZN(G1330gat));
  AOI21_X1  g588(.A(G50gat), .B1(new_n744_), .B2(new_n659_), .ZN(new_n790_));
  AND2_X1   g589(.A1(new_n659_), .A2(G50gat), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n757_), .B2(new_n791_), .ZN(G1331gat));
  NOR2_X1   g591(.A1(new_n350_), .A2(new_n386_), .ZN(new_n793_));
  AND3_X1   g592(.A1(new_n793_), .A2(new_n705_), .A3(new_n330_), .ZN(new_n794_));
  AOI21_X1  g593(.A(G57gat), .B1(new_n794_), .B2(new_n636_), .ZN(new_n795_));
  XOR2_X1   g594(.A(new_n795_), .B(KEYINPUT113), .Z(new_n796_));
  AND3_X1   g595(.A1(new_n793_), .A2(new_n705_), .A3(new_n708_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(KEYINPUT114), .B(G57gat), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n711_), .A2(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n796_), .B1(new_n797_), .B2(new_n799_), .ZN(G1332gat));
  INV_X1    g599(.A(G64gat), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n801_), .B1(new_n797_), .B2(new_n684_), .ZN(new_n802_));
  XOR2_X1   g601(.A(new_n802_), .B(KEYINPUT48), .Z(new_n803_));
  NAND3_X1  g602(.A1(new_n794_), .A2(new_n801_), .A3(new_n684_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(G1333gat));
  INV_X1    g604(.A(G71gat), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n806_), .B1(new_n797_), .B2(new_n723_), .ZN(new_n807_));
  XOR2_X1   g606(.A(KEYINPUT115), .B(KEYINPUT49), .Z(new_n808_));
  XNOR2_X1  g607(.A(new_n807_), .B(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n794_), .A2(new_n806_), .A3(new_n723_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(G1334gat));
  INV_X1    g610(.A(G78gat), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n812_), .B1(new_n797_), .B2(new_n659_), .ZN(new_n813_));
  XOR2_X1   g612(.A(new_n813_), .B(KEYINPUT50), .Z(new_n814_));
  NAND3_X1  g613(.A1(new_n794_), .A2(new_n812_), .A3(new_n659_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(G1335gat));
  AND3_X1   g615(.A1(new_n793_), .A2(new_n705_), .A3(new_n739_), .ZN(new_n817_));
  AOI21_X1  g616(.A(G85gat), .B1(new_n817_), .B2(new_n636_), .ZN(new_n818_));
  XOR2_X1   g617(.A(new_n818_), .B(KEYINPUT116), .Z(new_n819_));
  NAND2_X1  g618(.A1(new_n793_), .A2(new_n329_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n820_), .B1(new_n747_), .B2(new_n750_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n822_), .A2(new_n214_), .A3(new_n711_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n819_), .A2(new_n823_), .ZN(G1336gat));
  OAI21_X1  g623(.A(G92gat), .B1(new_n822_), .B2(new_n715_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n817_), .A2(new_n215_), .A3(new_n684_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(G1337gat));
  NAND4_X1  g626(.A1(new_n817_), .A2(new_n207_), .A3(new_n209_), .A4(new_n723_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n822_), .A2(new_n683_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n828_), .B1(new_n829_), .B2(new_n229_), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n830_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g630(.A1(new_n817_), .A2(new_n208_), .A3(new_n659_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n208_), .B1(new_n821_), .B2(new_n659_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT52), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n833_), .A2(new_n834_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n832_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(KEYINPUT53), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT53), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n839_), .B(new_n832_), .C1(new_n835_), .C2(new_n836_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n840_), .ZN(G1339gat));
  INV_X1    g640(.A(KEYINPUT59), .ZN(new_n842_));
  XOR2_X1   g641(.A(KEYINPUT117), .B(KEYINPUT54), .Z(new_n843_));
  XNOR2_X1  g642(.A(new_n843_), .B(KEYINPUT118), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n844_), .B1(new_n351_), .B2(new_n386_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT118), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n843_), .A2(new_n846_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n330_), .A2(new_n387_), .A3(new_n350_), .A4(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n845_), .A2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n353_), .A2(new_n359_), .A3(new_n362_), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n850_), .B(new_n383_), .C1(new_n379_), .C2(new_n359_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n377_), .A2(new_n851_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n340_), .A2(new_n344_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n334_), .A2(new_n336_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT119), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n335_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n334_), .A2(KEYINPUT119), .A3(new_n336_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n857_), .A2(new_n858_), .A3(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT120), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n857_), .A2(KEYINPUT120), .A3(new_n858_), .A4(new_n859_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(KEYINPUT121), .A2(KEYINPUT55), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n337_), .A2(KEYINPUT121), .A3(KEYINPUT55), .ZN(new_n865_));
  NAND2_X1  g664(.A1(KEYINPUT121), .A2(KEYINPUT55), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n334_), .A2(new_n335_), .A3(new_n336_), .A4(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n864_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n862_), .A2(new_n863_), .A3(new_n868_), .ZN(new_n869_));
  AND3_X1   g668(.A1(new_n869_), .A2(KEYINPUT56), .A3(new_n344_), .ZN(new_n870_));
  AOI21_X1  g669(.A(KEYINPUT56), .B1(new_n869_), .B2(new_n344_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n854_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(KEYINPUT122), .B(KEYINPUT58), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n749_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT58), .ZN(new_n875_));
  OAI21_X1  g674(.A(KEYINPUT123), .B1(new_n872_), .B2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n871_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n869_), .A2(KEYINPUT56), .A3(new_n344_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT123), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n879_), .A2(new_n880_), .A3(KEYINPUT58), .A4(new_n854_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n874_), .A2(new_n876_), .A3(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n853_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n386_), .A2(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n884_), .B1(new_n877_), .B2(new_n878_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n852_), .A2(new_n345_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n738_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT57), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n853_), .B1(new_n377_), .B2(new_n385_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n890_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n886_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n893_), .A2(KEYINPUT57), .A3(new_n738_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n882_), .A2(new_n889_), .A3(new_n894_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n849_), .B1(new_n895_), .B2(new_n329_), .ZN(new_n896_));
  NOR4_X1   g695(.A1(new_n684_), .A2(new_n683_), .A3(new_n711_), .A4(new_n659_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n842_), .B1(new_n896_), .B2(new_n898_), .ZN(new_n899_));
  AOI21_X1  g698(.A(KEYINPUT57), .B1(new_n893_), .B2(new_n738_), .ZN(new_n900_));
  AOI211_X1 g699(.A(new_n888_), .B(new_n707_), .C1(new_n891_), .C2(new_n892_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n737_), .B1(new_n902_), .B2(new_n882_), .ZN(new_n903_));
  OAI211_X1 g702(.A(KEYINPUT59), .B(new_n897_), .C1(new_n903_), .C2(new_n849_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n899_), .A2(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n603_), .B1(new_n386_), .B2(KEYINPUT124), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n906_), .B1(KEYINPUT124), .B2(new_n603_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n896_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n908_), .A2(new_n386_), .A3(new_n897_), .ZN(new_n909_));
  AOI22_X1  g708(.A1(new_n905_), .A2(new_n907_), .B1(new_n909_), .B2(new_n603_), .ZN(G1340gat));
  NOR2_X1   g709(.A1(new_n896_), .A2(new_n898_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n601_), .B1(new_n350_), .B2(KEYINPUT60), .ZN(new_n912_));
  OAI211_X1 g711(.A(new_n911_), .B(new_n912_), .C1(KEYINPUT60), .C2(new_n601_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n350_), .B1(new_n899_), .B2(new_n904_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n913_), .B1(new_n914_), .B2(new_n601_), .ZN(G1341gat));
  NAND3_X1  g714(.A1(new_n911_), .A2(new_n598_), .A3(new_n737_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n329_), .B1(new_n899_), .B2(new_n904_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n917_), .B2(new_n598_), .ZN(G1342gat));
  NAND3_X1  g717(.A1(new_n911_), .A2(new_n596_), .A3(new_n707_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n749_), .B1(new_n899_), .B2(new_n904_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n919_), .B1(new_n920_), .B2(new_n596_), .ZN(G1343gat));
  NAND4_X1  g720(.A1(new_n715_), .A2(new_n636_), .A3(new_n659_), .A4(new_n683_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n896_), .A2(new_n922_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(KEYINPUT125), .B(G141gat), .ZN(new_n924_));
  AND3_X1   g723(.A1(new_n923_), .A2(new_n386_), .A3(new_n924_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n924_), .B1(new_n923_), .B2(new_n386_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n925_), .A2(new_n926_), .ZN(G1344gat));
  INV_X1    g726(.A(new_n923_), .ZN(new_n928_));
  OAI21_X1  g727(.A(G148gat), .B1(new_n928_), .B2(new_n350_), .ZN(new_n929_));
  INV_X1    g728(.A(new_n350_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n923_), .A2(new_n541_), .A3(new_n930_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n929_), .A2(new_n931_), .ZN(G1345gat));
  XNOR2_X1  g731(.A(KEYINPUT61), .B(G155gat), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n933_), .B1(new_n928_), .B2(new_n329_), .ZN(new_n934_));
  INV_X1    g733(.A(new_n933_), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n923_), .A2(new_n737_), .A3(new_n935_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n934_), .A2(new_n936_), .ZN(G1346gat));
  OAI21_X1  g736(.A(G162gat), .B1(new_n928_), .B2(new_n749_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n923_), .A2(new_n528_), .A3(new_n707_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n938_), .A2(new_n939_), .ZN(G1347gat));
  NOR2_X1   g739(.A1(new_n715_), .A2(new_n686_), .ZN(new_n941_));
  INV_X1    g740(.A(new_n941_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n896_), .A2(new_n942_), .ZN(new_n943_));
  XNOR2_X1  g742(.A(KEYINPUT22), .B(G169gat), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n386_), .A2(new_n944_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(new_n945_), .B(KEYINPUT126), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n943_), .A2(new_n946_), .ZN(new_n947_));
  OAI211_X1 g746(.A(new_n386_), .B(new_n941_), .C1(new_n903_), .C2(new_n849_), .ZN(new_n948_));
  INV_X1    g747(.A(KEYINPUT62), .ZN(new_n949_));
  AND3_X1   g748(.A1(new_n948_), .A2(new_n949_), .A3(G169gat), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n949_), .B1(new_n948_), .B2(G169gat), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n947_), .B1(new_n950_), .B2(new_n951_), .ZN(G1348gat));
  NOR3_X1   g751(.A1(new_n896_), .A2(new_n350_), .A3(new_n942_), .ZN(new_n953_));
  INV_X1    g752(.A(G176gat), .ZN(new_n954_));
  XNOR2_X1  g753(.A(new_n953_), .B(new_n954_), .ZN(G1349gat));
  NOR4_X1   g754(.A1(new_n896_), .A2(new_n434_), .A3(new_n329_), .A4(new_n942_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n943_), .A2(new_n737_), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n956_), .B1(new_n456_), .B2(new_n957_), .ZN(G1350gat));
  NAND3_X1  g757(.A1(new_n943_), .A2(new_n435_), .A3(new_n707_), .ZN(new_n959_));
  NOR3_X1   g758(.A1(new_n896_), .A2(new_n749_), .A3(new_n942_), .ZN(new_n960_));
  OAI21_X1  g759(.A(new_n959_), .B1(new_n960_), .B2(new_n460_), .ZN(G1351gat));
  NAND3_X1  g760(.A1(new_n684_), .A2(new_n637_), .A3(new_n683_), .ZN(new_n962_));
  NOR2_X1   g761(.A1(new_n896_), .A2(new_n962_), .ZN(new_n963_));
  AND3_X1   g762(.A1(new_n963_), .A2(G197gat), .A3(new_n386_), .ZN(new_n964_));
  AOI21_X1  g763(.A(G197gat), .B1(new_n963_), .B2(new_n386_), .ZN(new_n965_));
  NOR2_X1   g764(.A1(new_n964_), .A2(new_n965_), .ZN(G1352gat));
  OR2_X1    g765(.A1(new_n896_), .A2(new_n962_), .ZN(new_n967_));
  OAI211_X1 g766(.A(KEYINPUT127), .B(G204gat), .C1(new_n967_), .C2(new_n350_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n969_));
  NAND3_X1  g768(.A1(new_n963_), .A2(new_n930_), .A3(new_n969_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n968_), .A2(new_n970_), .ZN(G1353gat));
  OR2_X1    g770(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n972_));
  AOI21_X1  g771(.A(new_n972_), .B1(new_n963_), .B2(new_n737_), .ZN(new_n973_));
  NOR2_X1   g772(.A1(new_n967_), .A2(new_n329_), .ZN(new_n974_));
  XOR2_X1   g773(.A(KEYINPUT63), .B(G211gat), .Z(new_n975_));
  AOI21_X1  g774(.A(new_n973_), .B1(new_n974_), .B2(new_n975_), .ZN(G1354gat));
  OAI21_X1  g775(.A(G218gat), .B1(new_n967_), .B2(new_n749_), .ZN(new_n977_));
  NAND3_X1  g776(.A1(new_n963_), .A2(new_n402_), .A3(new_n707_), .ZN(new_n978_));
  NAND2_X1  g777(.A1(new_n977_), .A2(new_n978_), .ZN(G1355gat));
endmodule


