//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 0 0 0 1 0 0 1 1 0 1 1 0 0 1 0 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 0 1 0 1 1 1 0 0 0 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n688_, new_n689_, new_n690_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n882_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n907_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n916_, new_n917_, new_n918_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G134gat), .B(G162gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT36), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT66), .B(KEYINPUT6), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G85gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT9), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n209_), .A2(new_n210_), .A3(G92gat), .ZN(new_n211_));
  XOR2_X1   g010(.A(G85gat), .B(G92gat), .Z(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT9), .ZN(new_n213_));
  XOR2_X1   g012(.A(KEYINPUT10), .B(G99gat), .Z(new_n214_));
  INV_X1    g013(.A(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n208_), .A2(new_n211_), .A3(new_n213_), .A4(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(G99gat), .A2(G106gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT7), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n208_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(new_n212_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT8), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT8), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n221_), .A2(new_n224_), .A3(new_n212_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n218_), .B1(new_n223_), .B2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G29gat), .B(G36gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(KEYINPUT72), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G43gat), .B(G50gat), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  OR2_X1    g030(.A1(new_n227_), .A2(KEYINPUT72), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n227_), .A2(KEYINPUT72), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n232_), .A2(new_n233_), .A3(new_n229_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n231_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT35), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G232gat), .A2(G233gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT34), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  AOI22_X1  g039(.A1(new_n226_), .A2(new_n236_), .B1(new_n237_), .B2(new_n240_), .ZN(new_n241_));
  AND3_X1   g040(.A1(new_n221_), .A2(new_n224_), .A3(new_n212_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n224_), .B1(new_n221_), .B2(new_n212_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n217_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT69), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  OAI211_X1 g045(.A(KEYINPUT69), .B(new_n217_), .C1(new_n242_), .C2(new_n243_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT15), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n235_), .A2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n231_), .A2(KEYINPUT15), .A3(new_n234_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n241_), .B1(new_n248_), .B2(new_n253_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n240_), .A2(new_n237_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  OAI221_X1 g055(.A(new_n241_), .B1(new_n237_), .B2(new_n240_), .C1(new_n248_), .C2(new_n253_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n205_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT73), .B(KEYINPUT36), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n204_), .A2(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n256_), .A2(new_n257_), .A3(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT74), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n256_), .A2(new_n257_), .A3(KEYINPUT74), .A4(new_n260_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n258_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT37), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G230gat), .A2(G233gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT64), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G57gat), .B(G64gat), .ZN(new_n270_));
  AND2_X1   g069(.A1(new_n270_), .A2(KEYINPUT67), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n270_), .A2(KEYINPUT67), .ZN(new_n272_));
  OR3_X1    g071(.A1(new_n271_), .A2(new_n272_), .A3(KEYINPUT11), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT11), .B1(new_n271_), .B2(new_n272_), .ZN(new_n274_));
  XOR2_X1   g073(.A(G71gat), .B(G78gat), .Z(new_n275_));
  NAND3_X1  g074(.A1(new_n273_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n274_), .A2(new_n275_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n226_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n278_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n244_), .A2(new_n280_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n269_), .B1(new_n279_), .B2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT68), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  OAI211_X1 g083(.A(KEYINPUT68), .B(new_n269_), .C1(new_n279_), .C2(new_n281_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  AND3_X1   g085(.A1(new_n276_), .A2(KEYINPUT12), .A3(new_n277_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n246_), .A2(new_n247_), .A3(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT70), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n244_), .A2(new_n280_), .ZN(new_n290_));
  XOR2_X1   g089(.A(KEYINPUT71), .B(KEYINPUT12), .Z(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT70), .ZN(new_n293_));
  NAND4_X1  g092(.A1(new_n246_), .A2(new_n293_), .A3(new_n287_), .A4(new_n247_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n281_), .A2(new_n269_), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n289_), .A2(new_n292_), .A3(new_n294_), .A4(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n286_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G120gat), .B(G148gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT5), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G176gat), .B(G204gat), .ZN(new_n300_));
  XOR2_X1   g099(.A(new_n299_), .B(new_n300_), .Z(new_n301_));
  NAND2_X1  g100(.A1(new_n297_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n301_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n286_), .A2(new_n296_), .A3(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(KEYINPUT13), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G231gat), .A2(G233gat), .ZN(new_n307_));
  XOR2_X1   g106(.A(new_n278_), .B(new_n307_), .Z(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT75), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G15gat), .B(G22gat), .ZN(new_n310_));
  INV_X1    g109(.A(G1gat), .ZN(new_n311_));
  INV_X1    g110(.A(G8gat), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT14), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n310_), .A2(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G1gat), .B(G8gat), .ZN(new_n315_));
  XOR2_X1   g114(.A(new_n314_), .B(new_n315_), .Z(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n309_), .B(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G127gat), .B(G155gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT16), .ZN(new_n320_));
  XOR2_X1   g119(.A(G183gat), .B(G211gat), .Z(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT17), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n318_), .A2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n322_), .B(KEYINPUT17), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n325_), .B1(new_n318_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n267_), .A2(new_n306_), .A3(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G225gat), .A2(G233gat), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  OR2_X1    g132(.A1(G155gat), .A2(G162gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G155gat), .A2(G162gat), .ZN(new_n335_));
  AND2_X1   g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT2), .ZN(new_n337_));
  AND3_X1   g136(.A1(KEYINPUT86), .A2(G141gat), .A3(G148gat), .ZN(new_n338_));
  AOI21_X1  g137(.A(KEYINPUT86), .B1(G141gat), .B2(G148gat), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n337_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  NOR4_X1   g139(.A1(KEYINPUT88), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT88), .ZN(new_n342_));
  NOR2_X1   g141(.A1(G141gat), .A2(G148gat), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT3), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n342_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n340_), .B1(new_n341_), .B2(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT89), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n350_));
  NAND4_X1  g149(.A1(KEYINPUT89), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n349_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n336_), .B1(new_n346_), .B2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT1), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n334_), .A2(new_n354_), .A3(new_n335_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G141gat), .A2(G148gat), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT86), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(KEYINPUT86), .A2(G141gat), .A3(G148gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n355_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT87), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n343_), .A2(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT87), .B1(G141gat), .B2(G148gat), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n363_), .B(new_n364_), .C1(new_n354_), .C2(new_n335_), .ZN(new_n365_));
  OR2_X1    g164(.A1(new_n361_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n353_), .A2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G113gat), .B(G120gat), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(G134gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(G127gat), .ZN(new_n371_));
  INV_X1    g170(.A(G127gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(G134gat), .ZN(new_n373_));
  AND3_X1   g172(.A1(new_n371_), .A2(new_n373_), .A3(KEYINPUT84), .ZN(new_n374_));
  AOI21_X1  g173(.A(KEYINPUT84), .B1(new_n371_), .B2(new_n373_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n369_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n371_), .A2(new_n373_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT84), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n371_), .A2(new_n373_), .A3(KEYINPUT84), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n379_), .A2(new_n380_), .A3(new_n368_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n376_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n367_), .A2(new_n383_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n361_), .A2(new_n365_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n343_), .A2(new_n344_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(KEYINPUT88), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n343_), .A2(new_n342_), .A3(new_n344_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  AND3_X1   g188(.A1(new_n349_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n389_), .A2(new_n390_), .A3(new_n340_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n385_), .B1(new_n391_), .B2(new_n336_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(new_n382_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n384_), .A2(new_n393_), .A3(KEYINPUT4), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n382_), .B1(new_n353_), .B2(new_n366_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT4), .ZN(new_n396_));
  AOI21_X1  g195(.A(KEYINPUT100), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT100), .ZN(new_n398_));
  NOR4_X1   g197(.A1(new_n392_), .A2(new_n398_), .A3(new_n382_), .A4(KEYINPUT4), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n333_), .B(new_n394_), .C1(new_n397_), .C2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT102), .ZN(new_n401_));
  AND3_X1   g200(.A1(new_n353_), .A2(new_n382_), .A3(new_n366_), .ZN(new_n402_));
  NOR3_X1   g201(.A1(new_n402_), .A2(new_n395_), .A3(new_n333_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G1gat), .B(G29gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(G85gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT0), .B(G57gat), .ZN(new_n407_));
  XOR2_X1   g206(.A(new_n406_), .B(new_n407_), .Z(new_n408_));
  NAND4_X1  g207(.A1(new_n400_), .A2(new_n401_), .A3(new_n404_), .A4(new_n408_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n402_), .A2(new_n395_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n332_), .B1(new_n410_), .B2(KEYINPUT4), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n398_), .B1(new_n384_), .B2(KEYINPUT4), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n395_), .A2(KEYINPUT100), .A3(new_n396_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n403_), .B1(new_n411_), .B2(new_n414_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n409_), .B1(new_n415_), .B2(new_n408_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n401_), .B1(new_n415_), .B2(new_n408_), .ZN(new_n417_));
  OAI21_X1  g216(.A(KEYINPUT104), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  OR2_X1    g217(.A1(G183gat), .A2(G190gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G183gat), .A2(G190gat), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT23), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT81), .B(KEYINPUT23), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n419_), .B(new_n422_), .C1(new_n423_), .C2(new_n420_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G169gat), .A2(G176gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(KEYINPUT22), .B(G169gat), .ZN(new_n426_));
  INV_X1    g225(.A(G176gat), .ZN(new_n427_));
  AND3_X1   g226(.A1(new_n426_), .A2(KEYINPUT82), .A3(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(KEYINPUT82), .B1(new_n426_), .B2(new_n427_), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n424_), .B(new_n425_), .C1(new_n428_), .C2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT24), .ZN(new_n431_));
  INV_X1    g230(.A(G169gat), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n431_), .A2(new_n432_), .A3(new_n427_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n425_), .A2(KEYINPUT24), .ZN(new_n434_));
  NOR2_X1   g233(.A1(G169gat), .A2(G176gat), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n433_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT25), .B(G183gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(KEYINPUT26), .B(G190gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  AND2_X1   g239(.A1(G183gat), .A2(G190gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n421_), .A2(KEYINPUT81), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT81), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(KEYINPUT23), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n441_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n420_), .A2(KEYINPUT23), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n437_), .B(new_n440_), .C1(new_n445_), .C2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n430_), .A2(new_n447_), .ZN(new_n448_));
  XOR2_X1   g247(.A(G71gat), .B(G99gat), .Z(new_n449_));
  XOR2_X1   g248(.A(KEYINPUT83), .B(G43gat), .Z(new_n450_));
  XOR2_X1   g249(.A(new_n449_), .B(new_n450_), .Z(new_n451_));
  OR2_X1    g250(.A1(new_n448_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G227gat), .A2(G233gat), .ZN(new_n453_));
  INV_X1    g252(.A(G15gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(KEYINPUT30), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(KEYINPUT31), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n448_), .A2(new_n451_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n452_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n457_), .B1(new_n452_), .B2(new_n458_), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT85), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT31), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n456_), .B(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n458_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n448_), .A2(new_n451_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n464_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT85), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n467_), .A2(new_n468_), .A3(new_n459_), .ZN(new_n469_));
  AND3_X1   g268(.A1(new_n462_), .A2(new_n383_), .A3(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n383_), .B1(new_n462_), .B2(new_n469_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n400_), .A2(new_n404_), .A3(new_n408_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT102), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n400_), .A2(new_n404_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n408_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT104), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n474_), .A2(new_n477_), .A3(new_n478_), .A4(new_n409_), .ZN(new_n479_));
  AND3_X1   g278(.A1(new_n418_), .A2(new_n472_), .A3(new_n479_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n367_), .A2(KEYINPUT29), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT28), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G22gat), .B(G50gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT28), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n481_), .B(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n483_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n484_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(G233gat), .ZN(new_n490_));
  AND2_X1   g289(.A1(new_n490_), .A2(KEYINPUT90), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n490_), .A2(KEYINPUT90), .ZN(new_n492_));
  OAI21_X1  g291(.A(G228gat), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT29), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n495_), .B1(new_n353_), .B2(new_n366_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT21), .ZN(new_n497_));
  INV_X1    g296(.A(G218gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(G211gat), .ZN(new_n499_));
  INV_X1    g298(.A(G211gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(G218gat), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n497_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n502_));
  AND2_X1   g301(.A1(G197gat), .A2(G204gat), .ZN(new_n503_));
  NOR2_X1   g302(.A1(G197gat), .A2(G204gat), .ZN(new_n504_));
  OAI21_X1  g303(.A(KEYINPUT91), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  OR2_X1    g304(.A1(G197gat), .A2(G204gat), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT91), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G197gat), .A2(G204gat), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n506_), .A2(new_n507_), .A3(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n502_), .A2(new_n505_), .A3(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT92), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT92), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n502_), .A2(new_n509_), .A3(new_n505_), .A4(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n506_), .A2(KEYINPUT21), .A3(new_n508_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n499_), .A2(new_n501_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n506_), .A2(new_n508_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n515_), .B1(new_n497_), .B2(new_n516_), .ZN(new_n517_));
  AOI22_X1  g316(.A1(new_n511_), .A2(new_n513_), .B1(new_n514_), .B2(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n494_), .B1(new_n496_), .B2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n511_), .A2(new_n513_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n517_), .A2(new_n514_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n522_), .B(new_n493_), .C1(new_n495_), .C2(new_n392_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G78gat), .B(G106gat), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n519_), .A2(new_n523_), .A3(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n525_), .B1(new_n519_), .B2(new_n523_), .ZN(new_n528_));
  NOR3_X1   g327(.A1(new_n489_), .A2(new_n527_), .A3(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n526_), .B1(new_n528_), .B2(KEYINPUT93), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT93), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n519_), .A2(new_n523_), .A3(new_n531_), .A4(new_n525_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(new_n489_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT94), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n533_), .A2(new_n489_), .A3(KEYINPUT94), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n529_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G8gat), .B(G36gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G64gat), .B(G92gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT20), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n420_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n422_), .ZN(new_n547_));
  NOR3_X1   g346(.A1(new_n436_), .A2(new_n546_), .A3(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT96), .ZN(new_n549_));
  INV_X1    g348(.A(G183gat), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n550_), .A2(KEYINPUT25), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n550_), .A2(KEYINPUT25), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n549_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n438_), .A2(KEYINPUT96), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n553_), .A2(new_n554_), .A3(new_n439_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n419_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n425_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n557_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n558_));
  AOI22_X1  g357(.A1(new_n548_), .A2(new_n555_), .B1(new_n556_), .B2(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n545_), .B1(new_n518_), .B2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n522_), .A2(new_n448_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G226gat), .A2(G233gat), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n562_), .B(KEYINPUT19), .Z(new_n563_));
  NAND3_X1  g362(.A1(new_n560_), .A2(new_n561_), .A3(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT97), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  XOR2_X1   g365(.A(new_n563_), .B(KEYINPUT95), .Z(new_n567_));
  NOR2_X1   g366(.A1(new_n522_), .A2(new_n448_), .ZN(new_n568_));
  OAI21_X1  g367(.A(KEYINPUT20), .B1(new_n518_), .B2(new_n559_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n567_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n560_), .A2(new_n561_), .A3(KEYINPUT97), .A4(new_n563_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n544_), .B1(new_n566_), .B2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n564_), .A2(new_n565_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n574_), .A2(new_n570_), .A3(new_n571_), .A4(new_n543_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n573_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT27), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n548_), .A2(new_n555_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n556_), .A2(new_n558_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n545_), .B1(new_n522_), .B2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n567_), .ZN(new_n582_));
  OAI211_X1 g381(.A(new_n581_), .B(new_n582_), .C1(new_n448_), .C2(new_n522_), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n560_), .A2(new_n561_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n583_), .B1(new_n584_), .B2(new_n563_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n577_), .B1(new_n585_), .B2(new_n544_), .ZN(new_n586_));
  AOI22_X1  g385(.A1(new_n576_), .A2(new_n577_), .B1(new_n575_), .B2(new_n586_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n480_), .A2(KEYINPUT105), .A3(new_n538_), .A4(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT105), .ZN(new_n589_));
  INV_X1    g388(.A(new_n529_), .ZN(new_n590_));
  AOI21_X1  g389(.A(KEYINPUT94), .B1(new_n533_), .B2(new_n489_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n537_), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n587_), .B(new_n590_), .C1(new_n591_), .C2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n418_), .A2(new_n472_), .A3(new_n479_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n589_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n588_), .A2(new_n595_), .ZN(new_n596_));
  NOR3_X1   g395(.A1(new_n568_), .A2(new_n569_), .A3(new_n567_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n563_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n598_));
  OAI211_X1 g397(.A(KEYINPUT32), .B(new_n543_), .C1(new_n597_), .C2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n543_), .A2(KEYINPUT32), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n574_), .A2(new_n570_), .A3(new_n571_), .A4(new_n600_), .ZN(new_n601_));
  AND2_X1   g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n602_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT103), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n570_), .A2(new_n571_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n543_), .B1(new_n606_), .B2(new_n574_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n575_), .ZN(new_n608_));
  OAI21_X1  g407(.A(KEYINPUT99), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT99), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n573_), .A2(new_n610_), .A3(new_n575_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n408_), .B1(new_n410_), .B2(new_n333_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n397_), .A2(new_n399_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n394_), .A2(new_n332_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n612_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(KEYINPUT101), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT101), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n617_), .B(new_n612_), .C1(new_n613_), .C2(new_n614_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n473_), .A2(KEYINPUT33), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT33), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n400_), .A2(new_n621_), .A3(new_n404_), .A4(new_n408_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n609_), .A2(new_n611_), .A3(new_n619_), .A4(new_n623_), .ZN(new_n624_));
  OAI211_X1 g423(.A(KEYINPUT103), .B(new_n602_), .C1(new_n416_), .C2(new_n417_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n605_), .A2(new_n624_), .A3(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(new_n538_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n418_), .A2(new_n479_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n590_), .B1(new_n592_), .B2(new_n591_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n629_), .A2(new_n630_), .A3(new_n587_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n472_), .B1(new_n627_), .B2(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n596_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n236_), .A2(new_n316_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(G229gat), .A2(G233gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT77), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n634_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n251_), .ZN(new_n638_));
  AOI21_X1  g437(.A(KEYINPUT15), .B1(new_n231_), .B2(new_n234_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n317_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT76), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n252_), .A2(KEYINPUT76), .A3(new_n317_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n637_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n317_), .A2(new_n235_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n635_), .B1(new_n634_), .B2(new_n645_), .ZN(new_n646_));
  NOR3_X1   g445(.A1(new_n644_), .A2(KEYINPUT80), .A3(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT80), .ZN(new_n648_));
  INV_X1    g447(.A(new_n637_), .ZN(new_n649_));
  AOI21_X1  g448(.A(KEYINPUT76), .B1(new_n252_), .B2(new_n317_), .ZN(new_n650_));
  AOI211_X1 g449(.A(new_n641_), .B(new_n316_), .C1(new_n250_), .C2(new_n251_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n649_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n646_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n648_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(G113gat), .B(G141gat), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT79), .ZN(new_n656_));
  XOR2_X1   g455(.A(G169gat), .B(G197gat), .Z(new_n657_));
  XNOR2_X1  g456(.A(new_n656_), .B(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  OAI22_X1  g458(.A1(new_n647_), .A2(new_n654_), .B1(KEYINPUT78), .B2(new_n659_), .ZN(new_n660_));
  OAI21_X1  g459(.A(KEYINPUT80), .B1(new_n644_), .B2(new_n646_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n652_), .A2(new_n653_), .A3(new_n648_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n659_), .A2(KEYINPUT78), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n661_), .A2(new_n662_), .A3(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n660_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n633_), .A2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n331_), .A2(new_n667_), .ZN(new_n668_));
  NOR3_X1   g467(.A1(new_n668_), .A2(G1gat), .A3(new_n629_), .ZN(new_n669_));
  OR2_X1    g468(.A1(new_n669_), .A2(KEYINPUT38), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(KEYINPUT38), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n633_), .A2(new_n265_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n672_), .A2(new_n665_), .A3(new_n306_), .A4(new_n329_), .ZN(new_n673_));
  OAI21_X1  g472(.A(G1gat), .B1(new_n673_), .B2(new_n629_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n670_), .A2(new_n671_), .A3(new_n674_), .ZN(G1324gat));
  OAI21_X1  g474(.A(G8gat), .B1(new_n673_), .B2(new_n587_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT39), .ZN(new_n677_));
  INV_X1    g476(.A(new_n668_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n587_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n678_), .A2(new_n312_), .A3(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n677_), .A2(new_n680_), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n681_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g481(.A(new_n472_), .ZN(new_n683_));
  OAI21_X1  g482(.A(G15gat), .B1(new_n673_), .B2(new_n683_), .ZN(new_n684_));
  XOR2_X1   g483(.A(new_n684_), .B(KEYINPUT41), .Z(new_n685_));
  NAND3_X1  g484(.A1(new_n678_), .A2(new_n454_), .A3(new_n472_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(G1326gat));
  OAI21_X1  g486(.A(G22gat), .B1(new_n673_), .B2(new_n538_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT42), .ZN(new_n689_));
  OR2_X1    g488(.A1(new_n538_), .A2(G22gat), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n689_), .B1(new_n668_), .B2(new_n690_), .ZN(G1327gat));
  INV_X1    g490(.A(new_n306_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n692_), .A2(new_n329_), .A3(new_n666_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n588_), .A2(new_n595_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n587_), .A2(new_n418_), .A3(new_n479_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n697_), .A2(new_n538_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n698_), .B1(new_n538_), .B2(new_n626_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n696_), .B1(new_n699_), .B2(new_n472_), .ZN(new_n700_));
  AOI211_X1 g499(.A(new_n694_), .B(new_n695_), .C1(new_n700_), .C2(new_n266_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n266_), .B1(new_n596_), .B2(new_n632_), .ZN(new_n702_));
  AOI21_X1  g501(.A(KEYINPUT43), .B1(new_n702_), .B2(KEYINPUT106), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n693_), .B1(new_n701_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  OAI211_X1 g505(.A(KEYINPUT44), .B(new_n693_), .C1(new_n701_), .C2(new_n703_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(G29gat), .B1(new_n708_), .B2(new_n629_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n328_), .A2(new_n265_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT107), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n667_), .A2(new_n711_), .A3(new_n306_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n629_), .A2(G29gat), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n713_), .B(KEYINPUT108), .Z(new_n714_));
  OAI21_X1  g513(.A(new_n709_), .B1(new_n712_), .B2(new_n714_), .ZN(G1328gat));
  NOR3_X1   g514(.A1(new_n712_), .A2(G36gat), .A3(new_n587_), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT45), .Z(new_n717_));
  NAND3_X1  g516(.A1(new_n706_), .A2(new_n679_), .A3(new_n707_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT109), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n718_), .A2(new_n719_), .A3(G36gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(new_n718_), .B2(G36gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n717_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT46), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  OAI211_X1 g523(.A(new_n717_), .B(KEYINPUT46), .C1(new_n720_), .C2(new_n721_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(G1329gat));
  NAND2_X1  g525(.A1(new_n472_), .A2(G43gat), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n712_), .A2(new_n683_), .ZN(new_n728_));
  OAI22_X1  g527(.A1(new_n708_), .A2(new_n727_), .B1(G43gat), .B2(new_n728_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g529(.A(new_n712_), .ZN(new_n731_));
  AOI21_X1  g530(.A(G50gat), .B1(new_n731_), .B2(new_n630_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n708_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n630_), .A2(G50gat), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n732_), .B1(new_n733_), .B2(new_n734_), .ZN(G1331gat));
  NAND4_X1  g534(.A1(new_n672_), .A2(new_n666_), .A3(new_n692_), .A4(new_n329_), .ZN(new_n736_));
  OAI21_X1  g535(.A(G57gat), .B1(new_n736_), .B2(new_n629_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n633_), .A2(new_n665_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n266_), .A2(new_n328_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n738_), .A2(new_n692_), .A3(new_n739_), .ZN(new_n740_));
  OR2_X1    g539(.A1(new_n629_), .A2(G57gat), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n737_), .B1(new_n740_), .B2(new_n741_), .ZN(G1332gat));
  OAI21_X1  g541(.A(G64gat), .B1(new_n736_), .B2(new_n587_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT48), .ZN(new_n744_));
  OR2_X1    g543(.A1(new_n587_), .A2(G64gat), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n744_), .B1(new_n740_), .B2(new_n745_), .ZN(G1333gat));
  OAI21_X1  g545(.A(G71gat), .B1(new_n736_), .B2(new_n683_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT49), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n683_), .A2(G71gat), .ZN(new_n749_));
  XOR2_X1   g548(.A(new_n749_), .B(KEYINPUT110), .Z(new_n750_));
  OAI21_X1  g549(.A(new_n748_), .B1(new_n740_), .B2(new_n750_), .ZN(G1334gat));
  OAI21_X1  g550(.A(G78gat), .B1(new_n736_), .B2(new_n538_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n752_), .B(new_n753_), .ZN(new_n754_));
  OR2_X1    g553(.A1(new_n538_), .A2(G78gat), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n754_), .B1(new_n740_), .B2(new_n755_), .ZN(G1335gat));
  NAND3_X1  g555(.A1(new_n738_), .A2(new_n711_), .A3(new_n692_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(G85gat), .B1(new_n758_), .B2(new_n628_), .ZN(new_n759_));
  OR2_X1    g558(.A1(new_n701_), .A2(new_n703_), .ZN(new_n760_));
  NOR3_X1   g559(.A1(new_n306_), .A2(new_n665_), .A3(new_n329_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n628_), .A2(new_n209_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n759_), .B1(new_n763_), .B2(new_n764_), .ZN(G1336gat));
  AOI21_X1  g564(.A(G92gat), .B1(new_n758_), .B2(new_n679_), .ZN(new_n766_));
  XOR2_X1   g565(.A(new_n766_), .B(KEYINPUT112), .Z(new_n767_));
  NAND2_X1  g566(.A1(new_n679_), .A2(G92gat), .ZN(new_n768_));
  XOR2_X1   g567(.A(new_n768_), .B(KEYINPUT113), .Z(new_n769_));
  AOI21_X1  g568(.A(new_n767_), .B1(new_n763_), .B2(new_n769_), .ZN(G1337gat));
  NAND3_X1  g569(.A1(new_n758_), .A2(new_n472_), .A3(new_n214_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n760_), .A2(new_n472_), .A3(new_n761_), .ZN(new_n772_));
  AND3_X1   g571(.A1(new_n772_), .A2(KEYINPUT114), .A3(G99gat), .ZN(new_n773_));
  AOI21_X1  g572(.A(KEYINPUT114), .B1(new_n772_), .B2(G99gat), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n771_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g575(.A1(new_n758_), .A2(new_n215_), .A3(new_n630_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT115), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n760_), .A2(new_n630_), .A3(new_n761_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(KEYINPUT116), .B(KEYINPUT52), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n779_), .A2(G106gat), .A3(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n781_), .B1(new_n779_), .B2(G106gat), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n778_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g584(.A1(new_n593_), .A2(new_n629_), .A3(new_n683_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n788_));
  INV_X1    g587(.A(new_n281_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n289_), .A2(new_n292_), .A3(new_n294_), .A4(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(new_n269_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n296_), .A2(new_n792_), .ZN(new_n793_));
  AOI22_X1  g592(.A1(new_n288_), .A2(KEYINPUT70), .B1(new_n290_), .B2(new_n291_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n794_), .A2(KEYINPUT55), .A3(new_n294_), .A4(new_n295_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n791_), .A2(new_n793_), .A3(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(new_n301_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT56), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n796_), .A2(KEYINPUT56), .A3(new_n301_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT117), .ZN(new_n802_));
  INV_X1    g601(.A(new_n664_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n663_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n304_), .B(new_n802_), .C1(new_n803_), .C2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n802_), .B1(new_n665_), .B2(new_n304_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n636_), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n634_), .B(new_n809_), .C1(new_n650_), .C2(new_n651_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n634_), .A2(new_n645_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n659_), .B1(new_n811_), .B2(new_n636_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n812_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n813_), .B(KEYINPUT118), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n644_), .A2(new_n658_), .A3(new_n646_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  AOI22_X1  g615(.A1(new_n801_), .A2(new_n808_), .B1(new_n305_), .B2(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n788_), .B1(new_n817_), .B2(new_n265_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n305_), .A2(new_n816_), .ZN(new_n819_));
  AND3_X1   g618(.A1(new_n796_), .A2(KEYINPUT56), .A3(new_n301_), .ZN(new_n820_));
  AOI21_X1  g619(.A(KEYINPUT56), .B1(new_n796_), .B2(new_n301_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n665_), .A2(new_n304_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT117), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n805_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n819_), .B1(new_n822_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n265_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(KEYINPUT57), .A3(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT58), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n816_), .A2(new_n304_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n829_), .B1(new_n822_), .B2(new_n830_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n801_), .A2(KEYINPUT58), .A3(new_n304_), .A4(new_n816_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n831_), .A2(new_n832_), .A3(new_n266_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n818_), .A2(new_n828_), .A3(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n328_), .ZN(new_n835_));
  OAI21_X1  g634(.A(KEYINPUT54), .B1(new_n330_), .B2(new_n665_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT54), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n739_), .A2(new_n837_), .A3(new_n666_), .A4(new_n306_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n787_), .B1(new_n835_), .B2(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(G113gat), .B1(new_n840_), .B2(new_n665_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT120), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n841_), .B(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT59), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n840_), .A2(KEYINPUT121), .A3(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(KEYINPUT121), .B1(new_n840_), .B2(new_n844_), .ZN(new_n847_));
  OAI22_X1  g646(.A1(new_n846_), .A2(new_n847_), .B1(new_n844_), .B2(new_n840_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n665_), .A2(G113gat), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n843_), .B1(new_n849_), .B2(new_n850_), .ZN(G1340gat));
  NAND2_X1  g650(.A1(new_n835_), .A2(new_n839_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n786_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT60), .ZN(new_n854_));
  AND2_X1   g653(.A1(new_n854_), .A2(G120gat), .ZN(new_n855_));
  AOI21_X1  g654(.A(G120gat), .B1(new_n692_), .B2(new_n854_), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n853_), .A2(new_n855_), .A3(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT122), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n857_), .B(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n692_), .B1(new_n840_), .B2(new_n844_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n852_), .A2(new_n844_), .A3(new_n786_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT121), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n860_), .B1(new_n863_), .B2(new_n845_), .ZN(new_n864_));
  OAI21_X1  g663(.A(G120gat), .B1(new_n864_), .B2(KEYINPUT123), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n306_), .B1(new_n853_), .B2(KEYINPUT59), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n866_), .B(KEYINPUT123), .C1(new_n846_), .C2(new_n847_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n859_), .B1(new_n865_), .B2(new_n868_), .ZN(G1341gat));
  OAI21_X1  g668(.A(G127gat), .B1(new_n848_), .B2(new_n328_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n840_), .A2(new_n372_), .A3(new_n329_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(G1342gat));
  OAI21_X1  g671(.A(G134gat), .B1(new_n848_), .B2(new_n267_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n840_), .A2(new_n370_), .A3(new_n265_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(G1343gat));
  AOI21_X1  g674(.A(new_n538_), .B1(new_n835_), .B2(new_n839_), .ZN(new_n876_));
  NOR3_X1   g675(.A1(new_n629_), .A2(new_n472_), .A3(new_n679_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n665_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n692_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g682(.A1(new_n878_), .A2(new_n328_), .ZN(new_n884_));
  XOR2_X1   g683(.A(KEYINPUT61), .B(G155gat), .Z(new_n885_));
  XNOR2_X1  g684(.A(new_n884_), .B(new_n885_), .ZN(G1346gat));
  OR3_X1    g685(.A1(new_n878_), .A2(G162gat), .A3(new_n827_), .ZN(new_n887_));
  OAI21_X1  g686(.A(G162gat), .B1(new_n878_), .B2(new_n267_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(G1347gat));
  INV_X1    g688(.A(KEYINPUT124), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n594_), .A2(new_n630_), .A3(new_n587_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n852_), .A2(new_n891_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n892_), .A2(new_n666_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(new_n426_), .ZN(new_n894_));
  OAI211_X1 g693(.A(KEYINPUT62), .B(G169gat), .C1(new_n892_), .C2(new_n666_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  AND2_X1   g695(.A1(new_n852_), .A2(new_n891_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n665_), .ZN(new_n898_));
  AOI21_X1  g697(.A(KEYINPUT62), .B1(new_n898_), .B2(G169gat), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n890_), .B1(new_n896_), .B2(new_n899_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT62), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n901_), .B1(new_n893_), .B2(new_n432_), .ZN(new_n902_));
  NAND4_X1  g701(.A1(new_n902_), .A2(KEYINPUT124), .A3(new_n894_), .A4(new_n895_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n900_), .A2(new_n903_), .ZN(G1348gat));
  AOI21_X1  g703(.A(new_n306_), .B1(KEYINPUT125), .B2(new_n427_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n897_), .A2(new_n905_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n427_), .A2(KEYINPUT125), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n906_), .B(new_n907_), .ZN(G1349gat));
  NAND2_X1  g707(.A1(new_n897_), .A2(new_n329_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n553_), .A2(new_n554_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  OR3_X1    g710(.A1(new_n909_), .A2(KEYINPUT126), .A3(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(KEYINPUT126), .B1(new_n909_), .B2(new_n911_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n909_), .A2(new_n550_), .ZN(new_n914_));
  AND3_X1   g713(.A1(new_n912_), .A2(new_n913_), .A3(new_n914_), .ZN(G1350gat));
  OAI21_X1  g714(.A(G190gat), .B1(new_n892_), .B2(new_n267_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n265_), .A2(new_n439_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(KEYINPUT127), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n916_), .B1(new_n892_), .B2(new_n918_), .ZN(G1351gat));
  NOR3_X1   g718(.A1(new_n628_), .A2(new_n472_), .A3(new_n587_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n876_), .A2(new_n920_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n921_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(new_n665_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g723(.A1(new_n922_), .A2(new_n692_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g725(.A1(new_n921_), .A2(new_n328_), .ZN(new_n927_));
  NOR3_X1   g726(.A1(new_n927_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n928_));
  XOR2_X1   g727(.A(KEYINPUT63), .B(G211gat), .Z(new_n929_));
  AOI21_X1  g728(.A(new_n928_), .B1(new_n927_), .B2(new_n929_), .ZN(G1354gat));
  OAI21_X1  g729(.A(G218gat), .B1(new_n921_), .B2(new_n267_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n265_), .A2(new_n498_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n931_), .B1(new_n921_), .B2(new_n932_), .ZN(G1355gat));
endmodule


