//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 1 1 0 1 0 1 0 0 0 1 0 0 1 1 1 0 0 0 0 1 1 0 0 0 1 0 1 1 1 1 1 1 0 0 1 1 1 1 1 0 1 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n705_, new_n706_,
    new_n707_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n722_, new_n723_, new_n724_, new_n725_, new_n727_,
    new_n728_, new_n729_, new_n731_, new_n732_, new_n733_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n742_,
    new_n743_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n833_, new_n834_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n843_, new_n844_, new_n845_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n877_, new_n879_, new_n880_, new_n881_, new_n882_,
    new_n884_, new_n886_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_, new_n896_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  INV_X1    g001(.A(G43gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G50gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT15), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n204_), .B(G50gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT15), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n207_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT6), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n214_));
  OR3_X1    g013(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n213_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  XOR2_X1   g015(.A(G85gat), .B(G92gat), .Z(new_n217_));
  INV_X1    g016(.A(KEYINPUT64), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT8), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n216_), .A2(new_n217_), .A3(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n218_), .A2(KEYINPUT8), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  XOR2_X1   g021(.A(KEYINPUT10), .B(G99gat), .Z(new_n223_));
  INV_X1    g022(.A(G106gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n217_), .A2(KEYINPUT9), .ZN(new_n226_));
  INV_X1    g025(.A(G85gat), .ZN(new_n227_));
  INV_X1    g026(.A(G92gat), .ZN(new_n228_));
  OR3_X1    g027(.A1(new_n227_), .A2(new_n228_), .A3(KEYINPUT9), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n225_), .A2(new_n226_), .A3(new_n229_), .A4(new_n213_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n221_), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n216_), .A2(new_n217_), .A3(new_n231_), .A4(new_n219_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n222_), .A2(new_n230_), .A3(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n211_), .A2(new_n233_), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n233_), .A2(new_n208_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G232gat), .A2(G233gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT34), .ZN(new_n237_));
  XOR2_X1   g036(.A(new_n237_), .B(KEYINPUT35), .Z(new_n238_));
  NAND3_X1  g037(.A1(new_n234_), .A2(new_n235_), .A3(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT70), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n234_), .A2(new_n235_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n242_), .A2(KEYINPUT35), .A3(new_n237_), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n234_), .A2(KEYINPUT70), .A3(new_n235_), .A4(new_n238_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n241_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT69), .B(G190gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(G218gat), .ZN(new_n247_));
  XOR2_X1   g046(.A(G134gat), .B(G162gat), .Z(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT36), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n249_), .A2(new_n250_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n245_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n251_), .B1(new_n245_), .B2(new_n252_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT101), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G57gat), .B(G64gat), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n258_), .A2(KEYINPUT11), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(KEYINPUT11), .ZN(new_n260_));
  XOR2_X1   g059(.A(G71gat), .B(G78gat), .Z(new_n261_));
  NAND3_X1  g060(.A1(new_n259_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n262_));
  OR2_X1    g061(.A1(new_n260_), .A2(new_n261_), .ZN(new_n263_));
  AND2_X1   g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n233_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(KEYINPUT65), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(KEYINPUT12), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G230gat), .A2(G233gat), .ZN(new_n268_));
  OR2_X1    g067(.A1(new_n233_), .A2(new_n264_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT65), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n270_), .B1(new_n233_), .B2(new_n264_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT12), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n267_), .A2(new_n268_), .A3(new_n269_), .A4(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n269_), .A2(new_n265_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n275_), .A2(G230gat), .A3(G233gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n274_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT66), .ZN(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT67), .B(G204gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G120gat), .B(G148gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT5), .B(G176gat), .ZN(new_n282_));
  XOR2_X1   g081(.A(new_n281_), .B(new_n282_), .Z(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT68), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT66), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n274_), .A2(new_n286_), .A3(new_n276_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n278_), .A2(new_n285_), .A3(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT13), .ZN(new_n289_));
  INV_X1    g088(.A(new_n283_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n274_), .A2(new_n276_), .A3(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n288_), .A2(new_n289_), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n289_), .B1(new_n288_), .B2(new_n291_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT71), .B(G22gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(G15gat), .ZN(new_n297_));
  INV_X1    g096(.A(G1gat), .ZN(new_n298_));
  INV_X1    g097(.A(G8gat), .ZN(new_n299_));
  OAI21_X1  g098(.A(KEYINPUT14), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n297_), .A2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT72), .B(KEYINPUT73), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G1gat), .B(G8gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n301_), .B(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(new_n206_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G229gat), .A2(G233gat), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n305_), .A2(new_n206_), .ZN(new_n310_));
  AND2_X1   g109(.A1(new_n207_), .A2(new_n210_), .ZN(new_n311_));
  OAI211_X1 g110(.A(new_n307_), .B(new_n310_), .C1(new_n311_), .C2(new_n305_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n309_), .A2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G113gat), .B(G141gat), .ZN(new_n314_));
  INV_X1    g113(.A(G169gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(G197gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n313_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n318_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n309_), .A2(new_n312_), .A3(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G231gat), .A2(G233gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n264_), .B(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(new_n305_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G127gat), .B(G155gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G183gat), .B(G211gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT17), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n331_), .A2(new_n332_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n326_), .A2(new_n333_), .A3(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT76), .ZN(new_n337_));
  OR2_X1    g136(.A1(new_n326_), .A2(KEYINPUT74), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n326_), .A2(KEYINPUT74), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n338_), .A2(new_n334_), .A3(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n337_), .A2(new_n340_), .ZN(new_n341_));
  NOR3_X1   g140(.A1(new_n295_), .A2(new_n323_), .A3(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT100), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n257_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G225gat), .A2(G233gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT81), .B(G127gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(G134gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G113gat), .B(G120gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  XOR2_X1   g148(.A(G155gat), .B(G162gat), .Z(new_n350_));
  INV_X1    g149(.A(KEYINPUT1), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(G141gat), .ZN(new_n353_));
  INV_X1    g152(.A(G148gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G141gat), .A2(G148gat), .ZN(new_n356_));
  NAND3_X1  g155(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n352_), .A2(new_n355_), .A3(new_n356_), .A4(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(KEYINPUT84), .A2(KEYINPUT2), .ZN(new_n359_));
  NOR2_X1   g158(.A1(KEYINPUT84), .A2(KEYINPUT2), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n359_), .B1(new_n360_), .B2(new_n356_), .ZN(new_n361_));
  OAI21_X1  g160(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT3), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n363_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(KEYINPUT84), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n361_), .A2(new_n362_), .A3(new_n364_), .A4(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT85), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n366_), .A2(new_n367_), .A3(new_n350_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n367_), .B1(new_n366_), .B2(new_n350_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n358_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  OR2_X1    g169(.A1(new_n349_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n349_), .A2(new_n370_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n371_), .A2(KEYINPUT4), .A3(new_n372_), .ZN(new_n373_));
  OR2_X1    g172(.A1(new_n372_), .A2(KEYINPUT4), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n345_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT0), .B(G57gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(G85gat), .ZN(new_n378_));
  XOR2_X1   g177(.A(G1gat), .B(G29gat), .Z(new_n379_));
  XOR2_X1   g178(.A(new_n378_), .B(new_n379_), .Z(new_n380_));
  NAND2_X1  g179(.A1(new_n371_), .A2(new_n372_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(new_n345_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n376_), .A2(new_n380_), .A3(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n380_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n382_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n384_), .B1(new_n385_), .B2(new_n375_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n383_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT27), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G226gat), .A2(G233gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT19), .ZN(new_n391_));
  AND2_X1   g190(.A1(KEYINPUT87), .A2(G197gat), .ZN(new_n392_));
  NOR2_X1   g191(.A1(KEYINPUT87), .A2(G197gat), .ZN(new_n393_));
  OAI21_X1  g192(.A(G204gat), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n317_), .A2(G204gat), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n394_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT21), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G211gat), .B(G218gat), .ZN(new_n399_));
  NOR3_X1   g198(.A1(new_n397_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n394_), .A2(new_n398_), .A3(new_n396_), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n402_), .A2(new_n399_), .ZN(new_n403_));
  NOR3_X1   g202(.A1(new_n392_), .A2(new_n393_), .A3(G204gat), .ZN(new_n404_));
  INV_X1    g203(.A(G204gat), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT88), .B1(new_n405_), .B2(G197gat), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT88), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n407_), .A2(new_n317_), .A3(G204gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n406_), .A2(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT21), .B1(new_n404_), .B2(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(KEYINPUT89), .B1(new_n403_), .B2(new_n410_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n410_), .A2(KEYINPUT89), .A3(new_n399_), .A4(new_n402_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n401_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(KEYINPUT26), .B(G190gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(KEYINPUT25), .B(G183gat), .ZN(new_n416_));
  AND2_X1   g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  OR2_X1    g216(.A1(G169gat), .A2(G176gat), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n418_), .A2(KEYINPUT24), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G169gat), .A2(G176gat), .ZN(new_n420_));
  AND3_X1   g219(.A1(new_n418_), .A2(KEYINPUT24), .A3(new_n420_), .ZN(new_n421_));
  NOR3_X1   g220(.A1(new_n417_), .A2(new_n419_), .A3(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT23), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n423_), .A2(G183gat), .A3(G190gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(KEYINPUT77), .ZN(new_n425_));
  INV_X1    g224(.A(G183gat), .ZN(new_n426_));
  INV_X1    g225(.A(G190gat), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT23), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT77), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n429_), .A2(new_n423_), .A3(G183gat), .A4(G190gat), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n425_), .A2(new_n428_), .A3(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n422_), .A2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(KEYINPUT78), .B(G169gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT22), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT79), .ZN(new_n435_));
  XOR2_X1   g234(.A(KEYINPUT80), .B(G176gat), .Z(new_n436_));
  INV_X1    g235(.A(KEYINPUT22), .ZN(new_n437_));
  AOI21_X1  g236(.A(KEYINPUT79), .B1(new_n437_), .B2(new_n315_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n438_), .B1(new_n433_), .B2(new_n437_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n435_), .A2(new_n436_), .A3(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n428_), .A2(new_n424_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n426_), .A2(new_n427_), .ZN(new_n442_));
  AOI22_X1  g241(.A1(new_n441_), .A2(new_n442_), .B1(G169gat), .B2(G176gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n440_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n432_), .A2(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT20), .B1(new_n414_), .B2(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n416_), .B(KEYINPUT91), .ZN(new_n447_));
  AOI22_X1  g246(.A1(new_n447_), .A2(new_n415_), .B1(new_n428_), .B2(new_n424_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n420_), .A2(KEYINPUT24), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(KEYINPUT92), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n419_), .B1(new_n450_), .B2(new_n418_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(KEYINPUT22), .B(G169gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n436_), .A2(new_n452_), .ZN(new_n453_));
  AOI22_X1  g252(.A1(new_n431_), .A2(new_n442_), .B1(G169gat), .B2(G176gat), .ZN(new_n454_));
  AOI22_X1  g253(.A1(new_n448_), .A2(new_n451_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT89), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n402_), .A2(new_n399_), .ZN(new_n457_));
  AND2_X1   g256(.A1(new_n406_), .A2(new_n408_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n393_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(KEYINPUT87), .A2(G197gat), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n459_), .A2(new_n405_), .A3(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n398_), .B1(new_n458_), .B2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n456_), .B1(new_n457_), .B2(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n400_), .B1(new_n463_), .B2(new_n412_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n455_), .A2(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n391_), .B1(new_n446_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT93), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n414_), .A2(new_n467_), .A3(new_n445_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT20), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n469_), .B1(new_n455_), .B2(new_n464_), .ZN(new_n470_));
  AOI22_X1  g269(.A1(new_n431_), .A2(new_n422_), .B1(new_n440_), .B2(new_n443_), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT93), .B1(new_n464_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n391_), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n468_), .A2(new_n470_), .A3(new_n472_), .A4(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT18), .B(G64gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(G92gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G8gat), .B(G36gat), .ZN(new_n477_));
  XOR2_X1   g276(.A(new_n476_), .B(new_n477_), .Z(new_n478_));
  NAND3_X1  g277(.A1(new_n466_), .A2(new_n474_), .A3(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(KEYINPUT99), .ZN(new_n480_));
  NOR3_X1   g279(.A1(new_n446_), .A2(new_n391_), .A3(new_n465_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT97), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT97), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n468_), .A2(new_n470_), .A3(new_n472_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n483_), .B1(new_n484_), .B2(new_n391_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n482_), .B1(new_n485_), .B2(new_n481_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n478_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n389_), .B1(new_n480_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n479_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n478_), .B1(new_n466_), .B2(new_n474_), .ZN(new_n491_));
  NOR3_X1   g290(.A1(new_n490_), .A2(KEYINPUT27), .A3(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n489_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G228gat), .A2(G233gat), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT29), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n366_), .A2(new_n350_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT85), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n366_), .A2(new_n367_), .A3(new_n350_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n498_), .B1(new_n502_), .B2(new_n358_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G78gat), .B(G106gat), .ZN(new_n504_));
  NOR3_X1   g303(.A1(new_n503_), .A2(new_n464_), .A3(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n504_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n370_), .A2(KEYINPUT29), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n506_), .B1(new_n414_), .B2(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n497_), .B1(new_n505_), .B2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT86), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n504_), .B1(new_n503_), .B2(new_n464_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n414_), .A2(new_n507_), .A3(new_n506_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n497_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n511_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n509_), .A2(new_n510_), .A3(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n502_), .A2(new_n498_), .A3(new_n358_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G22gat), .B(G50gat), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n509_), .A2(new_n510_), .A3(new_n514_), .A4(new_n516_), .ZN(new_n521_));
  AND3_X1   g320(.A1(new_n518_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n520_), .B1(new_n518_), .B2(new_n521_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n496_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  AND3_X1   g323(.A1(new_n511_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n513_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n516_), .B1(new_n527_), .B2(new_n510_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n521_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n519_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n518_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n530_), .A2(new_n495_), .A3(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G71gat), .B(G99gat), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G227gat), .A2(G233gat), .ZN(new_n535_));
  XOR2_X1   g334(.A(new_n535_), .B(KEYINPUT30), .Z(new_n536_));
  NAND2_X1  g335(.A1(new_n471_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n471_), .A2(new_n536_), .ZN(new_n539_));
  XOR2_X1   g338(.A(G15gat), .B(G43gat), .Z(new_n540_));
  NOR3_X1   g339(.A1(new_n538_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n540_), .ZN(new_n542_));
  OR2_X1    g341(.A1(new_n471_), .A2(new_n536_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n542_), .B1(new_n543_), .B2(new_n537_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n534_), .B1(new_n541_), .B2(new_n544_), .ZN(new_n545_));
  XOR2_X1   g344(.A(new_n349_), .B(KEYINPUT31), .Z(new_n546_));
  OAI21_X1  g345(.A(new_n540_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n543_), .A2(new_n542_), .A3(new_n537_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n547_), .A2(new_n533_), .A3(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n545_), .A2(new_n546_), .A3(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT82), .ZN(new_n551_));
  AND2_X1   g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n550_), .A2(new_n551_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT83), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n545_), .A2(new_n549_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n546_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n554_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  AOI211_X1 g356(.A(KEYINPUT83), .B(new_n546_), .C1(new_n545_), .C2(new_n549_), .ZN(new_n558_));
  OAI22_X1  g357(.A1(new_n552_), .A2(new_n553_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  AND3_X1   g358(.A1(new_n524_), .A2(new_n532_), .A3(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n559_), .B1(new_n524_), .B2(new_n532_), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n388_), .B(new_n494_), .C1(new_n560_), .C2(new_n561_), .ZN(new_n562_));
  NOR3_X1   g361(.A1(new_n522_), .A2(new_n523_), .A3(new_n496_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n495_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n564_));
  NOR3_X1   g363(.A1(new_n563_), .A2(new_n564_), .A3(new_n559_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n490_), .A2(new_n491_), .ZN(new_n566_));
  OR2_X1    g365(.A1(new_n566_), .A2(KEYINPUT94), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n386_), .B(KEYINPUT33), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n566_), .A2(KEYINPUT94), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n345_), .B1(new_n381_), .B2(KEYINPUT95), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n570_), .B1(KEYINPUT95), .B2(new_n381_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n373_), .A2(new_n345_), .A3(new_n374_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n571_), .A2(new_n380_), .A3(new_n572_), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n567_), .A2(new_n568_), .A3(new_n569_), .A4(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n478_), .A2(KEYINPUT32), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  AOI22_X1  g375(.A1(new_n576_), .A2(new_n486_), .B1(new_n383_), .B2(new_n386_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n466_), .A2(new_n474_), .A3(new_n575_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT96), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n577_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT98), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n577_), .A2(KEYINPUT98), .A3(new_n580_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n574_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n565_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n562_), .A2(new_n586_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n344_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n342_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(KEYINPUT100), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT102), .ZN(new_n592_));
  OAI21_X1  g391(.A(G1gat), .B1(new_n592_), .B2(new_n388_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n559_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n594_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n524_), .A2(new_n532_), .A3(new_n559_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n493_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  AOI22_X1  g396(.A1(new_n597_), .A2(new_n388_), .B1(new_n585_), .B2(new_n565_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT37), .ZN(new_n599_));
  NOR3_X1   g398(.A1(new_n254_), .A2(new_n255_), .A3(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n245_), .A2(new_n252_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n251_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(KEYINPUT37), .B1(new_n603_), .B2(new_n253_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n600_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NOR3_X1   g405(.A1(new_n598_), .A2(new_n589_), .A3(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n607_), .A2(new_n298_), .A3(new_n387_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT38), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n593_), .A2(new_n609_), .ZN(G1324gat));
  INV_X1    g409(.A(KEYINPUT103), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n588_), .A2(new_n611_), .A3(new_n590_), .A4(new_n493_), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n590_), .A2(new_n344_), .A3(new_n493_), .A4(new_n587_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(KEYINPUT103), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n612_), .A2(G8gat), .A3(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(KEYINPUT39), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT39), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n612_), .A2(new_n614_), .A3(new_n617_), .A4(G8gat), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n607_), .A2(new_n299_), .A3(new_n493_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(KEYINPUT104), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT104), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n619_), .A2(new_n623_), .A3(new_n620_), .ZN(new_n624_));
  AND3_X1   g423(.A1(new_n622_), .A2(KEYINPUT40), .A3(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(KEYINPUT40), .B1(new_n622_), .B2(new_n624_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n625_), .A2(new_n626_), .ZN(G1325gat));
  OAI21_X1  g426(.A(G15gat), .B1(new_n592_), .B2(new_n594_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n628_), .B(KEYINPUT41), .Z(new_n629_));
  INV_X1    g428(.A(G15gat), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n607_), .A2(new_n630_), .A3(new_n559_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n629_), .A2(new_n631_), .ZN(G1326gat));
  NOR2_X1   g431(.A1(new_n563_), .A2(new_n564_), .ZN(new_n633_));
  OAI21_X1  g432(.A(G22gat), .B1(new_n592_), .B2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT42), .ZN(new_n635_));
  INV_X1    g434(.A(G22gat), .ZN(new_n636_));
  INV_X1    g435(.A(new_n633_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n607_), .A2(new_n636_), .A3(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n635_), .A2(new_n638_), .ZN(G1327gat));
  NOR2_X1   g438(.A1(new_n605_), .A2(KEYINPUT43), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n587_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT107), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT106), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n643_), .B1(new_n600_), .B2(new_n604_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n599_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n603_), .A2(KEYINPUT37), .A3(new_n253_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n645_), .A2(new_n646_), .A3(KEYINPUT106), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n644_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n587_), .A2(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n642_), .B1(new_n650_), .B2(KEYINPUT43), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n648_), .B1(new_n562_), .B2(new_n586_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT43), .ZN(new_n653_));
  NOR3_X1   g452(.A1(new_n652_), .A2(KEYINPUT107), .A3(new_n653_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n641_), .B1(new_n651_), .B2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n341_), .ZN(new_n656_));
  NOR3_X1   g455(.A1(new_n295_), .A2(new_n323_), .A3(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT105), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n655_), .A2(KEYINPUT44), .A3(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT44), .ZN(new_n660_));
  INV_X1    g459(.A(new_n641_), .ZN(new_n661_));
  OAI211_X1 g460(.A(new_n642_), .B(KEYINPUT43), .C1(new_n598_), .C2(new_n648_), .ZN(new_n662_));
  OAI21_X1  g461(.A(KEYINPUT107), .B1(new_n652_), .B2(new_n653_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n661_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n658_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n660_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n659_), .A2(new_n666_), .A3(new_n387_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT108), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND4_X1  g468(.A1(new_n659_), .A2(new_n666_), .A3(KEYINPUT108), .A4(new_n387_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n669_), .A2(G29gat), .A3(new_n670_), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n587_), .A2(new_n256_), .A3(new_n657_), .ZN(new_n672_));
  INV_X1    g471(.A(G29gat), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n672_), .A2(new_n673_), .A3(new_n387_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n671_), .A2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(KEYINPUT109), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT109), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n671_), .A2(new_n677_), .A3(new_n674_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n678_), .ZN(G1328gat));
  INV_X1    g478(.A(KEYINPUT111), .ZN(new_n680_));
  INV_X1    g479(.A(G36gat), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n493_), .B(KEYINPUT110), .Z(new_n682_));
  NAND4_X1  g481(.A1(new_n672_), .A2(new_n680_), .A3(new_n681_), .A4(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n256_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n684_), .B1(new_n562_), .B2(new_n586_), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n685_), .A2(new_n681_), .A3(new_n657_), .A4(new_n682_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(KEYINPUT111), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n683_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT45), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n683_), .A2(KEYINPUT45), .A3(new_n687_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n659_), .A2(new_n666_), .A3(new_n493_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n692_), .B1(new_n693_), .B2(G36gat), .ZN(new_n694_));
  OAI21_X1  g493(.A(KEYINPUT46), .B1(new_n694_), .B2(KEYINPUT113), .ZN(new_n695_));
  OAI21_X1  g494(.A(KEYINPUT113), .B1(new_n694_), .B2(KEYINPUT112), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  OAI211_X1 g496(.A(KEYINPUT113), .B(KEYINPUT46), .C1(new_n694_), .C2(KEYINPUT112), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(G1329gat));
  AND2_X1   g498(.A1(new_n659_), .A2(new_n666_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n594_), .A2(new_n203_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n672_), .A2(new_n559_), .ZN(new_n702_));
  AOI22_X1  g501(.A1(new_n700_), .A2(new_n701_), .B1(new_n203_), .B2(new_n702_), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g503(.A(G50gat), .B1(new_n672_), .B2(new_n637_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n633_), .A2(new_n205_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n705_), .B1(new_n700_), .B2(new_n706_), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT114), .Z(G1331gat));
  INV_X1    g507(.A(new_n294_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(new_n292_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n337_), .A2(new_n323_), .A3(new_n340_), .ZN(new_n711_));
  AOI211_X1 g510(.A(new_n710_), .B(new_n711_), .C1(new_n562_), .C2(new_n586_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(new_n605_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(G57gat), .B1(new_n714_), .B2(new_n387_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n257_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n712_), .A2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT115), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n717_), .B(new_n718_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n719_), .A2(new_n388_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n715_), .B1(new_n720_), .B2(G57gat), .ZN(G1332gat));
  INV_X1    g520(.A(new_n682_), .ZN(new_n722_));
  OAI21_X1  g521(.A(G64gat), .B1(new_n719_), .B2(new_n722_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT48), .ZN(new_n724_));
  OR2_X1    g523(.A1(new_n722_), .A2(G64gat), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n724_), .B1(new_n713_), .B2(new_n725_), .ZN(G1333gat));
  OAI21_X1  g525(.A(G71gat), .B1(new_n719_), .B2(new_n594_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT49), .ZN(new_n728_));
  OR2_X1    g527(.A1(new_n594_), .A2(G71gat), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n728_), .B1(new_n713_), .B2(new_n729_), .ZN(G1334gat));
  OAI21_X1  g529(.A(G78gat), .B1(new_n719_), .B2(new_n633_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT50), .ZN(new_n732_));
  OR2_X1    g531(.A1(new_n633_), .A2(G78gat), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n713_), .B2(new_n733_), .ZN(G1335gat));
  NAND3_X1  g533(.A1(new_n295_), .A2(new_n323_), .A3(new_n341_), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n598_), .A2(new_n684_), .A3(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(G85gat), .B1(new_n736_), .B2(new_n387_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT116), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n664_), .A2(new_n735_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n388_), .A2(new_n227_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n738_), .B1(new_n739_), .B2(new_n740_), .ZN(G1336gat));
  AOI21_X1  g540(.A(G92gat), .B1(new_n736_), .B2(new_n493_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n722_), .A2(new_n228_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n739_), .B2(new_n743_), .ZN(G1337gat));
  NAND2_X1  g543(.A1(new_n739_), .A2(new_n559_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n559_), .A2(new_n223_), .ZN(new_n746_));
  AOI22_X1  g545(.A1(new_n745_), .A2(G99gat), .B1(new_n736_), .B2(new_n746_), .ZN(new_n747_));
  XOR2_X1   g546(.A(new_n747_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g547(.A1(new_n736_), .A2(new_n224_), .A3(new_n637_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT52), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n739_), .A2(new_n637_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(new_n751_), .B2(G106gat), .ZN(new_n752_));
  AOI211_X1 g551(.A(KEYINPUT52), .B(new_n224_), .C1(new_n739_), .C2(new_n637_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n749_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g554(.A1(new_n493_), .A2(new_n388_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT119), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n758_), .B(new_n310_), .C1(new_n311_), .C2(new_n305_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n305_), .B1(new_n207_), .B2(new_n210_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n305_), .A2(new_n206_), .ZN(new_n761_));
  OAI21_X1  g560(.A(KEYINPUT119), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n759_), .A2(new_n762_), .A3(new_n308_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n306_), .A2(new_n307_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n763_), .A2(new_n318_), .A3(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n765_), .A2(new_n321_), .A3(new_n291_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT122), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n766_), .B(new_n767_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n271_), .B(KEYINPUT12), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n268_), .B1(new_n769_), .B2(new_n269_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT55), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n274_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n769_), .A2(KEYINPUT55), .A3(new_n268_), .A4(new_n269_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(KEYINPUT56), .B1(new_n774_), .B2(new_n285_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT56), .ZN(new_n776_));
  AOI211_X1 g575(.A(new_n776_), .B(new_n284_), .C1(new_n772_), .C2(new_n773_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n768_), .B1(new_n775_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT58), .ZN(new_n779_));
  OR2_X1    g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n779_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n780_), .A2(new_n606_), .A3(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT121), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n783_), .A2(KEYINPUT57), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n288_), .A2(new_n291_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n765_), .A2(new_n321_), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n785_), .A2(KEYINPUT120), .A3(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(KEYINPUT120), .B1(new_n785_), .B2(new_n786_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n322_), .B(new_n291_), .C1(new_n775_), .C2(new_n777_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n784_), .B1(new_n791_), .B2(new_n684_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n784_), .ZN(new_n793_));
  AOI211_X1 g592(.A(new_n256_), .B(new_n793_), .C1(new_n789_), .C2(new_n790_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n782_), .B1(new_n792_), .B2(new_n794_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT123), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(new_n341_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT54), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n798_), .A2(KEYINPUT118), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT117), .ZN(new_n800_));
  INV_X1    g599(.A(new_n711_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n800_), .B1(new_n710_), .B2(new_n801_), .ZN(new_n802_));
  AOI211_X1 g601(.A(KEYINPUT117), .B(new_n711_), .C1(new_n709_), .C2(new_n292_), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n605_), .B(new_n799_), .C1(new_n802_), .C2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(KEYINPUT117), .B1(new_n295_), .B2(new_n711_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n710_), .A2(new_n800_), .A3(new_n801_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n606_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  XOR2_X1   g606(.A(KEYINPUT118), .B(KEYINPUT54), .Z(new_n808_));
  OAI21_X1  g607(.A(new_n804_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  AOI211_X1 g609(.A(new_n596_), .B(new_n757_), .C1(new_n797_), .C2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(G113gat), .B1(new_n811_), .B2(new_n322_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n809_), .B1(new_n795_), .B2(new_n341_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n813_), .A2(new_n596_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT59), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n814_), .A2(new_n815_), .A3(new_n756_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n797_), .A2(new_n810_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n818_), .A2(new_n560_), .A3(new_n756_), .ZN(new_n819_));
  AOI211_X1 g618(.A(new_n323_), .B(new_n817_), .C1(new_n819_), .C2(KEYINPUT59), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n812_), .B1(new_n820_), .B2(G113gat), .ZN(G1340gat));
  OAI211_X1 g620(.A(new_n295_), .B(new_n816_), .C1(new_n811_), .C2(new_n815_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(G120gat), .ZN(new_n823_));
  INV_X1    g622(.A(G120gat), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n824_), .B1(new_n710_), .B2(KEYINPUT60), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n811_), .B(new_n825_), .C1(KEYINPUT60), .C2(new_n824_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n823_), .A2(new_n826_), .ZN(G1341gat));
  AOI21_X1  g626(.A(G127gat), .B1(new_n811_), .B2(new_n656_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n817_), .B1(new_n819_), .B2(KEYINPUT59), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n656_), .A2(G127gat), .ZN(new_n830_));
  XOR2_X1   g629(.A(new_n830_), .B(KEYINPUT124), .Z(new_n831_));
  AOI21_X1  g630(.A(new_n828_), .B1(new_n829_), .B2(new_n831_), .ZN(G1342gat));
  AOI21_X1  g631(.A(G134gat), .B1(new_n811_), .B2(new_n257_), .ZN(new_n833_));
  AOI211_X1 g632(.A(new_n605_), .B(new_n817_), .C1(new_n819_), .C2(KEYINPUT59), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n833_), .B1(new_n834_), .B2(G134gat), .ZN(G1343gat));
  NAND2_X1  g634(.A1(new_n818_), .A2(new_n561_), .ZN(new_n836_));
  NOR3_X1   g635(.A1(new_n836_), .A2(new_n388_), .A3(new_n682_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n837_), .A2(new_n353_), .A3(new_n322_), .ZN(new_n838_));
  AOI211_X1 g637(.A(new_n388_), .B(new_n595_), .C1(new_n797_), .C2(new_n810_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n839_), .A2(new_n322_), .A3(new_n722_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(G141gat), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n838_), .A2(new_n841_), .ZN(G1344gat));
  NAND3_X1  g641(.A1(new_n837_), .A2(new_n354_), .A3(new_n295_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n839_), .A2(new_n295_), .A3(new_n722_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(G148gat), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n845_), .ZN(G1345gat));
  AOI21_X1  g645(.A(new_n595_), .B1(new_n797_), .B2(new_n810_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n847_), .A2(new_n387_), .A3(new_n656_), .A4(new_n722_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(KEYINPUT61), .B(G155gat), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n848_), .B(new_n849_), .ZN(G1346gat));
  INV_X1    g649(.A(G162gat), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n648_), .A2(new_n851_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n839_), .A2(new_n257_), .A3(new_n722_), .ZN(new_n853_));
  AOI22_X1  g652(.A1(new_n837_), .A2(new_n852_), .B1(new_n853_), .B2(new_n851_), .ZN(G1347gat));
  NAND2_X1  g653(.A1(new_n682_), .A2(new_n388_), .ZN(new_n855_));
  NOR4_X1   g654(.A1(new_n813_), .A2(new_n323_), .A3(new_n596_), .A4(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(KEYINPUT125), .B1(new_n856_), .B2(new_n315_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n813_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n855_), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n858_), .A2(new_n322_), .A3(new_n560_), .A4(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT125), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(new_n861_), .A3(G169gat), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n857_), .A2(new_n862_), .A3(KEYINPUT62), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n856_), .A2(new_n452_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT62), .ZN(new_n865_));
  OAI211_X1 g664(.A(KEYINPUT125), .B(new_n865_), .C1(new_n856_), .C2(new_n315_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n863_), .A2(new_n864_), .A3(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(KEYINPUT126), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT126), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n863_), .A2(new_n869_), .A3(new_n864_), .A4(new_n866_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n868_), .A2(new_n870_), .ZN(G1348gat));
  AOI21_X1  g670(.A(new_n596_), .B1(new_n797_), .B2(new_n810_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n872_), .A2(G176gat), .A3(new_n295_), .A4(new_n859_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n814_), .A2(new_n859_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n436_), .B1(new_n874_), .B2(new_n710_), .ZN(new_n875_));
  AND2_X1   g674(.A1(new_n873_), .A2(new_n875_), .ZN(G1349gat));
  NOR2_X1   g675(.A1(new_n874_), .A2(new_n341_), .ZN(new_n877_));
  MUX2_X1   g676(.A(G183gat), .B(new_n447_), .S(new_n877_), .Z(G1350gat));
  OAI21_X1  g677(.A(G190gat), .B1(new_n874_), .B2(new_n605_), .ZN(new_n879_));
  AND2_X1   g678(.A1(new_n879_), .A2(KEYINPUT127), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n879_), .A2(KEYINPUT127), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n257_), .A2(new_n415_), .ZN(new_n882_));
  OAI22_X1  g681(.A1(new_n880_), .A2(new_n881_), .B1(new_n874_), .B2(new_n882_), .ZN(G1351gat));
  NAND3_X1  g682(.A1(new_n847_), .A2(new_n322_), .A3(new_n859_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g684(.A1(new_n847_), .A2(new_n295_), .A3(new_n859_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(G204gat), .ZN(G1353gat));
  NAND3_X1  g686(.A1(new_n847_), .A2(new_n656_), .A3(new_n859_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(KEYINPUT63), .B(G211gat), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n890_), .B1(new_n888_), .B2(new_n891_), .ZN(G1354gat));
  NOR2_X1   g691(.A1(new_n836_), .A2(new_n855_), .ZN(new_n893_));
  INV_X1    g692(.A(G218gat), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n605_), .A2(new_n894_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n847_), .A2(new_n257_), .A3(new_n859_), .ZN(new_n896_));
  AOI22_X1  g695(.A1(new_n893_), .A2(new_n895_), .B1(new_n896_), .B2(new_n894_), .ZN(G1355gat));
endmodule


