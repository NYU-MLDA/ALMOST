//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 1 1 1 1 1 1 0 0 1 0 1 0 0 1 1 1 0 0 0 0 0 0 0 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 0 0 0 0 1 0 1 1 1 0 1 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n641_, new_n642_, new_n643_, new_n645_, new_n646_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n663_, new_n664_, new_n665_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n683_, new_n684_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n792_, new_n793_, new_n794_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n813_, new_n814_, new_n815_, new_n816_, new_n818_,
    new_n819_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n845_, new_n846_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_;
  NOR2_X1   g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G169gat), .A2(G176gat), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n203_), .A2(KEYINPUT24), .A3(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n206_), .A2(KEYINPUT78), .ZN(new_n207_));
  OR2_X1    g006(.A1(new_n203_), .A2(KEYINPUT24), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT23), .ZN(new_n210_));
  AND2_X1   g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n206_), .A2(KEYINPUT78), .ZN(new_n212_));
  INV_X1    g011(.A(G190gat), .ZN(new_n213_));
  OR3_X1    g012(.A1(new_n213_), .A2(KEYINPUT77), .A3(KEYINPUT26), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT25), .B(G183gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT26), .B1(new_n213_), .B2(KEYINPUT77), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n214_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n207_), .A2(new_n211_), .A3(new_n212_), .A4(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n210_), .B1(G183gat), .B2(G190gat), .ZN(new_n219_));
  INV_X1    g018(.A(G176gat), .ZN(new_n220_));
  INV_X1    g019(.A(G169gat), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT22), .B1(new_n221_), .B2(KEYINPUT79), .ZN(new_n222_));
  OR2_X1    g021(.A1(new_n221_), .A2(KEYINPUT22), .ZN(new_n223_));
  OAI211_X1 g022(.A(new_n220_), .B(new_n222_), .C1(new_n223_), .C2(KEYINPUT79), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n219_), .A2(new_n204_), .A3(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n218_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT30), .ZN(new_n227_));
  XOR2_X1   g026(.A(KEYINPUT80), .B(KEYINPUT81), .Z(new_n228_));
  XNOR2_X1  g027(.A(new_n227_), .B(new_n228_), .ZN(new_n229_));
  XOR2_X1   g028(.A(G71gat), .B(G99gat), .Z(new_n230_));
  NAND2_X1  g029(.A1(G227gat), .A2(G233gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n230_), .B(new_n231_), .ZN(new_n232_));
  XOR2_X1   g031(.A(G15gat), .B(G43gat), .Z(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n229_), .B(new_n234_), .ZN(new_n235_));
  OR2_X1    g034(.A1(new_n235_), .A2(KEYINPUT83), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(KEYINPUT83), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G127gat), .B(G134gat), .ZN(new_n238_));
  INV_X1    g037(.A(G113gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(G120gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n242_));
  XOR2_X1   g041(.A(new_n241_), .B(new_n242_), .Z(new_n243_));
  NAND3_X1  g042(.A1(new_n236_), .A2(new_n237_), .A3(new_n243_), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n237_), .A2(new_n243_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  XOR2_X1   g045(.A(G211gat), .B(G218gat), .Z(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT85), .B(G197gat), .ZN(new_n249_));
  INV_X1    g048(.A(G204gat), .ZN(new_n250_));
  OR3_X1    g049(.A1(new_n249_), .A2(KEYINPUT86), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(G197gat), .ZN(new_n252_));
  OAI21_X1  g051(.A(KEYINPUT86), .B1(new_n249_), .B2(new_n250_), .ZN(new_n253_));
  AND3_X1   g052(.A1(new_n251_), .A2(new_n252_), .A3(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT87), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n248_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT21), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n251_), .A2(new_n252_), .A3(new_n253_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n257_), .B1(new_n258_), .B2(KEYINPUT87), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n256_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G197gat), .A2(G204gat), .ZN(new_n261_));
  OAI211_X1 g060(.A(KEYINPUT21), .B(new_n261_), .C1(new_n249_), .C2(G204gat), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n262_), .B(new_n248_), .C1(new_n258_), .C2(KEYINPUT21), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n260_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G155gat), .A2(G162gat), .ZN(new_n265_));
  OR2_X1    g064(.A1(G155gat), .A2(G162gat), .ZN(new_n266_));
  NOR2_X1   g065(.A1(G141gat), .A2(G148gat), .ZN(new_n267_));
  XOR2_X1   g066(.A(new_n267_), .B(KEYINPUT3), .Z(new_n268_));
  NAND2_X1  g067(.A1(G141gat), .A2(G148gat), .ZN(new_n269_));
  XOR2_X1   g068(.A(new_n269_), .B(KEYINPUT2), .Z(new_n270_));
  OAI211_X1 g069(.A(new_n265_), .B(new_n266_), .C1(new_n268_), .C2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n265_), .A2(KEYINPUT1), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT84), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n265_), .A2(KEYINPUT84), .A3(KEYINPUT1), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n274_), .A2(new_n275_), .A3(new_n266_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n265_), .A2(KEYINPUT1), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n269_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n271_), .B1(new_n267_), .B2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT29), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n264_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(G50gat), .ZN(new_n282_));
  INV_X1    g081(.A(G50gat), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n264_), .A2(new_n283_), .A3(new_n280_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n282_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G78gat), .B(G106gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n279_), .A2(KEYINPUT29), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT28), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G228gat), .A2(G233gat), .ZN(new_n290_));
  INV_X1    g089(.A(G22gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n289_), .B(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n286_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n282_), .A2(new_n294_), .A3(new_n284_), .ZN(new_n295_));
  AND3_X1   g094(.A1(new_n287_), .A2(new_n293_), .A3(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n293_), .B1(new_n287_), .B2(new_n295_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT20), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G226gat), .A2(G233gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT19), .ZN(new_n301_));
  AOI211_X1 g100(.A(new_n299_), .B(new_n301_), .C1(new_n264_), .C2(new_n226_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n247_), .B1(new_n254_), .B2(new_n257_), .ZN(new_n303_));
  AOI22_X1  g102(.A1(new_n259_), .A2(new_n256_), .B1(new_n303_), .B2(new_n262_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT22), .B(G169gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(new_n220_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n219_), .A2(new_n204_), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT88), .ZN(new_n308_));
  OR2_X1    g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n308_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT26), .B(G190gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n215_), .A2(new_n311_), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n211_), .A2(new_n205_), .ZN(new_n313_));
  AOI22_X1  g112(.A1(new_n309_), .A2(new_n310_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n304_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n226_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n260_), .A2(new_n316_), .A3(new_n263_), .ZN(new_n317_));
  OAI211_X1 g116(.A(new_n317_), .B(KEYINPUT20), .C1(new_n304_), .C2(new_n314_), .ZN(new_n318_));
  AOI22_X1  g117(.A1(new_n302_), .A2(new_n315_), .B1(new_n318_), .B2(new_n301_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G64gat), .B(G92gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G8gat), .B(G36gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT90), .B1(new_n319_), .B2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n318_), .A2(new_n301_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n299_), .B1(new_n264_), .B2(new_n226_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n301_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n327_), .A2(new_n328_), .A3(new_n315_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n326_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT90), .ZN(new_n331_));
  INV_X1    g130(.A(new_n324_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n330_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  AND2_X1   g132(.A1(new_n325_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n319_), .A2(new_n324_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n241_), .B(new_n279_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G225gat), .A2(G233gat), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT4), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n241_), .A2(new_n341_), .A3(new_n279_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n342_), .B1(new_n336_), .B2(new_n341_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n340_), .B1(new_n343_), .B2(new_n339_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G1gat), .B(G29gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(G85gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT0), .ZN(new_n347_));
  INV_X1    g146(.A(G57gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(KEYINPUT33), .B1(new_n344_), .B2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n337_), .A2(new_n338_), .ZN(new_n351_));
  OAI211_X1 g150(.A(new_n342_), .B(new_n339_), .C1(new_n336_), .C2(new_n341_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n351_), .A2(new_n352_), .A3(new_n349_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n350_), .A2(new_n353_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n351_), .A2(new_n352_), .A3(KEYINPUT33), .A4(new_n349_), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n334_), .A2(new_n335_), .A3(new_n354_), .A4(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n324_), .A2(KEYINPUT32), .ZN(new_n357_));
  XOR2_X1   g156(.A(new_n357_), .B(KEYINPUT91), .Z(new_n358_));
  NAND3_X1  g157(.A1(new_n319_), .A2(KEYINPUT92), .A3(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n326_), .A2(new_n329_), .A3(new_n358_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT92), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n359_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n351_), .A2(new_n352_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n349_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(new_n353_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n313_), .A2(new_n312_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n304_), .A2(new_n368_), .A3(new_n307_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n327_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(new_n301_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT93), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n370_), .A2(KEYINPUT93), .A3(new_n301_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT94), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n375_), .B1(new_n318_), .B2(new_n301_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n314_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n299_), .B1(new_n377_), .B2(new_n264_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n378_), .A2(KEYINPUT94), .A3(new_n328_), .A4(new_n317_), .ZN(new_n379_));
  AOI22_X1  g178(.A1(new_n373_), .A2(new_n374_), .B1(new_n376_), .B2(new_n379_), .ZN(new_n380_));
  OAI211_X1 g179(.A(new_n363_), .B(new_n367_), .C1(new_n380_), .C2(new_n357_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n298_), .B1(new_n356_), .B2(new_n381_), .ZN(new_n382_));
  OAI211_X1 g181(.A(KEYINPUT27), .B(new_n335_), .C1(new_n380_), .C2(new_n324_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n325_), .A2(new_n335_), .A3(new_n333_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT27), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NOR3_X1   g185(.A1(new_n296_), .A2(new_n297_), .A3(new_n367_), .ZN(new_n387_));
  AND3_X1   g186(.A1(new_n383_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n246_), .B1(new_n382_), .B2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT95), .ZN(new_n390_));
  AND2_X1   g189(.A1(new_n383_), .A2(new_n386_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n298_), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n367_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n246_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n393_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT95), .ZN(new_n397_));
  OAI211_X1 g196(.A(new_n397_), .B(new_n246_), .C1(new_n382_), .C2(new_n388_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n390_), .A2(new_n396_), .A3(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G120gat), .B(G148gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT5), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(G176gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(G204gat), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT69), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(G106gat), .ZN(new_n406_));
  INV_X1    g205(.A(G99gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT10), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT10), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(G99gat), .ZN(new_n410_));
  AND3_X1   g209(.A1(new_n408_), .A2(new_n410_), .A3(KEYINPUT64), .ZN(new_n411_));
  AOI21_X1  g210(.A(KEYINPUT64), .B1(new_n408_), .B2(new_n410_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n406_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(G85gat), .ZN(new_n414_));
  INV_X1    g213(.A(G92gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G85gat), .A2(G92gat), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n416_), .A2(KEYINPUT9), .A3(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n417_), .A2(KEYINPUT9), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G99gat), .A2(G106gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(KEYINPUT6), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT6), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n422_), .A2(G99gat), .A3(G106gat), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n419_), .B1(new_n421_), .B2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n413_), .A2(new_n418_), .A3(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n421_), .A2(new_n423_), .ZN(new_n426_));
  OAI21_X1  g225(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT7), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n428_), .A2(new_n407_), .A3(new_n406_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n426_), .A2(new_n427_), .A3(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT8), .ZN(new_n431_));
  AND3_X1   g230(.A1(new_n416_), .A2(KEYINPUT65), .A3(new_n417_), .ZN(new_n432_));
  AND3_X1   g231(.A1(new_n430_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n431_), .B1(new_n430_), .B2(new_n432_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n425_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT66), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT66), .ZN(new_n437_));
  OAI211_X1 g236(.A(new_n425_), .B(new_n437_), .C1(new_n433_), .C2(new_n434_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  AND2_X1   g238(.A1(G57gat), .A2(G64gat), .ZN(new_n440_));
  NOR2_X1   g239(.A1(G57gat), .A2(G64gat), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT11), .ZN(new_n443_));
  AOI22_X1  g242(.A1(new_n442_), .A2(new_n443_), .B1(G71gat), .B2(G78gat), .ZN(new_n444_));
  OAI21_X1  g243(.A(KEYINPUT67), .B1(new_n442_), .B2(new_n443_), .ZN(new_n445_));
  INV_X1    g244(.A(G71gat), .ZN(new_n446_));
  INV_X1    g245(.A(G78gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT67), .ZN(new_n449_));
  OAI211_X1 g248(.A(new_n449_), .B(KEYINPUT11), .C1(new_n440_), .C2(new_n441_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n444_), .A2(new_n445_), .A3(new_n448_), .A4(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(G71gat), .A2(G78gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G57gat), .B(G64gat), .ZN(new_n453_));
  OAI211_X1 g252(.A(new_n448_), .B(new_n452_), .C1(new_n453_), .C2(KEYINPUT11), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n449_), .B1(new_n453_), .B2(KEYINPUT11), .ZN(new_n455_));
  INV_X1    g254(.A(new_n450_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n454_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  AND2_X1   g256(.A1(new_n451_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n439_), .A2(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n458_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n461_));
  OAI211_X1 g260(.A(G230gat), .B(G233gat), .C1(new_n460_), .C2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n435_), .A2(new_n458_), .A3(KEYINPUT12), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT68), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n435_), .A2(new_n458_), .A3(KEYINPUT68), .A4(KEYINPUT12), .ZN(new_n466_));
  AOI22_X1  g265(.A1(new_n465_), .A2(new_n466_), .B1(new_n439_), .B2(new_n459_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G230gat), .A2(G233gat), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT12), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n469_), .B1(new_n439_), .B2(new_n459_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n467_), .A2(new_n468_), .A3(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n405_), .B1(new_n462_), .B2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n471_), .A2(new_n462_), .A3(new_n403_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT70), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT70), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n471_), .A2(new_n462_), .A3(new_n475_), .A4(new_n403_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n472_), .B1(new_n474_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT71), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  AOI211_X1 g278(.A(KEYINPUT71), .B(new_n472_), .C1(new_n474_), .C2(new_n476_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT13), .ZN(new_n481_));
  OR3_X1    g280(.A1(new_n479_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n481_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G113gat), .B(G141gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(new_n221_), .ZN(new_n487_));
  INV_X1    g286(.A(G197gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  AND2_X1   g288(.A1(G229gat), .A2(G233gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(KEYINPUT73), .B(G8gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(G1gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT14), .ZN(new_n493_));
  XOR2_X1   g292(.A(G15gat), .B(G22gat), .Z(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n493_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(G1gat), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n494_), .B1(new_n492_), .B2(KEYINPUT14), .ZN(new_n498_));
  INV_X1    g297(.A(G1gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n497_), .A2(G8gat), .A3(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(G8gat), .B1(new_n497_), .B2(new_n500_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G29gat), .B(G36gat), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n504_), .A2(G43gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(G43gat), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n505_), .A2(G50gat), .A3(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(G50gat), .B1(new_n505_), .B2(new_n506_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NOR3_X1   g309(.A1(new_n502_), .A2(new_n503_), .A3(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n509_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(new_n507_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n497_), .A2(new_n500_), .ZN(new_n514_));
  INV_X1    g313(.A(G8gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n513_), .B1(new_n516_), .B2(new_n501_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n490_), .B1(new_n511_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT15), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n519_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n512_), .A2(new_n507_), .A3(KEYINPUT15), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n522_), .A2(new_n501_), .A3(new_n516_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n510_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n490_), .B(KEYINPUT75), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n523_), .A2(new_n524_), .A3(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n518_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT76), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n489_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n489_), .ZN(new_n531_));
  AOI211_X1 g330(.A(KEYINPUT76), .B(new_n531_), .C1(new_n518_), .C2(new_n527_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n485_), .A2(new_n533_), .ZN(new_n534_));
  AND2_X1   g333(.A1(new_n399_), .A2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G127gat), .B(G155gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT16), .ZN(new_n537_));
  INV_X1    g336(.A(G183gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(G211gat), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n541_), .A2(KEYINPUT74), .A3(KEYINPUT17), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n516_), .A2(new_n501_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G231gat), .A2(G233gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(new_n459_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n541_), .A2(KEYINPUT17), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n542_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n548_), .B1(new_n542_), .B2(new_n546_), .ZN(new_n549_));
  AOI22_X1  g348(.A1(new_n439_), .A2(new_n510_), .B1(new_n522_), .B2(new_n435_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G232gat), .A2(G233gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT34), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n550_), .B1(KEYINPUT35), .B2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(KEYINPUT35), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G190gat), .B(G218gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT72), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(G134gat), .ZN(new_n558_));
  INV_X1    g357(.A(G162gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n555_), .B1(KEYINPUT36), .B2(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n560_), .B(KEYINPUT36), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n562_), .B1(new_n563_), .B2(new_n555_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT37), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n535_), .A2(new_n549_), .A3(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT96), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n568_), .A2(new_n499_), .A3(new_n367_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT97), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT38), .ZN(new_n571_));
  OR3_X1    g370(.A1(new_n569_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n570_), .B1(new_n569_), .B2(new_n571_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n564_), .B(KEYINPUT98), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n535_), .A2(new_n574_), .A3(new_n549_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n499_), .B1(new_n575_), .B2(new_n367_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n569_), .B1(new_n571_), .B2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n572_), .A2(new_n573_), .A3(new_n577_), .ZN(G1324gat));
  INV_X1    g377(.A(new_n391_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n515_), .B1(new_n575_), .B2(new_n579_), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n580_), .B(KEYINPUT39), .Z(new_n581_));
  INV_X1    g380(.A(new_n491_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n568_), .A2(new_n582_), .A3(new_n579_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT40), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n581_), .A2(new_n583_), .A3(KEYINPUT40), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(G1325gat));
  INV_X1    g387(.A(G15gat), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n568_), .A2(new_n589_), .A3(new_n395_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n575_), .ZN(new_n591_));
  OAI21_X1  g390(.A(G15gat), .B1(new_n591_), .B2(new_n246_), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n592_), .A2(KEYINPUT99), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(KEYINPUT99), .ZN(new_n594_));
  AND3_X1   g393(.A1(new_n593_), .A2(KEYINPUT41), .A3(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(KEYINPUT41), .B1(new_n593_), .B2(new_n594_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n590_), .B1(new_n595_), .B2(new_n596_), .ZN(G1326gat));
  XOR2_X1   g396(.A(new_n298_), .B(KEYINPUT100), .Z(new_n598_));
  AOI21_X1  g397(.A(new_n291_), .B1(new_n575_), .B2(new_n598_), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n599_), .B(KEYINPUT42), .Z(new_n600_));
  NAND3_X1  g399(.A1(new_n568_), .A2(new_n291_), .A3(new_n598_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(G1327gat));
  NOR2_X1   g401(.A1(new_n574_), .A2(new_n549_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n535_), .A2(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(G29gat), .B1(new_n604_), .B2(new_n367_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT102), .ZN(new_n606_));
  INV_X1    g405(.A(new_n533_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n549_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n484_), .A2(new_n607_), .A3(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT101), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT43), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n399_), .A2(new_n611_), .A3(new_n565_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n611_), .B1(new_n399_), .B2(new_n565_), .ZN(new_n613_));
  OAI211_X1 g412(.A(new_n606_), .B(new_n610_), .C1(new_n612_), .C2(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(KEYINPUT44), .B1(new_n614_), .B2(KEYINPUT103), .ZN(new_n615_));
  AOI21_X1  g414(.A(KEYINPUT102), .B1(KEYINPUT103), .B2(KEYINPUT44), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n399_), .A2(new_n565_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(KEYINPUT43), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n399_), .A2(new_n611_), .A3(new_n565_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n616_), .B1(new_n620_), .B2(new_n610_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n615_), .A2(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n622_), .A2(new_n394_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n605_), .B1(new_n623_), .B2(G29gat), .ZN(G1328gat));
  OAI21_X1  g423(.A(new_n579_), .B1(new_n615_), .B2(new_n621_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(G36gat), .ZN(new_n626_));
  INV_X1    g425(.A(G36gat), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n604_), .A2(KEYINPUT45), .A3(new_n627_), .A4(new_n579_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT45), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n535_), .A2(new_n627_), .A3(new_n603_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n629_), .B1(new_n630_), .B2(new_n391_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n628_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n626_), .A2(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(KEYINPUT46), .B1(new_n634_), .B2(KEYINPUT104), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n632_), .B1(new_n625_), .B2(G36gat), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT104), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT46), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n636_), .A2(new_n637_), .A3(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n635_), .A2(new_n639_), .ZN(G1329gat));
  OAI21_X1  g439(.A(new_n395_), .B1(new_n615_), .B2(new_n621_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n246_), .A2(G43gat), .ZN(new_n642_));
  AOI22_X1  g441(.A1(new_n641_), .A2(G43gat), .B1(new_n604_), .B2(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g443(.A(G50gat), .B1(new_n622_), .B2(new_n392_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n604_), .A2(new_n283_), .A3(new_n598_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(G1331gat));
  NOR2_X1   g446(.A1(new_n608_), .A2(new_n607_), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n399_), .A2(new_n574_), .A3(new_n485_), .A4(new_n648_), .ZN(new_n649_));
  NOR3_X1   g448(.A1(new_n649_), .A2(new_n348_), .A3(new_n394_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n399_), .A2(new_n533_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT105), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n485_), .A2(new_n549_), .A3(new_n566_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n651_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n654_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(new_n367_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n650_), .B1(new_n656_), .B2(new_n348_), .ZN(G1332gat));
  INV_X1    g456(.A(G64gat), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n655_), .A2(new_n658_), .A3(new_n579_), .ZN(new_n659_));
  OAI21_X1  g458(.A(G64gat), .B1(new_n649_), .B2(new_n391_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT48), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n659_), .A2(new_n661_), .ZN(G1333gat));
  NAND3_X1  g461(.A1(new_n655_), .A2(new_n446_), .A3(new_n395_), .ZN(new_n663_));
  OAI21_X1  g462(.A(G71gat), .B1(new_n649_), .B2(new_n246_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT49), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n663_), .A2(new_n665_), .ZN(G1334gat));
  NAND3_X1  g465(.A1(new_n655_), .A2(new_n447_), .A3(new_n598_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n598_), .ZN(new_n668_));
  OAI21_X1  g467(.A(G78gat), .B1(new_n649_), .B2(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT50), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n667_), .A2(new_n670_), .ZN(G1335gat));
  NAND3_X1  g470(.A1(new_n651_), .A2(new_n485_), .A3(new_n603_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n414_), .B1(new_n672_), .B2(new_n394_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT106), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n484_), .A2(new_n549_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n620_), .A2(new_n533_), .A3(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT107), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n620_), .A2(KEYINPUT107), .A3(new_n533_), .A4(new_n675_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n394_), .A2(new_n414_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n674_), .B1(new_n680_), .B2(new_n681_), .ZN(G1336gat));
  NAND3_X1  g481(.A1(new_n680_), .A2(G92gat), .A3(new_n579_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n415_), .B1(new_n672_), .B2(new_n391_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n683_), .A2(new_n684_), .ZN(G1337gat));
  NOR2_X1   g484(.A1(new_n411_), .A2(new_n412_), .ZN(new_n686_));
  NOR3_X1   g485(.A1(new_n672_), .A2(new_n686_), .A3(new_n246_), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n687_), .B(KEYINPUT108), .Z(new_n688_));
  NAND3_X1  g487(.A1(new_n678_), .A2(new_n395_), .A3(new_n679_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(G99gat), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI21_X1  g491(.A(G106gat), .B1(new_n676_), .B2(new_n392_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT110), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  OAI211_X1 g494(.A(KEYINPUT110), .B(G106gat), .C1(new_n676_), .C2(new_n392_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n695_), .A2(KEYINPUT52), .A3(new_n696_), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n672_), .A2(G106gat), .A3(new_n392_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT109), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT52), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n693_), .A2(new_n694_), .A3(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n697_), .A2(new_n699_), .A3(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(KEYINPUT53), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT53), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n697_), .A2(new_n704_), .A3(new_n699_), .A4(new_n701_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(G1339gat));
  AOI21_X1  g505(.A(new_n533_), .B1(new_n474_), .B2(new_n476_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n468_), .B1(new_n467_), .B2(new_n470_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT55), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n471_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n467_), .A2(KEYINPUT55), .A3(new_n468_), .A4(new_n470_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n405_), .ZN(new_n713_));
  AOI21_X1  g512(.A(KEYINPUT56), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT56), .ZN(new_n715_));
  AOI211_X1 g514(.A(new_n715_), .B(new_n405_), .C1(new_n710_), .C2(new_n711_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n707_), .B1(new_n714_), .B2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(KEYINPUT111), .ZN(new_n718_));
  OR3_X1    g517(.A1(new_n511_), .A2(new_n517_), .A3(new_n525_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n523_), .A2(new_n524_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(new_n525_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n531_), .B1(new_n719_), .B2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n528_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n722_), .B1(new_n723_), .B2(new_n531_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n724_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT111), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n707_), .B(new_n726_), .C1(new_n714_), .C2(new_n716_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n718_), .A2(new_n725_), .A3(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(new_n574_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT57), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n714_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n716_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT112), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n732_), .A2(new_n733_), .A3(new_n734_), .ZN(new_n735_));
  AOI22_X1  g534(.A1(new_n716_), .A2(KEYINPUT112), .B1(new_n474_), .B2(new_n476_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n735_), .A2(new_n724_), .A3(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT113), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n738_), .A2(KEYINPUT58), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n739_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n735_), .A2(new_n736_), .A3(new_n741_), .A4(new_n724_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n740_), .A2(new_n565_), .A3(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n728_), .A2(new_n574_), .A3(KEYINPUT57), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n731_), .A2(new_n743_), .A3(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(KEYINPUT114), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT114), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n731_), .A2(new_n743_), .A3(new_n747_), .A4(new_n744_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n746_), .A2(new_n608_), .A3(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n484_), .A2(new_n566_), .A3(new_n648_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT54), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n749_), .A2(KEYINPUT115), .A3(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(KEYINPUT115), .B1(new_n749_), .B2(new_n751_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n393_), .A2(new_n367_), .A3(new_n395_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n754_), .A2(KEYINPUT116), .A3(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n749_), .A2(new_n751_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT115), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n749_), .A2(KEYINPUT115), .A3(new_n751_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n760_), .A2(new_n761_), .A3(new_n756_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT116), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n757_), .A2(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(G113gat), .B1(new_n765_), .B2(new_n607_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT117), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n752_), .A2(new_n753_), .A3(new_n755_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT59), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n767_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n745_), .A2(new_n608_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n751_), .A2(new_n771_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n772_), .A2(new_n756_), .A3(new_n773_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT119), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n762_), .A2(KEYINPUT117), .A3(KEYINPUT59), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n770_), .A2(new_n775_), .A3(new_n776_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n533_), .A2(new_n239_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n766_), .B1(new_n777_), .B2(new_n778_), .ZN(G1340gat));
  NAND4_X1  g578(.A1(new_n770_), .A2(new_n485_), .A3(new_n775_), .A4(new_n776_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(G120gat), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT60), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n782_), .B1(new_n484_), .B2(G120gat), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n765_), .B(new_n783_), .C1(new_n782_), .C2(G120gat), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n781_), .A2(new_n784_), .ZN(G1341gat));
  AOI21_X1  g584(.A(G127gat), .B1(new_n765_), .B2(new_n549_), .ZN(new_n786_));
  INV_X1    g585(.A(G127gat), .ZN(new_n787_));
  OAI21_X1  g586(.A(KEYINPUT120), .B1(new_n608_), .B2(new_n787_), .ZN(new_n788_));
  AND4_X1   g587(.A1(new_n775_), .A2(new_n770_), .A3(new_n776_), .A4(new_n788_), .ZN(new_n789_));
  OR2_X1    g588(.A1(new_n787_), .A2(KEYINPUT120), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n786_), .B1(new_n789_), .B2(new_n790_), .ZN(G1342gat));
  INV_X1    g590(.A(new_n574_), .ZN(new_n792_));
  AOI21_X1  g591(.A(G134gat), .B1(new_n765_), .B2(new_n792_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n565_), .A2(G134gat), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n793_), .B1(new_n777_), .B2(new_n794_), .ZN(G1343gat));
  NOR2_X1   g594(.A1(new_n395_), .A2(new_n392_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  NOR3_X1   g596(.A1(new_n752_), .A2(new_n753_), .A3(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(new_n367_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n800_), .A2(new_n607_), .A3(new_n391_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(G141gat), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n799_), .A2(new_n579_), .ZN(new_n803_));
  INV_X1    g602(.A(G141gat), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n803_), .A2(new_n804_), .A3(new_n607_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n802_), .A2(new_n805_), .ZN(G1344gat));
  NAND3_X1  g605(.A1(new_n800_), .A2(new_n485_), .A3(new_n391_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(KEYINPUT121), .B(G148gat), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n808_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n803_), .A2(new_n485_), .A3(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n811_), .ZN(G1345gat));
  XNOR2_X1  g611(.A(KEYINPUT61), .B(G155gat), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n813_), .B1(new_n803_), .B2(new_n549_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n813_), .ZN(new_n815_));
  NOR4_X1   g614(.A1(new_n799_), .A2(new_n579_), .A3(new_n608_), .A4(new_n815_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n814_), .A2(new_n816_), .ZN(G1346gat));
  NAND2_X1  g616(.A1(new_n803_), .A2(new_n792_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n566_), .A2(new_n559_), .ZN(new_n819_));
  AOI22_X1  g618(.A1(new_n818_), .A2(new_n559_), .B1(new_n803_), .B2(new_n819_), .ZN(G1347gat));
  INV_X1    g619(.A(KEYINPUT62), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n598_), .B1(new_n751_), .B2(new_n771_), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n246_), .A2(new_n391_), .A3(new_n367_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n824_), .A2(new_n533_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n821_), .B1(new_n825_), .B2(new_n221_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n305_), .ZN(new_n827_));
  OAI211_X1 g626(.A(KEYINPUT62), .B(G169gat), .C1(new_n824_), .C2(new_n533_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n826_), .A2(new_n827_), .A3(new_n828_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n829_), .B(KEYINPUT122), .ZN(G1348gat));
  NAND4_X1  g629(.A1(new_n760_), .A2(new_n392_), .A3(new_n761_), .A4(new_n823_), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n831_), .A2(new_n220_), .A3(new_n484_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT123), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n832_), .A2(new_n833_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n824_), .ZN(new_n836_));
  AOI21_X1  g635(.A(G176gat), .B1(new_n836_), .B2(new_n485_), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n834_), .A2(new_n835_), .A3(new_n837_), .ZN(G1349gat));
  INV_X1    g637(.A(KEYINPUT124), .ZN(new_n839_));
  OR3_X1    g638(.A1(new_n831_), .A2(new_n839_), .A3(new_n608_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n839_), .B1(new_n831_), .B2(new_n608_), .ZN(new_n841_));
  AND3_X1   g640(.A1(new_n840_), .A2(new_n538_), .A3(new_n841_), .ZN(new_n842_));
  NOR3_X1   g641(.A1(new_n824_), .A2(new_n215_), .A3(new_n608_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n842_), .A2(new_n843_), .ZN(G1350gat));
  NAND3_X1  g643(.A1(new_n836_), .A2(new_n792_), .A3(new_n311_), .ZN(new_n845_));
  OAI21_X1  g644(.A(G190gat), .B1(new_n824_), .B2(new_n566_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(G1351gat));
  NOR2_X1   g646(.A1(new_n391_), .A2(new_n367_), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n754_), .A2(new_n607_), .A3(new_n796_), .A4(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT125), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n488_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT126), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n852_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n760_), .A2(new_n761_), .A3(new_n796_), .A4(new_n848_), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n850_), .B(new_n852_), .C1(new_n854_), .C2(new_n533_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n851_), .B1(new_n853_), .B2(new_n856_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n854_), .A2(new_n533_), .ZN(new_n858_));
  AOI21_X1  g657(.A(G197gat), .B1(new_n858_), .B2(KEYINPUT125), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n850_), .B1(new_n854_), .B2(new_n533_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(KEYINPUT126), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n859_), .A2(new_n855_), .A3(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n857_), .A2(new_n862_), .ZN(G1352gat));
  INV_X1    g662(.A(new_n854_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n485_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n250_), .A2(KEYINPUT127), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n865_), .B(new_n866_), .ZN(G1353gat));
  AOI211_X1 g666(.A(KEYINPUT63), .B(G211gat), .C1(new_n864_), .C2(new_n549_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(KEYINPUT63), .B(G211gat), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n854_), .A2(new_n608_), .A3(new_n869_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n868_), .A2(new_n870_), .ZN(G1354gat));
  INV_X1    g670(.A(G218gat), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n854_), .A2(new_n872_), .A3(new_n566_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n864_), .A2(new_n792_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n873_), .B1(new_n874_), .B2(new_n872_), .ZN(G1355gat));
endmodule


