//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 0 0 0 0 0 0 0 1 0 0 0 0 0 0 1 0 1 0 0 1 0 1 0 1 1 0 0 1 0 1 0 1 0 1 0 0 1 1 0 1 0 1 1 0 0 0 1 0 1 0 1 1 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n591_, new_n592_, new_n593_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n663_, new_n664_, new_n665_, new_n666_, new_n668_,
    new_n669_, new_n670_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n812_, new_n813_, new_n814_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n822_,
    new_n823_, new_n825_, new_n826_, new_n827_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n865_, new_n866_, new_n868_, new_n869_, new_n870_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n882_, new_n883_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  NOR2_X1   g001(.A1(new_n202_), .A2(KEYINPUT23), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT73), .B(KEYINPUT23), .ZN(new_n204_));
  INV_X1    g003(.A(new_n202_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT74), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n203_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n208_), .B1(new_n207_), .B2(new_n206_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT25), .B(G183gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT26), .B(G190gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  XOR2_X1   g011(.A(G169gat), .B(G176gat), .Z(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT24), .ZN(new_n214_));
  OR3_X1    g013(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n209_), .A2(new_n212_), .A3(new_n214_), .A4(new_n215_), .ZN(new_n216_));
  MUX2_X1   g015(.A(KEYINPUT23), .B(new_n204_), .S(new_n205_), .Z(new_n217_));
  INV_X1    g016(.A(G183gat), .ZN(new_n218_));
  INV_X1    g017(.A(G190gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n217_), .A2(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n222_));
  INV_X1    g021(.A(G169gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n222_), .B(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n221_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n216_), .A2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(KEYINPUT30), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT75), .B(G43gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G227gat), .A2(G233gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(G15gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(G71gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n230_), .B(new_n233_), .ZN(new_n234_));
  XOR2_X1   g033(.A(G127gat), .B(G134gat), .Z(new_n235_));
  XOR2_X1   g034(.A(G113gat), .B(G120gat), .Z(new_n236_));
  OR2_X1    g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT76), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n238_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n235_), .A2(new_n236_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n239_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT31), .ZN(new_n243_));
  INV_X1    g042(.A(G99gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  OR2_X1    g044(.A1(new_n234_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n234_), .A2(new_n245_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT28), .ZN(new_n249_));
  NOR2_X1   g048(.A1(G155gat), .A2(G162gat), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT77), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n250_), .B(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n252_), .B1(G155gat), .B2(G162gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G141gat), .A2(G148gat), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT78), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  AND2_X1   g055(.A1(new_n256_), .A2(KEYINPUT2), .ZN(new_n257_));
  OR2_X1    g056(.A1(G141gat), .A2(G148gat), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n258_), .A2(KEYINPUT3), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(KEYINPUT3), .ZN(new_n260_));
  OAI211_X1 g059(.A(new_n259_), .B(new_n260_), .C1(new_n256_), .C2(KEYINPUT2), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n253_), .B1(new_n257_), .B2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G155gat), .A2(G162gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT1), .ZN(new_n264_));
  OAI211_X1 g063(.A(new_n258_), .B(new_n254_), .C1(new_n252_), .C2(new_n264_), .ZN(new_n265_));
  AND2_X1   g064(.A1(new_n262_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT29), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n249_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n262_), .A2(new_n265_), .ZN(new_n269_));
  NOR3_X1   g068(.A1(new_n269_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n268_), .A2(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G22gat), .B(G50gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n271_), .A2(new_n272_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(KEYINPUT79), .B1(new_n273_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n273_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT79), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G211gat), .B(G218gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT80), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G197gat), .B(G204gat), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT21), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  AND2_X1   g083(.A1(new_n282_), .A2(new_n283_), .ZN(new_n285_));
  OR3_X1    g084(.A1(new_n281_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n281_), .A2(new_n284_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT81), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G228gat), .A2(G233gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n269_), .A2(KEYINPUT29), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n290_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G78gat), .B(G106gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT82), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n292_), .A2(new_n288_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n296_), .A2(G228gat), .A3(G233gat), .ZN(new_n297_));
  AND3_X1   g096(.A1(new_n293_), .A2(new_n295_), .A3(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n295_), .B1(new_n293_), .B2(new_n297_), .ZN(new_n299_));
  OAI22_X1  g098(.A1(new_n276_), .A2(new_n279_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n293_), .A2(new_n297_), .ZN(new_n301_));
  AND2_X1   g100(.A1(new_n301_), .A2(new_n294_), .ZN(new_n302_));
  OR3_X1    g101(.A1(new_n302_), .A2(new_n298_), .A3(new_n277_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n300_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT33), .ZN(new_n305_));
  OR2_X1    g104(.A1(new_n266_), .A2(new_n242_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n237_), .A2(new_n241_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n262_), .A2(new_n265_), .A3(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G225gat), .A2(G233gat), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n310_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT87), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n306_), .A2(new_n314_), .A3(KEYINPUT4), .A4(new_n308_), .ZN(new_n315_));
  OAI211_X1 g114(.A(KEYINPUT4), .B(new_n308_), .C1(new_n266_), .C2(new_n242_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT87), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n266_), .A2(new_n242_), .ZN(new_n318_));
  XOR2_X1   g117(.A(KEYINPUT88), .B(KEYINPUT4), .Z(new_n319_));
  AND3_X1   g118(.A1(new_n318_), .A2(KEYINPUT89), .A3(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(KEYINPUT89), .B1(new_n318_), .B2(new_n319_), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n315_), .B(new_n317_), .C1(new_n320_), .C2(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n313_), .B1(new_n322_), .B2(new_n312_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G1gat), .B(G29gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(G85gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT0), .B(G57gat), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n325_), .B(new_n326_), .Z(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n305_), .B1(new_n323_), .B2(new_n328_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n327_), .B1(new_n310_), .B2(new_n312_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n330_), .B1(new_n322_), .B2(new_n312_), .ZN(new_n331_));
  AND2_X1   g130(.A1(new_n329_), .A2(new_n331_), .ZN(new_n332_));
  AND2_X1   g131(.A1(new_n315_), .A2(new_n317_), .ZN(new_n333_));
  OR2_X1    g132(.A1(new_n320_), .A2(new_n321_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n311_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  OAI211_X1 g134(.A(KEYINPUT33), .B(new_n327_), .C1(new_n335_), .C2(new_n313_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT83), .B(KEYINPUT24), .ZN(new_n337_));
  OR3_X1    g136(.A1(new_n337_), .A2(G169gat), .A3(G176gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n213_), .A2(new_n337_), .ZN(new_n339_));
  AND4_X1   g138(.A1(new_n217_), .A2(new_n338_), .A3(new_n212_), .A4(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n209_), .A2(new_n220_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n340_), .B1(new_n341_), .B2(new_n225_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n288_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT84), .ZN(new_n344_));
  OR3_X1    g143(.A1(new_n342_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n344_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT20), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n288_), .B(KEYINPUT81), .ZN(new_n349_));
  INV_X1    g148(.A(new_n227_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n348_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n347_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G226gat), .A2(G233gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT19), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n348_), .B1(new_n290_), .B2(new_n227_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n342_), .A2(new_n343_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT85), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n354_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n357_), .A2(new_n358_), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n356_), .A2(new_n360_), .A3(new_n361_), .A4(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G8gat), .B(G36gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT18), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G64gat), .B(G92gat), .ZN(new_n366_));
  XOR2_X1   g165(.A(new_n365_), .B(new_n366_), .Z(new_n367_));
  NAND3_X1  g166(.A1(new_n355_), .A2(new_n363_), .A3(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n367_), .ZN(new_n369_));
  OAI211_X1 g168(.A(KEYINPUT20), .B(new_n361_), .C1(new_n349_), .C2(new_n350_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n362_), .ZN(new_n371_));
  NOR3_X1   g170(.A1(new_n370_), .A2(new_n371_), .A3(new_n359_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n361_), .B1(new_n347_), .B2(new_n351_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n369_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT86), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n368_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n375_), .B1(new_n368_), .B2(new_n374_), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n332_), .B(new_n336_), .C1(new_n376_), .C2(new_n377_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n327_), .B1(new_n335_), .B2(new_n313_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n323_), .A2(new_n328_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n367_), .A2(KEYINPUT32), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n355_), .A2(new_n363_), .A3(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT90), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n356_), .A2(new_n357_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(new_n354_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n387_), .B1(new_n352_), .B2(new_n354_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n388_), .A2(KEYINPUT32), .A3(new_n367_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n355_), .A2(KEYINPUT90), .A3(new_n363_), .A4(new_n382_), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n381_), .A2(new_n385_), .A3(new_n389_), .A4(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n304_), .B1(new_n378_), .B2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n388_), .A2(new_n369_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n393_), .A2(KEYINPUT27), .A3(new_n368_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n368_), .A2(new_n374_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT27), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n394_), .A2(new_n397_), .ZN(new_n398_));
  AND2_X1   g197(.A1(new_n300_), .A2(new_n303_), .ZN(new_n399_));
  NOR3_X1   g198(.A1(new_n398_), .A2(new_n399_), .A3(new_n381_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n248_), .B1(new_n392_), .B2(new_n400_), .ZN(new_n401_));
  AND2_X1   g200(.A1(new_n394_), .A2(new_n397_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(new_n399_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n248_), .A2(new_n381_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n401_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G85gat), .A2(G92gat), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n408_), .A2(KEYINPUT9), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G99gat), .A2(G106gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT6), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT6), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n412_), .A2(G99gat), .A3(G106gat), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n409_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n414_));
  OR2_X1    g213(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n415_));
  INV_X1    g214(.A(G106gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n415_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(G85gat), .ZN(new_n419_));
  INV_X1    g218(.A(G92gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  AND2_X1   g220(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n422_));
  NOR2_X1   g221(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n421_), .B(new_n408_), .C1(new_n422_), .C2(new_n423_), .ZN(new_n424_));
  AND3_X1   g223(.A1(new_n414_), .A2(new_n418_), .A3(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n421_), .A2(new_n408_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n412_), .B1(G99gat), .B2(G106gat), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n410_), .A2(KEYINPUT6), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT7), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n431_), .A2(new_n244_), .A3(new_n416_), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n427_), .B1(new_n430_), .B2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT8), .ZN(new_n436_));
  OAI211_X1 g235(.A(new_n433_), .B(new_n432_), .C1(new_n428_), .C2(new_n429_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT8), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n437_), .A2(new_n438_), .A3(new_n427_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n425_), .B1(new_n436_), .B2(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G57gat), .B(G64gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G71gat), .B(G78gat), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n441_), .A2(new_n442_), .A3(KEYINPUT11), .ZN(new_n443_));
  INV_X1    g242(.A(new_n442_), .ZN(new_n444_));
  INV_X1    g243(.A(G64gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(G57gat), .ZN(new_n446_));
  INV_X1    g245(.A(G57gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(G64gat), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n446_), .A2(new_n448_), .A3(KEYINPUT11), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n444_), .A2(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n441_), .A2(KEYINPUT11), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n443_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  AND2_X1   g251(.A1(KEYINPUT65), .A2(KEYINPUT12), .ZN(new_n453_));
  NOR2_X1   g252(.A1(KEYINPUT65), .A2(KEYINPUT12), .ZN(new_n454_));
  OAI22_X1  g253(.A1(new_n440_), .A2(new_n452_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n414_), .A2(new_n418_), .A3(new_n424_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n433_), .ZN(new_n457_));
  NOR3_X1   g256(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n411_), .A2(new_n413_), .ZN(new_n460_));
  AOI211_X1 g259(.A(KEYINPUT8), .B(new_n426_), .C1(new_n459_), .C2(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n438_), .B1(new_n437_), .B2(new_n427_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n456_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n452_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n454_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n463_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n466_));
  OAI211_X1 g265(.A(new_n452_), .B(new_n456_), .C1(new_n461_), .C2(new_n462_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G230gat), .A2(G233gat), .ZN(new_n468_));
  AND3_X1   g267(.A1(new_n467_), .A2(KEYINPUT66), .A3(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(KEYINPUT66), .B1(new_n467_), .B2(new_n468_), .ZN(new_n470_));
  OAI211_X1 g269(.A(new_n455_), .B(new_n466_), .C1(new_n469_), .C2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n468_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n440_), .A2(new_n452_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n467_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n472_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  AND2_X1   g274(.A1(new_n471_), .A2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G120gat), .B(G148gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT5), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G176gat), .B(G204gat), .ZN(new_n479_));
  XOR2_X1   g278(.A(new_n478_), .B(new_n479_), .Z(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n476_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT67), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  OR2_X1    g283(.A1(new_n476_), .A2(new_n481_), .ZN(new_n485_));
  AND2_X1   g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  XOR2_X1   g285(.A(KEYINPUT68), .B(KEYINPUT13), .Z(new_n487_));
  AND2_X1   g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT68), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n489_), .A2(KEYINPUT13), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n486_), .A2(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n488_), .A2(new_n491_), .ZN(new_n492_));
  XOR2_X1   g291(.A(G29gat), .B(G36gat), .Z(new_n493_));
  XOR2_X1   g292(.A(G43gat), .B(G50gat), .Z(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT15), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G15gat), .B(G22gat), .ZN(new_n497_));
  INV_X1    g296(.A(G1gat), .ZN(new_n498_));
  INV_X1    g297(.A(G8gat), .ZN(new_n499_));
  OAI21_X1  g298(.A(KEYINPUT14), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n497_), .A2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G1gat), .B(G8gat), .ZN(new_n502_));
  XOR2_X1   g301(.A(new_n501_), .B(new_n502_), .Z(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n496_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n495_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n505_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G229gat), .A2(G233gat), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n507_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(KEYINPUT72), .ZN(new_n511_));
  AOI21_X1  g310(.A(KEYINPUT70), .B1(new_n503_), .B2(new_n495_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT71), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n504_), .A2(new_n506_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(new_n509_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n511_), .A2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G113gat), .B(G141gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G169gat), .B(G197gat), .ZN(new_n519_));
  XOR2_X1   g318(.A(new_n518_), .B(new_n519_), .Z(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n517_), .A2(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n511_), .A2(new_n516_), .A3(new_n520_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n492_), .A2(new_n525_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n407_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G232gat), .A2(G233gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT34), .ZN(new_n529_));
  OAI22_X1  g328(.A1(new_n463_), .A2(new_n506_), .B1(KEYINPUT35), .B2(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n530_), .B1(new_n496_), .B2(new_n463_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n529_), .A2(KEYINPUT35), .ZN(new_n532_));
  XOR2_X1   g331(.A(new_n531_), .B(new_n532_), .Z(new_n533_));
  XNOR2_X1  g332(.A(G190gat), .B(G218gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G134gat), .B(G162gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n536_), .A2(KEYINPUT36), .ZN(new_n537_));
  AND2_X1   g336(.A1(new_n536_), .A2(KEYINPUT36), .ZN(new_n538_));
  NOR3_X1   g337(.A1(new_n533_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n533_), .A2(new_n537_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT37), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G231gat), .A2(G233gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n503_), .B(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(new_n452_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  XOR2_X1   g345(.A(G127gat), .B(G155gat), .Z(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(KEYINPUT16), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G183gat), .B(G211gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT17), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n551_), .A2(KEYINPUT69), .ZN(new_n552_));
  OR3_X1    g351(.A1(new_n546_), .A2(new_n550_), .A3(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n550_), .A2(new_n551_), .ZN(new_n554_));
  OAI211_X1 g353(.A(new_n546_), .B(new_n554_), .C1(new_n550_), .C2(new_n552_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n542_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n527_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n381_), .ZN(new_n559_));
  NOR3_X1   g358(.A1(new_n558_), .A2(G1gat), .A3(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(KEYINPUT91), .B(KEYINPUT38), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  NOR4_X1   g361(.A1(new_n248_), .A2(new_n398_), .A3(new_n381_), .A4(new_n304_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n336_), .A2(new_n329_), .A3(new_n331_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n395_), .A2(KEYINPUT86), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n368_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n564_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  AND4_X1   g366(.A1(new_n381_), .A2(new_n385_), .A3(new_n389_), .A4(new_n390_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n399_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n399_), .A2(new_n381_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(new_n402_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n563_), .B1(new_n572_), .B2(new_n248_), .ZN(new_n573_));
  NOR3_X1   g372(.A1(new_n573_), .A2(new_n556_), .A3(new_n541_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n526_), .B(KEYINPUT92), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(G1gat), .B1(new_n576_), .B2(new_n559_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n562_), .A2(new_n577_), .ZN(G1324gat));
  NAND2_X1  g377(.A1(new_n398_), .A2(new_n499_), .ZN(new_n579_));
  OR3_X1    g378(.A1(new_n558_), .A2(KEYINPUT93), .A3(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(KEYINPUT93), .B1(new_n558_), .B2(new_n579_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(G8gat), .B1(new_n576_), .B2(new_n402_), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n583_), .A2(KEYINPUT39), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT39), .ZN(new_n585_));
  OAI211_X1 g384(.A(new_n585_), .B(G8gat), .C1(new_n576_), .C2(new_n402_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n582_), .B1(new_n584_), .B2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT40), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(G1325gat));
  OAI21_X1  g389(.A(G15gat), .B1(new_n576_), .B2(new_n248_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT41), .ZN(new_n592_));
  NOR3_X1   g391(.A1(new_n558_), .A2(G15gat), .A3(new_n248_), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n592_), .A2(new_n593_), .ZN(G1326gat));
  OAI21_X1  g393(.A(G22gat), .B1(new_n576_), .B2(new_n399_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT42), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n399_), .A2(G22gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT94), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n596_), .B1(new_n558_), .B2(new_n598_), .ZN(G1327gat));
  INV_X1    g398(.A(new_n541_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n556_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n527_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(G29gat), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n604_), .A2(new_n605_), .A3(new_n381_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n542_), .ZN(new_n607_));
  OAI21_X1  g406(.A(KEYINPUT43), .B1(new_n573_), .B2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT43), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n407_), .A2(new_n609_), .A3(new_n542_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n610_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n575_), .A2(new_n556_), .ZN(new_n612_));
  OR2_X1    g411(.A1(KEYINPUT95), .A2(KEYINPUT44), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n611_), .A2(new_n612_), .A3(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n613_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n615_));
  NOR3_X1   g414(.A1(new_n614_), .A2(new_n615_), .A3(new_n559_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n606_), .B1(new_n616_), .B2(new_n605_), .ZN(G1328gat));
  INV_X1    g416(.A(KEYINPUT46), .ZN(new_n618_));
  NOR3_X1   g417(.A1(new_n614_), .A2(new_n615_), .A3(new_n402_), .ZN(new_n619_));
  INV_X1    g418(.A(G36gat), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n603_), .A2(G36gat), .A3(new_n402_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(KEYINPUT96), .B(KEYINPUT45), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(KEYINPUT97), .Z(new_n624_));
  XNOR2_X1  g423(.A(new_n622_), .B(new_n624_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n618_), .B1(new_n621_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n624_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n622_), .B(new_n627_), .ZN(new_n628_));
  OAI211_X1 g427(.A(new_n628_), .B(KEYINPUT46), .C1(new_n620_), .C2(new_n619_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n626_), .A2(new_n629_), .ZN(G1329gat));
  NOR3_X1   g429(.A1(new_n603_), .A2(G43gat), .A3(new_n248_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n614_), .A2(new_n615_), .A3(new_n248_), .ZN(new_n633_));
  INV_X1    g432(.A(G43gat), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n632_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(KEYINPUT98), .B(KEYINPUT47), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n637_), .ZN(new_n638_));
  OAI211_X1 g437(.A(new_n632_), .B(new_n636_), .C1(new_n633_), .C2(new_n634_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(G1330gat));
  AOI21_X1  g439(.A(G50gat), .B1(new_n604_), .B2(new_n304_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n614_), .A2(new_n615_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n304_), .A2(G50gat), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n641_), .B1(new_n642_), .B2(new_n643_), .ZN(G1331gat));
  INV_X1    g443(.A(new_n492_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n645_), .A2(new_n524_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n574_), .A2(new_n646_), .ZN(new_n647_));
  XOR2_X1   g446(.A(KEYINPUT100), .B(G57gat), .Z(new_n648_));
  NOR3_X1   g447(.A1(new_n647_), .A2(new_n559_), .A3(new_n648_), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n649_), .B(KEYINPUT101), .Z(new_n650_));
  AND2_X1   g449(.A1(new_n407_), .A2(new_n646_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(new_n557_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  OR2_X1    g452(.A1(new_n653_), .A2(KEYINPUT99), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(KEYINPUT99), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n654_), .A2(new_n381_), .A3(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n650_), .B1(new_n447_), .B2(new_n656_), .ZN(G1332gat));
  OAI21_X1  g456(.A(G64gat), .B1(new_n647_), .B2(new_n402_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(KEYINPUT102), .B(KEYINPUT48), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n658_), .B(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n653_), .A2(new_n445_), .A3(new_n398_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(G1333gat));
  OAI21_X1  g461(.A(G71gat), .B1(new_n647_), .B2(new_n248_), .ZN(new_n663_));
  XOR2_X1   g462(.A(KEYINPUT103), .B(KEYINPUT49), .Z(new_n664_));
  XNOR2_X1  g463(.A(new_n663_), .B(new_n664_), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n248_), .A2(G71gat), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n665_), .B1(new_n652_), .B2(new_n666_), .ZN(G1334gat));
  OAI21_X1  g466(.A(G78gat), .B1(new_n647_), .B2(new_n399_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT50), .ZN(new_n669_));
  OR2_X1    g468(.A1(new_n399_), .A2(G78gat), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n669_), .B1(new_n652_), .B2(new_n670_), .ZN(G1335gat));
  NAND2_X1  g470(.A1(new_n646_), .A2(new_n556_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n672_), .B1(new_n608_), .B2(new_n610_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n673_), .A2(new_n381_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n651_), .A2(new_n602_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n381_), .A2(new_n419_), .ZN(new_n676_));
  OAI22_X1  g475(.A1(new_n674_), .A2(new_n419_), .B1(new_n675_), .B2(new_n676_), .ZN(G1336gat));
  AND2_X1   g476(.A1(new_n673_), .A2(new_n398_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n398_), .A2(new_n420_), .ZN(new_n679_));
  OAI22_X1  g478(.A1(new_n678_), .A2(new_n420_), .B1(new_n675_), .B2(new_n679_), .ZN(G1337gat));
  INV_X1    g479(.A(new_n248_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n244_), .B1(new_n673_), .B2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n415_), .A2(new_n417_), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n675_), .A2(new_n683_), .A3(new_n248_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n682_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT104), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(KEYINPUT51), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n685_), .B(new_n687_), .ZN(G1338gat));
  AOI211_X1 g487(.A(new_n399_), .B(new_n672_), .C1(new_n608_), .C2(new_n610_), .ZN(new_n689_));
  OAI21_X1  g488(.A(KEYINPUT105), .B1(new_n689_), .B2(new_n416_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n672_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n609_), .B1(new_n407_), .B2(new_n542_), .ZN(new_n692_));
  AOI211_X1 g491(.A(KEYINPUT43), .B(new_n607_), .C1(new_n401_), .C2(new_n406_), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n304_), .B(new_n691_), .C1(new_n692_), .C2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT105), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n694_), .A2(new_n695_), .A3(G106gat), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n690_), .A2(KEYINPUT52), .A3(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT52), .ZN(new_n698_));
  OAI211_X1 g497(.A(KEYINPUT105), .B(new_n698_), .C1(new_n689_), .C2(new_n416_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n675_), .A2(G106gat), .A3(new_n399_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(KEYINPUT106), .B(KEYINPUT53), .ZN(new_n702_));
  AND4_X1   g501(.A1(new_n697_), .A2(new_n699_), .A3(new_n701_), .A4(new_n702_), .ZN(new_n703_));
  AOI211_X1 g502(.A(new_n695_), .B(KEYINPUT52), .C1(new_n694_), .C2(G106gat), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n704_), .A2(new_n700_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n702_), .B1(new_n705_), .B2(new_n697_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n703_), .A2(new_n706_), .ZN(G1339gat));
  INV_X1    g506(.A(KEYINPUT107), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n708_), .B1(new_n524_), .B2(new_n556_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n525_), .A2(KEYINPUT107), .A3(new_n601_), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n645_), .A2(new_n607_), .A3(new_n709_), .A4(new_n710_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(KEYINPUT108), .B(KEYINPUT54), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n711_), .B(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT57), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n515_), .A2(new_n508_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n507_), .A2(KEYINPUT115), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n507_), .A2(KEYINPUT115), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(new_n509_), .ZN(new_n718_));
  OAI211_X1 g517(.A(new_n715_), .B(new_n521_), .C1(new_n716_), .C2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(new_n523_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n486_), .A2(new_n720_), .ZN(new_n721_));
  XOR2_X1   g520(.A(KEYINPUT109), .B(KEYINPUT55), .Z(new_n722_));
  NAND2_X1  g521(.A1(new_n467_), .A2(new_n468_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT66), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n467_), .A2(KEYINPUT66), .A3(new_n468_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n463_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n453_), .A2(new_n454_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n729_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n728_), .A2(new_n730_), .ZN(new_n731_));
  AOI211_X1 g530(.A(KEYINPUT110), .B(new_n722_), .C1(new_n727_), .C2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT110), .ZN(new_n733_));
  INV_X1    g532(.A(new_n722_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n471_), .B2(new_n734_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n732_), .A2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT112), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n455_), .A2(new_n467_), .A3(new_n466_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT111), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n455_), .A2(KEYINPUT111), .A3(new_n467_), .A4(new_n466_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n740_), .A2(new_n472_), .A3(new_n741_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n727_), .A2(KEYINPUT55), .A3(new_n731_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n736_), .A2(new_n737_), .A3(new_n744_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n469_), .A2(new_n470_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n455_), .A2(new_n466_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n734_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(KEYINPUT110), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n471_), .A2(new_n733_), .A3(new_n734_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n471_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n468_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n753_));
  AOI22_X1  g552(.A1(KEYINPUT55), .A2(new_n752_), .B1(new_n753_), .B2(new_n741_), .ZN(new_n754_));
  AOI21_X1  g553(.A(KEYINPUT112), .B1(new_n751_), .B2(new_n754_), .ZN(new_n755_));
  OAI211_X1 g554(.A(KEYINPUT56), .B(new_n480_), .C1(new_n745_), .C2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT114), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT56), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n758_), .A2(KEYINPUT114), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n737_), .B1(new_n736_), .B2(new_n744_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n751_), .A2(KEYINPUT112), .A3(new_n754_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n481_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n759_), .B1(new_n762_), .B2(KEYINPUT113), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n480_), .B1(new_n745_), .B2(new_n755_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT113), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n764_), .A2(new_n765_), .A3(new_n758_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n757_), .A2(new_n763_), .A3(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n484_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n525_), .A2(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n721_), .B1(new_n767_), .B2(new_n769_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n714_), .B1(new_n770_), .B2(new_n541_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT117), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n768_), .A2(new_n720_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n762_), .A2(KEYINPUT56), .ZN(new_n774_));
  INV_X1    g573(.A(new_n756_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n773_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT58), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  OAI211_X1 g577(.A(KEYINPUT58), .B(new_n773_), .C1(new_n774_), .C2(new_n775_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n778_), .A2(new_n542_), .A3(new_n779_), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n771_), .A2(new_n772_), .A3(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n772_), .B1(new_n771_), .B2(new_n780_), .ZN(new_n782_));
  NOR3_X1   g581(.A1(new_n770_), .A2(new_n714_), .A3(new_n541_), .ZN(new_n783_));
  NOR3_X1   g582(.A1(new_n781_), .A2(new_n782_), .A3(new_n783_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n713_), .B1(new_n784_), .B2(new_n601_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  NOR3_X1   g585(.A1(new_n403_), .A2(new_n559_), .A3(new_n248_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n787_), .B(KEYINPUT116), .ZN(new_n788_));
  OR2_X1    g587(.A1(new_n788_), .A2(KEYINPUT59), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n771_), .A2(new_n780_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n556_), .B1(new_n790_), .B2(new_n783_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n713_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n793_), .A2(new_n788_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT59), .ZN(new_n795_));
  OAI22_X1  g594(.A1(new_n786_), .A2(new_n789_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(G113gat), .B1(new_n796_), .B2(new_n525_), .ZN(new_n797_));
  INV_X1    g596(.A(G113gat), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n794_), .A2(new_n798_), .A3(new_n524_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n797_), .A2(new_n799_), .ZN(G1340gat));
  OAI21_X1  g599(.A(G120gat), .B1(new_n796_), .B2(new_n645_), .ZN(new_n801_));
  INV_X1    g600(.A(G120gat), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n802_), .B1(new_n645_), .B2(KEYINPUT60), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n794_), .B(new_n803_), .C1(KEYINPUT60), .C2(new_n802_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n801_), .A2(new_n804_), .ZN(G1341gat));
  AND2_X1   g604(.A1(new_n601_), .A2(G127gat), .ZN(new_n806_));
  OAI221_X1 g605(.A(new_n806_), .B1(new_n794_), .B2(new_n795_), .C1(new_n786_), .C2(new_n789_), .ZN(new_n807_));
  NOR3_X1   g606(.A1(new_n793_), .A2(new_n556_), .A3(new_n788_), .ZN(new_n808_));
  OR3_X1    g607(.A1(new_n808_), .A2(KEYINPUT118), .A3(G127gat), .ZN(new_n809_));
  OAI21_X1  g608(.A(KEYINPUT118), .B1(new_n808_), .B2(G127gat), .ZN(new_n810_));
  AND3_X1   g609(.A1(new_n807_), .A2(new_n809_), .A3(new_n810_), .ZN(G1342gat));
  OAI21_X1  g610(.A(G134gat), .B1(new_n796_), .B2(new_n607_), .ZN(new_n812_));
  INV_X1    g611(.A(G134gat), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n794_), .A2(new_n813_), .A3(new_n541_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(new_n814_), .ZN(G1343gat));
  NAND2_X1  g614(.A1(new_n792_), .A2(new_n248_), .ZN(new_n816_));
  NOR3_X1   g615(.A1(new_n398_), .A2(new_n399_), .A3(new_n559_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n816_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n524_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n820_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g620(.A1(new_n819_), .A2(new_n492_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(KEYINPUT119), .B(G148gat), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n822_), .B(new_n823_), .ZN(G1345gat));
  NAND4_X1  g623(.A1(new_n792_), .A2(new_n248_), .A3(new_n601_), .A4(new_n817_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n825_), .B(KEYINPUT120), .ZN(new_n826_));
  XNOR2_X1  g625(.A(KEYINPUT61), .B(G155gat), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n826_), .B(new_n827_), .ZN(G1346gat));
  NOR3_X1   g627(.A1(new_n816_), .A2(new_n600_), .A3(new_n818_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT121), .ZN(new_n830_));
  OR3_X1    g629(.A1(new_n829_), .A2(new_n830_), .A3(G162gat), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n830_), .B1(new_n829_), .B2(G162gat), .ZN(new_n832_));
  INV_X1    g631(.A(G162gat), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n607_), .A2(new_n833_), .ZN(new_n834_));
  AOI22_X1  g633(.A1(new_n831_), .A2(new_n832_), .B1(new_n819_), .B2(new_n834_), .ZN(G1347gat));
  NAND3_X1  g634(.A1(new_n405_), .A2(new_n399_), .A3(new_n398_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n783_), .B1(new_n790_), .B2(KEYINPUT117), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n771_), .A2(new_n772_), .A3(new_n780_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n601_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n713_), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n524_), .B(new_n837_), .C1(new_n840_), .C2(new_n841_), .ZN(new_n842_));
  XOR2_X1   g641(.A(KEYINPUT22), .B(G169gat), .Z(new_n843_));
  OR2_X1    g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT62), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT122), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n842_), .A2(new_n846_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n785_), .A2(KEYINPUT122), .A3(new_n524_), .A4(new_n837_), .ZN(new_n848_));
  AND4_X1   g647(.A1(new_n845_), .A2(new_n847_), .A3(G169gat), .A4(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n223_), .B1(new_n842_), .B2(new_n846_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n845_), .B1(new_n850_), .B2(new_n848_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n844_), .B1(new_n849_), .B2(new_n851_), .ZN(G1348gat));
  NOR2_X1   g651(.A1(new_n786_), .A2(new_n836_), .ZN(new_n853_));
  AOI21_X1  g652(.A(G176gat), .B1(new_n853_), .B2(new_n492_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n793_), .A2(new_n836_), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n492_), .A2(G176gat), .ZN(new_n856_));
  AOI21_X1  g655(.A(KEYINPUT123), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  AND3_X1   g656(.A1(new_n855_), .A2(KEYINPUT123), .A3(new_n856_), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n854_), .A2(new_n857_), .A3(new_n858_), .ZN(G1349gat));
  NOR3_X1   g658(.A1(new_n793_), .A2(new_n556_), .A3(new_n836_), .ZN(new_n860_));
  OR2_X1    g659(.A1(new_n860_), .A2(KEYINPUT124), .ZN(new_n861_));
  AOI21_X1  g660(.A(G183gat), .B1(new_n860_), .B2(KEYINPUT124), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n556_), .A2(new_n210_), .ZN(new_n863_));
  AOI22_X1  g662(.A1(new_n861_), .A2(new_n862_), .B1(new_n853_), .B2(new_n863_), .ZN(G1350gat));
  NAND3_X1  g663(.A1(new_n853_), .A2(new_n211_), .A3(new_n541_), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n786_), .A2(new_n607_), .A3(new_n836_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(new_n219_), .B2(new_n866_), .ZN(G1351gat));
  NAND2_X1  g666(.A1(new_n570_), .A2(new_n398_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n816_), .A2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n524_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n492_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g672(.A(new_n868_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n556_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n792_), .A2(new_n248_), .A3(new_n874_), .A4(new_n875_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(KEYINPUT125), .ZN(new_n877_));
  NOR2_X1   g676(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n877_), .B(new_n878_), .ZN(G1354gat));
  NOR3_X1   g678(.A1(new_n816_), .A2(new_n600_), .A3(new_n868_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(KEYINPUT126), .ZN(new_n881_));
  XNOR2_X1  g680(.A(KEYINPUT127), .B(G218gat), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n607_), .A2(new_n882_), .ZN(new_n883_));
  AOI22_X1  g682(.A1(new_n881_), .A2(new_n882_), .B1(new_n869_), .B2(new_n883_), .ZN(G1355gat));
endmodule


