//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 0 1 1 1 0 1 1 0 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 0 0 1 1 0 1 1 1 0 1 0 0 1 1 0 0 1 1 1 1 1 1 1 0 1 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n737_, new_n738_, new_n739_, new_n740_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n761_, new_n762_, new_n764_,
    new_n765_, new_n766_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n784_,
    new_n785_, new_n786_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n883_, new_n885_, new_n886_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n918_, new_n919_, new_n920_, new_n922_, new_n923_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n934_, new_n935_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n943_, new_n944_, new_n945_;
  XNOR2_X1  g000(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G232gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT35), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT73), .ZN(new_n207_));
  AND2_X1   g006(.A1(G85gat), .A2(G92gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G85gat), .A2(G92gat), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT6), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n211_), .B(new_n212_), .ZN(new_n213_));
  OR3_X1    g012(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n210_), .B1(new_n213_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT67), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n217_), .A2(new_n218_), .A3(KEYINPUT8), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(KEYINPUT8), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n220_), .B(new_n210_), .C1(new_n213_), .C2(new_n216_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n219_), .A2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G29gat), .B(G36gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  XOR2_X1   g023(.A(G43gat), .B(G50gat), .Z(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G43gat), .B(G50gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n223_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n226_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  XOR2_X1   g029(.A(KEYINPUT10), .B(G99gat), .Z(new_n231_));
  INV_X1    g030(.A(KEYINPUT64), .ZN(new_n232_));
  INV_X1    g031(.A(G106gat), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n231_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT10), .B(G99gat), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT64), .B1(new_n235_), .B2(G106gat), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n213_), .B1(new_n234_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(G85gat), .ZN(new_n238_));
  INV_X1    g037(.A(G92gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G85gat), .A2(G92gat), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n240_), .A2(KEYINPUT65), .A3(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT9), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n210_), .A2(KEYINPUT65), .A3(KEYINPUT9), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n209_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n237_), .B1(new_n246_), .B2(KEYINPUT66), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n242_), .A2(new_n243_), .ZN(new_n248_));
  AOI21_X1  g047(.A(KEYINPUT9), .B1(new_n210_), .B2(KEYINPUT65), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n240_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT66), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n222_), .B(new_n230_), .C1(new_n247_), .C2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  AND3_X1   g053(.A1(new_n226_), .A2(KEYINPUT15), .A3(new_n228_), .ZN(new_n255_));
  AOI21_X1  g054(.A(KEYINPUT15), .B1(new_n226_), .B2(new_n228_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n250_), .A2(new_n251_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n246_), .A2(KEYINPUT66), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n258_), .A2(new_n259_), .A3(new_n237_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n257_), .B1(new_n260_), .B2(new_n222_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n207_), .B1(new_n254_), .B2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n204_), .A2(new_n205_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT75), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n222_), .B1(new_n247_), .B2(new_n252_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n257_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n264_), .B1(new_n267_), .B2(new_n253_), .ZN(new_n268_));
  OAI211_X1 g067(.A(new_n206_), .B(new_n262_), .C1(new_n268_), .C2(new_n207_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n206_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n254_), .A2(new_n261_), .ZN(new_n271_));
  OAI211_X1 g070(.A(KEYINPUT73), .B(new_n270_), .C1(new_n271_), .C2(new_n264_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G190gat), .B(G218gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G134gat), .B(G162gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n269_), .A2(new_n272_), .A3(KEYINPUT36), .A4(new_n275_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n275_), .A2(KEYINPUT36), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n269_), .A2(new_n272_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n277_), .B1(new_n278_), .B2(KEYINPUT74), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT74), .ZN(new_n280_));
  INV_X1    g079(.A(new_n277_), .ZN(new_n281_));
  AOI211_X1 g080(.A(new_n280_), .B(new_n281_), .C1(new_n269_), .C2(new_n272_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n276_), .B1(new_n279_), .B2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT37), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT37), .ZN(new_n285_));
  OAI211_X1 g084(.A(new_n276_), .B(new_n285_), .C1(new_n279_), .C2(new_n282_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G57gat), .B(G64gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G71gat), .B(G78gat), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n288_), .A2(new_n289_), .A3(KEYINPUT11), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n288_), .A2(KEYINPUT11), .ZN(new_n291_));
  INV_X1    g090(.A(new_n289_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n288_), .A2(KEYINPUT11), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n290_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT68), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G15gat), .B(G22gat), .ZN(new_n299_));
  INV_X1    g098(.A(G1gat), .ZN(new_n300_));
  INV_X1    g099(.A(G8gat), .ZN(new_n301_));
  OAI21_X1  g100(.A(KEYINPUT14), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n299_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G1gat), .B(G8gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G231gat), .A2(G233gat), .ZN(new_n306_));
  XOR2_X1   g105(.A(new_n306_), .B(KEYINPUT76), .Z(new_n307_));
  XOR2_X1   g106(.A(new_n305_), .B(new_n307_), .Z(new_n308_));
  XNOR2_X1  g107(.A(new_n298_), .B(new_n308_), .ZN(new_n309_));
  XOR2_X1   g108(.A(G127gat), .B(G155gat), .Z(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G183gat), .B(G211gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT17), .ZN(new_n315_));
  AND2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n314_), .A2(new_n315_), .ZN(new_n317_));
  NOR3_X1   g116(.A1(new_n309_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  XOR2_X1   g117(.A(new_n318_), .B(KEYINPUT78), .Z(new_n319_));
  INV_X1    g118(.A(new_n308_), .ZN(new_n320_));
  OR2_X1    g119(.A1(new_n320_), .A2(new_n295_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n295_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n321_), .A2(new_n317_), .A3(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n319_), .A2(new_n323_), .ZN(new_n324_));
  OR3_X1    g123(.A1(new_n287_), .A2(KEYINPUT79), .A3(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(KEYINPUT79), .B1(new_n287_), .B2(new_n324_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT12), .ZN(new_n328_));
  OR2_X1    g127(.A1(new_n295_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n265_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT69), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT69), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n265_), .A2(new_n333_), .A3(new_n330_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G230gat), .A2(G233gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n265_), .A2(new_n297_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n265_), .A2(new_n297_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n337_), .B1(new_n338_), .B2(new_n328_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n335_), .A2(new_n336_), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n337_), .ZN(new_n341_));
  OAI211_X1 g140(.A(G230gat), .B(G233gat), .C1(new_n341_), .C2(new_n338_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n340_), .A2(new_n342_), .ZN(new_n343_));
  XOR2_X1   g142(.A(G120gat), .B(G148gat), .Z(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G176gat), .B(G204gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n343_), .A2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n340_), .A2(new_n342_), .A3(new_n348_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT71), .B(KEYINPUT13), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(KEYINPUT71), .A2(KEYINPUT13), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n350_), .A2(new_n351_), .A3(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n354_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n257_), .A2(new_n305_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n359_), .B1(new_n305_), .B2(new_n230_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G229gat), .A2(G233gat), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  OR3_X1    g161(.A1(new_n360_), .A2(KEYINPUT80), .A3(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT80), .B1(new_n360_), .B2(new_n362_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n305_), .B(new_n230_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(new_n362_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n363_), .A2(new_n364_), .A3(new_n366_), .ZN(new_n367_));
  XOR2_X1   g166(.A(G113gat), .B(G141gat), .Z(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT81), .ZN(new_n369_));
  XOR2_X1   g168(.A(G169gat), .B(G197gat), .Z(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n367_), .B(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n358_), .A2(new_n373_), .ZN(new_n374_));
  AND3_X1   g173(.A1(KEYINPUT84), .A2(G183gat), .A3(G190gat), .ZN(new_n375_));
  AOI21_X1  g174(.A(KEYINPUT84), .B1(G183gat), .B2(G190gat), .ZN(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT23), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(G183gat), .ZN(new_n378_));
  INV_X1    g177(.A(G190gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G183gat), .A2(G190gat), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT23), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n377_), .A2(new_n380_), .A3(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G169gat), .A2(G176gat), .ZN(new_n385_));
  INV_X1    g184(.A(G169gat), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n386_), .A2(KEYINPUT85), .A3(KEYINPUT22), .ZN(new_n387_));
  INV_X1    g186(.A(G176gat), .ZN(new_n388_));
  AND2_X1   g187(.A1(KEYINPUT85), .A2(KEYINPUT22), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n387_), .B(new_n388_), .C1(new_n386_), .C2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT86), .ZN(new_n391_));
  AND2_X1   g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n390_), .A2(new_n391_), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n384_), .B(new_n385_), .C1(new_n392_), .C2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n379_), .A2(KEYINPUT26), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT26), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(G190gat), .ZN(new_n397_));
  AND2_X1   g196(.A1(new_n395_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n378_), .A2(KEYINPUT25), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT82), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT25), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(G183gat), .ZN(new_n403_));
  AND2_X1   g202(.A1(new_n399_), .A2(new_n403_), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n398_), .B(new_n401_), .C1(new_n404_), .C2(new_n400_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n386_), .A2(new_n388_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n406_), .A2(KEYINPUT24), .A3(new_n385_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT83), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n406_), .A2(KEYINPUT83), .A3(KEYINPUT24), .A4(new_n385_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n382_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n381_), .A2(KEYINPUT23), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  OR3_X1    g213(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n405_), .A2(new_n411_), .A3(new_n414_), .A4(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G71gat), .B(G99gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(G43gat), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n394_), .A2(new_n416_), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(G127gat), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n421_), .A2(G134gat), .ZN(new_n422_));
  INV_X1    g221(.A(G134gat), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n423_), .A2(G127gat), .ZN(new_n424_));
  INV_X1    g223(.A(G113gat), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n425_), .A2(G120gat), .ZN(new_n426_));
  INV_X1    g225(.A(G120gat), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n427_), .A2(G113gat), .ZN(new_n428_));
  OAI22_X1  g227(.A1(new_n422_), .A2(new_n424_), .B1(new_n426_), .B2(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G127gat), .B(G134gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G113gat), .B(G120gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT87), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n429_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n430_), .A2(new_n431_), .A3(KEYINPUT87), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(KEYINPUT31), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n418_), .B1(new_n394_), .B2(new_n416_), .ZN(new_n438_));
  NOR3_X1   g237(.A1(new_n420_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G227gat), .A2(G233gat), .ZN(new_n441_));
  INV_X1    g240(.A(G15gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n441_), .B(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT30), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT88), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n437_), .B1(new_n420_), .B2(new_n438_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n440_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n445_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n446_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n448_), .B1(new_n449_), .B2(new_n439_), .ZN(new_n450_));
  AND2_X1   g249(.A1(new_n447_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT29), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT89), .ZN(new_n453_));
  INV_X1    g252(.A(G155gat), .ZN(new_n454_));
  INV_X1    g253(.A(G162gat), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n453_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(KEYINPUT89), .B1(G155gat), .B2(G162gat), .ZN(new_n457_));
  AND2_X1   g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G155gat), .A2(G162gat), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT1), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n458_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(G141gat), .ZN(new_n463_));
  INV_X1    g262(.A(G148gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G141gat), .A2(G148gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n462_), .A2(new_n468_), .ZN(new_n469_));
  AND3_X1   g268(.A1(new_n456_), .A2(new_n457_), .A3(new_n459_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT90), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT3), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n472_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT2), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n466_), .A2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n476_));
  OAI21_X1  g275(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n473_), .A2(new_n475_), .A3(new_n476_), .A4(new_n477_), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n470_), .A2(new_n471_), .A3(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n471_), .B1(new_n470_), .B2(new_n478_), .ZN(new_n480_));
  OAI211_X1 g279(.A(new_n452_), .B(new_n469_), .C1(new_n479_), .C2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT28), .ZN(new_n482_));
  AND4_X1   g281(.A1(new_n475_), .A2(new_n473_), .A3(new_n476_), .A4(new_n477_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n456_), .A2(new_n457_), .A3(new_n459_), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT90), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n470_), .A2(new_n471_), .A3(new_n478_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT28), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n487_), .A2(new_n488_), .A3(new_n452_), .A4(new_n469_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G22gat), .B(G50gat), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  AND3_X1   g290(.A1(new_n482_), .A2(new_n489_), .A3(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n491_), .B1(new_n482_), .B2(new_n489_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  OR2_X1    g293(.A1(G197gat), .A2(G204gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G197gat), .A2(G204gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT21), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n495_), .A2(KEYINPUT21), .A3(new_n496_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G211gat), .B(G218gat), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n499_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  OR2_X1    g301(.A1(new_n500_), .A2(new_n501_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G228gat), .A2(G233gat), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n467_), .B1(new_n458_), .B2(new_n461_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n506_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n504_), .B(new_n505_), .C1(new_n507_), .C2(new_n452_), .ZN(new_n508_));
  AND2_X1   g307(.A1(new_n502_), .A2(new_n503_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n469_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n510_));
  XOR2_X1   g309(.A(KEYINPUT91), .B(KEYINPUT29), .Z(new_n511_));
  AOI21_X1  g310(.A(new_n509_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n508_), .B1(new_n512_), .B2(new_n505_), .ZN(new_n513_));
  XOR2_X1   g312(.A(G78gat), .B(G106gat), .Z(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n514_), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n508_), .B(new_n516_), .C1(new_n512_), .C2(new_n505_), .ZN(new_n517_));
  AND3_X1   g316(.A1(new_n494_), .A2(new_n515_), .A3(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n492_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n493_), .ZN(new_n520_));
  AOI22_X1  g319(.A1(new_n515_), .A2(new_n517_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n518_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G1gat), .B(G29gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G57gat), .B(G85gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT96), .ZN(new_n529_));
  INV_X1    g328(.A(new_n436_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n529_), .B1(new_n507_), .B2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n510_), .A2(KEYINPUT96), .A3(new_n436_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n429_), .A2(new_n432_), .ZN(new_n533_));
  AOI22_X1  g332(.A1(new_n531_), .A2(new_n532_), .B1(new_n533_), .B2(new_n507_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G225gat), .A2(G233gat), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n528_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n507_), .A2(new_n533_), .ZN(new_n537_));
  NOR3_X1   g336(.A1(new_n507_), .A2(new_n530_), .A3(new_n529_), .ZN(new_n538_));
  AOI21_X1  g337(.A(KEYINPUT96), .B1(new_n510_), .B2(new_n436_), .ZN(new_n539_));
  OAI211_X1 g338(.A(KEYINPUT4), .B(new_n537_), .C1(new_n538_), .C2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n535_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n510_), .A2(new_n436_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n541_), .B1(new_n542_), .B2(KEYINPUT4), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n540_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n536_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n528_), .ZN(new_n547_));
  AOI22_X1  g346(.A1(new_n540_), .A2(new_n544_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n546_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n399_), .A2(new_n403_), .A3(new_n395_), .A4(new_n397_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(new_n407_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(KEYINPUT93), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n377_), .A2(new_n383_), .A3(new_n415_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT93), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n550_), .A2(new_n555_), .A3(new_n407_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n552_), .A2(new_n554_), .A3(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n414_), .A2(new_n380_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n385_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(KEYINPUT22), .B(G169gat), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n559_), .B1(new_n560_), .B2(new_n388_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n558_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n557_), .A2(new_n509_), .A3(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G226gat), .A2(G233gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n563_), .A2(KEYINPUT20), .A3(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n509_), .B1(new_n394_), .B2(new_n416_), .ZN(new_n569_));
  OR2_X1    g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(G8gat), .B(G36gat), .Z(new_n571_));
  XNOR2_X1  g370(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G64gat), .B(G92gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(KEYINPUT32), .ZN(new_n577_));
  AND3_X1   g376(.A1(new_n550_), .A2(new_n555_), .A3(new_n407_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n555_), .B1(new_n550_), .B2(new_n407_), .ZN(new_n579_));
  NOR3_X1   g378(.A1(new_n578_), .A2(new_n579_), .A3(new_n553_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n561_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n581_), .B1(new_n414_), .B2(new_n380_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n504_), .B1(new_n580_), .B2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n394_), .A2(new_n416_), .A3(new_n509_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n583_), .A2(KEYINPUT20), .A3(new_n584_), .ZN(new_n585_));
  AND3_X1   g384(.A1(new_n585_), .A2(KEYINPUT94), .A3(new_n566_), .ZN(new_n586_));
  AOI21_X1  g385(.A(KEYINPUT94), .B1(new_n585_), .B2(new_n566_), .ZN(new_n587_));
  OAI211_X1 g386(.A(new_n570_), .B(new_n577_), .C1(new_n586_), .C2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(KEYINPUT98), .B(KEYINPUT20), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n563_), .A2(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n566_), .B1(new_n590_), .B2(new_n569_), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n583_), .A2(KEYINPUT20), .A3(new_n584_), .A4(new_n567_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n577_), .ZN(new_n594_));
  AOI21_X1  g393(.A(KEYINPUT99), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT99), .ZN(new_n596_));
  AOI211_X1 g395(.A(new_n596_), .B(new_n577_), .C1(new_n591_), .C2(new_n592_), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n549_), .B(new_n588_), .C1(new_n595_), .C2(new_n597_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n570_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(new_n575_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n542_), .A2(KEYINPUT4), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n601_), .A2(new_n541_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n540_), .A2(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n547_), .B1(new_n534_), .B2(new_n541_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n547_), .A2(KEYINPUT33), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n605_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n606_));
  AOI22_X1  g405(.A1(new_n603_), .A2(new_n604_), .B1(new_n606_), .B2(new_n545_), .ZN(new_n607_));
  OAI211_X1 g406(.A(new_n576_), .B(new_n570_), .C1(new_n586_), .C2(new_n587_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT33), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n543_), .B1(new_n534_), .B2(KEYINPUT4), .ZN(new_n610_));
  OAI211_X1 g409(.A(new_n537_), .B(new_n535_), .C1(new_n538_), .C2(new_n539_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(new_n547_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n609_), .B1(new_n610_), .B2(new_n612_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n600_), .A2(new_n607_), .A3(new_n608_), .A4(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n523_), .B1(new_n598_), .B2(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(KEYINPUT27), .B1(new_n600_), .B2(new_n608_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n611_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n528_), .B1(new_n610_), .B2(new_n617_), .ZN(new_n618_));
  OAI211_X1 g417(.A(new_n618_), .B(new_n546_), .C1(new_n518_), .C2(new_n521_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT27), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n620_), .B1(new_n593_), .B2(new_n575_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n608_), .A2(new_n621_), .ZN(new_n622_));
  NOR3_X1   g421(.A1(new_n616_), .A2(new_n619_), .A3(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n451_), .B1(new_n615_), .B2(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n616_), .A2(new_n622_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n451_), .A2(new_n549_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n625_), .A2(new_n522_), .A3(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n624_), .A2(new_n627_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n374_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n327_), .A2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT100), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT100), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n327_), .A2(new_n632_), .A3(new_n629_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n631_), .A2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n634_), .A2(new_n300_), .A3(new_n549_), .ZN(new_n635_));
  XOR2_X1   g434(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n636_));
  INV_X1    g435(.A(KEYINPUT103), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n600_), .A2(new_n608_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(new_n620_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n622_), .ZN(new_n640_));
  AND4_X1   g439(.A1(new_n522_), .A2(new_n639_), .A3(new_n640_), .A4(new_n626_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n604_), .A2(new_n603_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n606_), .A2(new_n545_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n613_), .A2(new_n642_), .A3(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n588_), .B1(new_n595_), .B2(new_n597_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n545_), .A2(new_n611_), .ZN(new_n646_));
  AOI22_X1  g445(.A1(new_n646_), .A2(new_n528_), .B1(new_n545_), .B2(new_n536_), .ZN(new_n647_));
  OAI22_X1  g446(.A1(new_n638_), .A2(new_n644_), .B1(new_n645_), .B2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(new_n522_), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n639_), .A2(new_n647_), .A3(new_n523_), .A4(new_n640_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n641_), .B1(new_n651_), .B2(new_n451_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n324_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n283_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n652_), .A2(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n637_), .B1(new_n656_), .B2(new_n374_), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n374_), .A2(new_n628_), .A3(new_n653_), .A4(new_n654_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n658_), .A2(KEYINPUT103), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n549_), .B1(new_n657_), .B2(new_n659_), .ZN(new_n660_));
  AOI22_X1  g459(.A1(new_n635_), .A2(new_n636_), .B1(new_n660_), .B2(G1gat), .ZN(new_n661_));
  INV_X1    g460(.A(new_n636_), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n634_), .A2(new_n300_), .A3(new_n662_), .A4(new_n549_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n663_), .A2(KEYINPUT102), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n663_), .A2(KEYINPUT102), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n661_), .B1(new_n664_), .B2(new_n665_), .ZN(G1324gat));
  NOR2_X1   g465(.A1(new_n625_), .A2(G8gat), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n631_), .A2(new_n633_), .A3(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT104), .ZN(new_n669_));
  OAI21_X1  g468(.A(G8gat), .B1(new_n658_), .B2(new_n625_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT39), .ZN(new_n671_));
  XNOR2_X1  g470(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n672_));
  AND3_X1   g471(.A1(new_n669_), .A2(new_n671_), .A3(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n672_), .B1(new_n669_), .B2(new_n671_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n673_), .A2(new_n674_), .ZN(G1325gat));
  INV_X1    g474(.A(new_n451_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n676_), .B1(new_n657_), .B2(new_n659_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT106), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n677_), .A2(new_n678_), .A3(G15gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n656_), .A2(new_n637_), .A3(new_n374_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n658_), .A2(KEYINPUT103), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n451_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(KEYINPUT106), .B1(new_n682_), .B2(new_n442_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n679_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT41), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n327_), .A2(new_n442_), .A3(new_n676_), .A4(new_n629_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n679_), .A2(new_n683_), .A3(KEYINPUT41), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n686_), .A2(new_n687_), .A3(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(KEYINPUT107), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT107), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n686_), .A2(new_n691_), .A3(new_n687_), .A4(new_n688_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n690_), .A2(new_n692_), .ZN(G1326gat));
  OAI21_X1  g492(.A(new_n523_), .B1(new_n657_), .B2(new_n659_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(G22gat), .ZN(new_n695_));
  XNOR2_X1  g494(.A(KEYINPUT108), .B(KEYINPUT42), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n695_), .B(new_n696_), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n522_), .A2(G22gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n697_), .B1(new_n630_), .B2(new_n698_), .ZN(G1327gat));
  NOR3_X1   g498(.A1(new_n652_), .A2(new_n653_), .A3(new_n654_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(new_n374_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(G29gat), .B1(new_n702_), .B2(new_n549_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n374_), .A2(new_n324_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n284_), .A2(new_n286_), .ZN(new_n705_));
  OAI21_X1  g504(.A(KEYINPUT43), .B1(new_n652_), .B2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT43), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n628_), .A2(new_n707_), .A3(new_n287_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n704_), .B1(new_n706_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n710_), .A2(KEYINPUT109), .A3(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT109), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n713_), .B1(new_n709_), .B2(KEYINPUT44), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n709_), .A2(KEYINPUT44), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n716_), .A2(new_n718_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n549_), .A2(G29gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n703_), .B1(new_n719_), .B2(new_n720_), .ZN(G1328gat));
  NOR2_X1   g520(.A1(new_n718_), .A2(new_n625_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n715_), .A2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(G36gat), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT110), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT46), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n701_), .A2(G36gat), .A3(new_n625_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT45), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n724_), .A2(new_n725_), .A3(new_n726_), .A4(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n725_), .A2(new_n726_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(KEYINPUT110), .A2(KEYINPUT46), .ZN(new_n732_));
  INV_X1    g531(.A(G36gat), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n733_), .B1(new_n715_), .B2(new_n722_), .ZN(new_n734_));
  OAI211_X1 g533(.A(new_n731_), .B(new_n732_), .C1(new_n734_), .C2(new_n728_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n730_), .A2(new_n735_), .ZN(G1329gat));
  NAND4_X1  g535(.A1(new_n715_), .A2(G43gat), .A3(new_n676_), .A4(new_n717_), .ZN(new_n737_));
  AOI21_X1  g536(.A(G43gat), .B1(new_n702_), .B2(new_n676_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g540(.A1(new_n716_), .A2(new_n522_), .A3(new_n718_), .ZN(new_n742_));
  INV_X1    g541(.A(G50gat), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n523_), .A2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT111), .ZN(new_n745_));
  OAI22_X1  g544(.A1(new_n742_), .A2(new_n743_), .B1(new_n701_), .B2(new_n745_), .ZN(G1331gat));
  NOR2_X1   g545(.A1(new_n357_), .A2(new_n372_), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n656_), .A2(G57gat), .A3(new_n549_), .A4(new_n747_), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT112), .Z(new_n749_));
  AND2_X1   g548(.A1(new_n628_), .A2(new_n747_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n327_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(G57gat), .B1(new_n752_), .B2(new_n549_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n749_), .A2(new_n753_), .ZN(G1332gat));
  NAND2_X1  g553(.A1(new_n656_), .A2(new_n747_), .ZN(new_n755_));
  OAI21_X1  g554(.A(G64gat), .B1(new_n755_), .B2(new_n625_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT48), .ZN(new_n757_));
  OR2_X1    g556(.A1(new_n625_), .A2(G64gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n757_), .B1(new_n751_), .B2(new_n758_), .ZN(G1333gat));
  OAI21_X1  g558(.A(G71gat), .B1(new_n755_), .B2(new_n451_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT49), .ZN(new_n761_));
  OR2_X1    g560(.A1(new_n451_), .A2(G71gat), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n761_), .B1(new_n751_), .B2(new_n762_), .ZN(G1334gat));
  OAI21_X1  g562(.A(G78gat), .B1(new_n755_), .B2(new_n522_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT50), .ZN(new_n765_));
  OR2_X1    g564(.A1(new_n522_), .A2(G78gat), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n765_), .B1(new_n751_), .B2(new_n766_), .ZN(G1335gat));
  NAND2_X1  g566(.A1(new_n747_), .A2(new_n324_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  AOI221_X4 g568(.A(KEYINPUT43), .B1(new_n284_), .B2(new_n286_), .C1(new_n624_), .C2(new_n627_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n707_), .B1(new_n628_), .B2(new_n287_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n769_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT113), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n706_), .A2(new_n708_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n775_), .A2(KEYINPUT113), .A3(new_n769_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(G85gat), .B1(new_n778_), .B2(new_n647_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n700_), .A2(new_n747_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n781_), .A2(new_n238_), .A3(new_n549_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n779_), .A2(new_n782_), .ZN(G1336gat));
  OAI21_X1  g582(.A(G92gat), .B1(new_n778_), .B2(new_n625_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n625_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n781_), .A2(new_n239_), .A3(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(G1337gat));
  NOR3_X1   g586(.A1(new_n780_), .A2(new_n235_), .A3(new_n451_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT113), .B1(new_n775_), .B2(new_n769_), .ZN(new_n789_));
  AOI211_X1 g588(.A(new_n773_), .B(new_n768_), .C1(new_n706_), .C2(new_n708_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n676_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(G99gat), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n788_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n791_), .A2(KEYINPUT114), .A3(G99gat), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n794_), .A2(KEYINPUT115), .A3(KEYINPUT51), .A4(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n451_), .B1(new_n774_), .B2(new_n776_), .ZN(new_n797_));
  INV_X1    g596(.A(G99gat), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n793_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n788_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n799_), .A2(new_n795_), .A3(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n802_));
  OR2_X1    g601(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n801_), .A2(new_n802_), .A3(new_n803_), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n796_), .A2(new_n804_), .ZN(G1338gat));
  OAI21_X1  g604(.A(G106gat), .B1(new_n772_), .B2(new_n522_), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n806_), .B(KEYINPUT52), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n781_), .A2(new_n233_), .A3(new_n523_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n809_), .B(new_n810_), .ZN(G1339gat));
  OR2_X1    g610(.A1(new_n367_), .A2(new_n371_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n365_), .A2(new_n361_), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n813_), .B(new_n371_), .C1(new_n360_), .C2(new_n361_), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n812_), .A2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n351_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n336_), .B1(new_n335_), .B2(new_n339_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n340_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n335_), .A2(new_n339_), .A3(KEYINPUT55), .A4(new_n336_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n349_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT56), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n821_), .A2(KEYINPUT56), .A3(new_n349_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n816_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(KEYINPUT58), .B1(new_n826_), .B2(KEYINPUT118), .ZN(new_n827_));
  AOI21_X1  g626(.A(KEYINPUT56), .B1(new_n821_), .B2(new_n349_), .ZN(new_n828_));
  AOI211_X1 g627(.A(new_n823_), .B(new_n348_), .C1(new_n819_), .C2(new_n820_), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n351_), .B(new_n815_), .C1(new_n828_), .C2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT118), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT58), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n830_), .A2(new_n831_), .A3(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n827_), .A2(new_n287_), .A3(new_n833_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n372_), .A2(new_n351_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n835_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n815_), .A2(new_n352_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n283_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT57), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n834_), .A2(new_n839_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n838_), .A2(KEYINPUT57), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n324_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n372_), .B1(new_n354_), .B2(new_n356_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n705_), .A2(new_n653_), .A3(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT54), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n844_), .B(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n842_), .A2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT59), .ZN(new_n849_));
  NOR4_X1   g648(.A1(new_n785_), .A2(new_n647_), .A3(new_n523_), .A4(new_n451_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT119), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  OR2_X1    g651(.A1(new_n850_), .A2(new_n851_), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n848_), .A2(new_n849_), .A3(new_n852_), .A4(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT57), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n836_), .A2(new_n837_), .ZN(new_n856_));
  OAI211_X1 g655(.A(KEYINPUT117), .B(new_n855_), .C1(new_n856_), .C2(new_n283_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT117), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n858_), .B1(new_n838_), .B2(KEYINPUT57), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n857_), .A2(new_n834_), .A3(new_n859_), .A4(new_n839_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n324_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n847_), .ZN(new_n862_));
  AND2_X1   g661(.A1(new_n862_), .A2(new_n850_), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n372_), .B(new_n854_), .C1(new_n863_), .C2(new_n849_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(G113gat), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n863_), .A2(new_n425_), .A3(new_n372_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(G1340gat));
  OAI211_X1 g666(.A(new_n358_), .B(new_n854_), .C1(new_n863_), .C2(new_n849_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(G120gat), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n427_), .B1(new_n357_), .B2(KEYINPUT60), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n863_), .B(new_n870_), .C1(KEYINPUT60), .C2(new_n427_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n871_), .ZN(G1341gat));
  OAI211_X1 g671(.A(new_n653_), .B(new_n854_), .C1(new_n863_), .C2(new_n849_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(G127gat), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n863_), .A2(new_n421_), .A3(new_n653_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(G1342gat));
  OAI211_X1 g675(.A(new_n287_), .B(new_n854_), .C1(new_n863_), .C2(new_n849_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(G134gat), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n863_), .A2(new_n423_), .A3(new_n283_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1343gat));
  NOR3_X1   g679(.A1(new_n676_), .A2(new_n647_), .A3(new_n522_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n862_), .A2(new_n625_), .A3(new_n881_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n882_), .A2(new_n373_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(new_n463_), .ZN(G1344gat));
  NOR2_X1   g683(.A1(new_n882_), .A2(new_n357_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(KEYINPUT120), .B(G148gat), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n885_), .B(new_n886_), .ZN(G1345gat));
  NOR2_X1   g686(.A1(new_n882_), .A2(new_n324_), .ZN(new_n888_));
  XOR2_X1   g687(.A(KEYINPUT61), .B(G155gat), .Z(new_n889_));
  XNOR2_X1  g688(.A(new_n888_), .B(new_n889_), .ZN(G1346gat));
  OAI21_X1  g689(.A(G162gat), .B1(new_n882_), .B2(new_n705_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n283_), .A2(new_n455_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n882_), .B2(new_n892_), .ZN(G1347gat));
  NAND2_X1  g692(.A1(new_n785_), .A2(new_n626_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n522_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n848_), .A2(new_n372_), .A3(new_n897_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n898_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n899_));
  INV_X1    g698(.A(new_n560_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n899_), .B1(new_n900_), .B2(new_n898_), .ZN(new_n901_));
  AOI21_X1  g700(.A(KEYINPUT62), .B1(new_n898_), .B2(G169gat), .ZN(new_n902_));
  OR2_X1    g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1348gat));
  NAND3_X1  g702(.A1(new_n848_), .A2(new_n358_), .A3(new_n897_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n388_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT121), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n523_), .B1(new_n861_), .B2(new_n847_), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n894_), .A2(new_n357_), .A3(new_n388_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n906_), .B1(new_n907_), .B2(new_n908_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n846_), .B1(new_n860_), .B2(new_n324_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n908_), .ZN(new_n911_));
  NOR4_X1   g710(.A1(new_n910_), .A2(KEYINPUT121), .A3(new_n523_), .A4(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n905_), .B1(new_n909_), .B2(new_n912_), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT122), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(new_n915_));
  OAI211_X1 g714(.A(new_n905_), .B(KEYINPUT122), .C1(new_n909_), .C2(new_n912_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(G1349gat));
  NAND2_X1  g716(.A1(new_n848_), .A2(new_n897_), .ZN(new_n918_));
  NOR3_X1   g717(.A1(new_n918_), .A2(new_n324_), .A3(new_n404_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n907_), .A2(new_n653_), .A3(new_n895_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n919_), .B1(new_n920_), .B2(new_n378_), .ZN(G1350gat));
  OAI21_X1  g720(.A(G190gat), .B1(new_n918_), .B2(new_n705_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n283_), .A2(new_n398_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n922_), .B1(new_n918_), .B2(new_n923_), .ZN(G1351gat));
  NOR3_X1   g723(.A1(new_n625_), .A2(new_n619_), .A3(new_n676_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n862_), .A2(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n926_), .ZN(new_n927_));
  AOI21_X1  g726(.A(G197gat), .B1(new_n927_), .B2(new_n372_), .ZN(new_n928_));
  NAND4_X1  g727(.A1(new_n862_), .A2(G197gat), .A3(new_n372_), .A4(new_n925_), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT123), .ZN(new_n930_));
  AND2_X1   g729(.A1(new_n929_), .A2(new_n930_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n929_), .A2(new_n930_), .ZN(new_n932_));
  NOR3_X1   g731(.A1(new_n928_), .A2(new_n931_), .A3(new_n932_), .ZN(G1352gat));
  NOR2_X1   g732(.A1(new_n926_), .A2(new_n357_), .ZN(new_n934_));
  XOR2_X1   g733(.A(KEYINPUT124), .B(G204gat), .Z(new_n935_));
  XNOR2_X1  g734(.A(new_n934_), .B(new_n935_), .ZN(G1353gat));
  NAND2_X1  g735(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n937_));
  NAND4_X1  g736(.A1(new_n862_), .A2(new_n653_), .A3(new_n925_), .A4(new_n937_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(KEYINPUT125), .B(KEYINPUT126), .ZN(new_n939_));
  NOR2_X1   g738(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n939_), .B(new_n940_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n938_), .B(new_n941_), .ZN(G1354gat));
  AOI21_X1  g741(.A(G218gat), .B1(new_n927_), .B2(new_n283_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n287_), .A2(G218gat), .ZN(new_n944_));
  XOR2_X1   g743(.A(new_n944_), .B(KEYINPUT127), .Z(new_n945_));
  AOI21_X1  g744(.A(new_n943_), .B1(new_n927_), .B2(new_n945_), .ZN(G1355gat));
endmodule


