//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 0 1 1 1 1 1 1 1 0 1 1 1 1 0 1 0 0 0 0 0 0 1 0 0 0 1 0 0 0 0 1 0 0 0 1 1 1 0 1 1 1 1 1 0 1 1 0 0 1 1 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n604_, new_n605_,
    new_n606_, new_n608_, new_n609_, new_n610_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n648_, new_n649_, new_n650_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n663_, new_n664_, new_n665_, new_n667_,
    new_n668_, new_n669_, new_n671_, new_n672_, new_n673_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n685_, new_n686_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n811_, new_n812_, new_n814_, new_n815_,
    new_n817_, new_n818_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n851_,
    new_n852_, new_n853_, new_n855_, new_n856_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_;
  INV_X1    g000(.A(KEYINPUT38), .ZN(new_n202_));
  NOR2_X1   g001(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(G169gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G183gat), .A2(G190gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n206_), .ZN(new_n208_));
  OR2_X1    g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n204_), .B1(new_n207_), .B2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT25), .B(G183gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT26), .B(G190gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  XOR2_X1   g013(.A(new_n214_), .B(KEYINPUT82), .Z(new_n215_));
  NOR3_X1   g014(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n216_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n205_), .B(KEYINPUT23), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n211_), .B1(new_n215_), .B2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G211gat), .B(G218gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(KEYINPUT91), .ZN(new_n225_));
  XOR2_X1   g024(.A(G197gat), .B(G204gat), .Z(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT21), .ZN(new_n227_));
  OR2_X1    g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(G197gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n229_), .A2(KEYINPUT89), .A3(G204gat), .ZN(new_n230_));
  OAI211_X1 g029(.A(KEYINPUT21), .B(new_n230_), .C1(new_n226_), .C2(KEYINPUT89), .ZN(new_n231_));
  XOR2_X1   g030(.A(KEYINPUT90), .B(KEYINPUT21), .Z(new_n232_));
  OAI211_X1 g031(.A(new_n225_), .B(new_n231_), .C1(new_n226_), .C2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n228_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n223_), .A2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT95), .ZN(new_n236_));
  XNOR2_X1  g035(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G226gat), .A2(G233gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT20), .ZN(new_n240_));
  INV_X1    g039(.A(new_n234_), .ZN(new_n241_));
  AND2_X1   g040(.A1(new_n221_), .A2(new_n209_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n204_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n214_), .A2(new_n221_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n220_), .ZN(new_n245_));
  OAI22_X1  g044(.A1(new_n242_), .A2(new_n243_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n240_), .B1(new_n241_), .B2(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n236_), .A2(new_n239_), .A3(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n240_), .B1(new_n234_), .B2(new_n246_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n250_), .B1(new_n234_), .B2(new_n223_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n239_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n249_), .A2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G8gat), .B(G36gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT18), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G64gat), .B(G92gat), .ZN(new_n257_));
  XOR2_X1   g056(.A(new_n256_), .B(new_n257_), .Z(new_n258_));
  XNOR2_X1  g057(.A(new_n254_), .B(new_n258_), .ZN(new_n259_));
  OR2_X1    g058(.A1(G141gat), .A2(G148gat), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT3), .B1(new_n260_), .B2(KEYINPUT87), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n260_), .A2(KEYINPUT87), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT3), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT2), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G141gat), .A2(G148gat), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n261_), .B(new_n264_), .C1(new_n265_), .C2(new_n266_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(G155gat), .A2(G162gat), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G155gat), .A2(G162gat), .ZN(new_n270_));
  AND2_X1   g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n267_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(KEYINPUT1), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT86), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  OAI211_X1 g074(.A(new_n275_), .B(new_n269_), .C1(KEYINPUT1), .C2(new_n270_), .ZN(new_n276_));
  AOI22_X1  g075(.A1(new_n276_), .A2(new_n260_), .B1(new_n265_), .B2(new_n271_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n266_), .B(KEYINPUT85), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n272_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G127gat), .B(G134gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G113gat), .B(G120gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT96), .ZN(new_n283_));
  OR2_X1    g082(.A1(new_n279_), .A2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n282_), .B(KEYINPUT83), .ZN(new_n285_));
  AOI21_X1  g084(.A(KEYINPUT97), .B1(new_n279_), .B2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT97), .ZN(new_n288_));
  NOR3_X1   g087(.A1(new_n279_), .A2(new_n288_), .A3(new_n283_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n287_), .A2(KEYINPUT4), .A3(new_n290_), .ZN(new_n291_));
  AND2_X1   g090(.A1(new_n279_), .A2(new_n285_), .ZN(new_n292_));
  OR2_X1    g091(.A1(new_n292_), .A2(KEYINPUT4), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G225gat), .A2(G233gat), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G1gat), .B(G29gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(G85gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT0), .B(G57gat), .ZN(new_n300_));
  XOR2_X1   g099(.A(new_n299_), .B(new_n300_), .Z(new_n301_));
  AOI21_X1  g100(.A(new_n289_), .B1(new_n286_), .B2(new_n284_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n302_), .A2(new_n296_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n297_), .A2(KEYINPUT33), .A3(new_n301_), .A4(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n294_), .A2(new_n295_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n301_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n307_), .B1(new_n302_), .B2(new_n295_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT99), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  OAI211_X1 g109(.A(KEYINPUT99), .B(new_n307_), .C1(new_n302_), .C2(new_n295_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n306_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  AND3_X1   g111(.A1(new_n259_), .A2(new_n305_), .A3(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n297_), .A2(new_n301_), .A3(new_n304_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT33), .ZN(new_n315_));
  AND3_X1   g114(.A1(new_n314_), .A2(KEYINPUT98), .A3(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(KEYINPUT98), .B1(new_n314_), .B2(new_n315_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n313_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n258_), .A2(KEYINPUT32), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n239_), .B1(new_n236_), .B2(new_n248_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n251_), .A2(new_n252_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n320_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT100), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT100), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n325_), .B(new_n320_), .C1(new_n321_), .C2(new_n322_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n254_), .ZN(new_n327_));
  AOI22_X1  g126(.A1(new_n324_), .A2(new_n326_), .B1(new_n327_), .B2(new_n319_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n295_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n307_), .B1(new_n329_), .B2(new_n303_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n314_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n328_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT101), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT101), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n328_), .A2(new_n331_), .A3(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n318_), .A2(new_n333_), .A3(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G78gat), .B(G106gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT92), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n241_), .B1(new_n279_), .B2(KEYINPUT29), .ZN(new_n339_));
  AOI22_X1  g138(.A1(new_n234_), .A2(KEYINPUT88), .B1(G228gat), .B2(G233gat), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n339_), .A2(new_n341_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n338_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n344_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n346_), .A2(new_n342_), .A3(new_n337_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT28), .ZN(new_n348_));
  INV_X1    g147(.A(new_n279_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT29), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n348_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  NOR3_X1   g150(.A1(new_n279_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G22gat), .B(G50gat), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  OR3_X1    g153(.A1(new_n351_), .A2(new_n352_), .A3(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n354_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n345_), .A2(new_n347_), .A3(new_n355_), .A4(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n338_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n346_), .A2(new_n342_), .A3(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n345_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n355_), .A2(new_n356_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n360_), .A2(KEYINPUT93), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(KEYINPUT93), .B1(new_n360_), .B2(new_n361_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n357_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n336_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n258_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n254_), .B(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT27), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n370_), .B1(new_n327_), .B2(new_n258_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n368_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n372_));
  AOI22_X1  g171(.A1(new_n369_), .A2(new_n370_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n331_), .A2(KEYINPUT102), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT102), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n375_), .B1(new_n314_), .B2(new_n330_), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n365_), .B(new_n373_), .C1(new_n374_), .C2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n367_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G227gat), .A2(G233gat), .ZN(new_n379_));
  INV_X1    g178(.A(G15gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT30), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n223_), .B(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G71gat), .B(G99gat), .ZN(new_n384_));
  INV_X1    g183(.A(G43gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n383_), .B(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n285_), .B(KEYINPUT31), .ZN(new_n388_));
  AND2_X1   g187(.A1(new_n388_), .A2(KEYINPUT84), .ZN(new_n389_));
  OR2_X1    g188(.A1(new_n387_), .A2(new_n389_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n388_), .A2(KEYINPUT84), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n387_), .B1(new_n391_), .B2(new_n389_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n373_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n395_), .A2(new_n365_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n374_), .A2(new_n376_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n397_), .A2(new_n394_), .ZN(new_n398_));
  AOI22_X1  g197(.A1(new_n378_), .A2(new_n394_), .B1(new_n396_), .B2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT67), .B(G71gat), .ZN(new_n400_));
  OR2_X1    g199(.A1(new_n400_), .A2(G78gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(G78gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G57gat), .B(G64gat), .ZN(new_n403_));
  AOI22_X1  g202(.A1(new_n401_), .A2(new_n402_), .B1(KEYINPUT11), .B2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(KEYINPUT11), .ZN(new_n405_));
  INV_X1    g204(.A(G78gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n400_), .B(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n404_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT12), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT70), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT9), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT64), .B(G85gat), .ZN(new_n414_));
  INV_X1    g213(.A(G92gat), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n413_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT65), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  OAI211_X1 g217(.A(KEYINPUT65), .B(new_n413_), .C1(new_n414_), .C2(new_n415_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(G85gat), .A2(G92gat), .ZN(new_n420_));
  AND2_X1   g219(.A1(G85gat), .A2(G92gat), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n420_), .B1(new_n421_), .B2(KEYINPUT9), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n418_), .A2(new_n419_), .A3(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G99gat), .A2(G106gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(KEYINPUT6), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT6), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n426_), .A2(G99gat), .A3(G106gat), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n425_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(G106gat), .ZN(new_n429_));
  XOR2_X1   g228(.A(KEYINPUT10), .B(G99gat), .Z(new_n430_));
  AOI21_X1  g229(.A(new_n428_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G85gat), .B(G92gat), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NOR3_X1   g235(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n425_), .A2(new_n427_), .ZN(new_n439_));
  AOI211_X1 g238(.A(new_n433_), .B(new_n434_), .C1(new_n438_), .C2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT7), .ZN(new_n441_));
  INV_X1    g240(.A(G99gat), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n441_), .A2(new_n442_), .A3(new_n429_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n426_), .B1(G99gat), .B2(G106gat), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n424_), .A2(KEYINPUT6), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n435_), .B(new_n443_), .C1(new_n444_), .C2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n434_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n432_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(KEYINPUT69), .B1(new_n440_), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n443_), .A2(new_n435_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n447_), .B1(new_n428_), .B2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(new_n433_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT69), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n446_), .A2(new_n432_), .A3(new_n447_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n452_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  AOI221_X4 g254(.A(new_n412_), .B1(new_n423_), .B2(new_n431_), .C1(new_n449_), .C2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n449_), .A2(new_n455_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n423_), .A2(new_n431_), .ZN(new_n458_));
  AOI21_X1  g257(.A(KEYINPUT70), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n411_), .B1(new_n456_), .B2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G230gat), .A2(G233gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n452_), .A2(new_n454_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n408_), .A2(new_n458_), .A3(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT12), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n458_), .A2(new_n462_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n409_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n460_), .A2(new_n461_), .A3(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT71), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n460_), .A2(new_n467_), .A3(KEYINPUT71), .A4(new_n461_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n466_), .A2(KEYINPUT68), .A3(new_n463_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n461_), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n472_), .B(new_n473_), .C1(KEYINPUT68), .C2(new_n466_), .ZN(new_n474_));
  XOR2_X1   g273(.A(G120gat), .B(G148gat), .Z(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G176gat), .B(G204gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n470_), .A2(new_n471_), .A3(new_n474_), .A4(new_n480_), .ZN(new_n481_));
  AND2_X1   g280(.A1(new_n481_), .A2(KEYINPUT73), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n481_), .A2(KEYINPUT73), .ZN(new_n483_));
  AND3_X1   g282(.A1(new_n470_), .A2(new_n471_), .A3(new_n474_), .ZN(new_n484_));
  OAI22_X1  g283(.A1(new_n482_), .A2(new_n483_), .B1(new_n484_), .B2(new_n480_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT13), .ZN(new_n486_));
  OR2_X1    g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n485_), .A2(new_n486_), .ZN(new_n488_));
  AND2_X1   g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G229gat), .A2(G233gat), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT14), .ZN(new_n492_));
  XNOR2_X1  g291(.A(KEYINPUT77), .B(G8gat), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n492_), .B1(new_n493_), .B2(G1gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT78), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G15gat), .B(G22gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G1gat), .B(G8gat), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n497_), .B(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G29gat), .B(G36gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT74), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G43gat), .B(G50gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n502_), .B(new_n503_), .ZN(new_n504_));
  AND2_X1   g303(.A1(new_n500_), .A2(new_n504_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n500_), .A2(new_n504_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n491_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n504_), .B(KEYINPUT15), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n497_), .B(new_n498_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n500_), .A2(new_n504_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n510_), .A2(new_n511_), .A3(new_n490_), .ZN(new_n512_));
  XOR2_X1   g311(.A(G113gat), .B(G141gat), .Z(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT81), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G169gat), .B(G197gat), .ZN(new_n515_));
  XOR2_X1   g314(.A(new_n514_), .B(new_n515_), .Z(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n507_), .A2(new_n512_), .A3(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n517_), .B1(new_n507_), .B2(new_n512_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n489_), .A2(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n399_), .A2(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n508_), .B1(new_n456_), .B2(new_n459_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT75), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G232gat), .A2(G233gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT34), .ZN(new_n528_));
  OAI21_X1  g327(.A(KEYINPUT76), .B1(new_n528_), .B2(KEYINPUT35), .ZN(new_n529_));
  INV_X1    g328(.A(new_n465_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n529_), .B1(new_n530_), .B2(new_n504_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n526_), .A2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n532_), .A2(KEYINPUT35), .A3(new_n528_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n528_), .A2(KEYINPUT35), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n526_), .A2(new_n534_), .A3(new_n531_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G190gat), .B(G218gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G134gat), .B(G162gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(new_n539_), .B(KEYINPUT36), .Z(new_n540_));
  NAND2_X1  g339(.A1(new_n536_), .A2(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n539_), .A2(KEYINPUT36), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n533_), .A2(new_n542_), .A3(new_n535_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT37), .ZN(new_n544_));
  AND3_X1   g343(.A1(new_n541_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n544_), .B1(new_n541_), .B2(new_n543_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G231gat), .A2(G233gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n500_), .B(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(new_n408_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n509_), .B(new_n548_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(new_n409_), .ZN(new_n552_));
  XOR2_X1   g351(.A(G127gat), .B(G155gat), .Z(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT16), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G183gat), .B(G211gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT17), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT79), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n550_), .A2(new_n552_), .A3(new_n558_), .ZN(new_n559_));
  AND2_X1   g358(.A1(new_n550_), .A2(new_n552_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT17), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n556_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  OAI211_X1 g362(.A(KEYINPUT80), .B(new_n559_), .C1(new_n560_), .C2(new_n563_), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n559_), .A2(KEYINPUT80), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n547_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n524_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n397_), .ZN(new_n570_));
  OR4_X1    g369(.A1(new_n202_), .A2(new_n569_), .A3(G1gat), .A4(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n541_), .A2(new_n543_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n399_), .A2(new_n573_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n523_), .A2(new_n567_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(G1gat), .B1(new_n576_), .B2(new_n570_), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n570_), .A2(G1gat), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n202_), .B1(new_n569_), .B2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n571_), .A2(new_n577_), .A3(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT103), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n571_), .A2(KEYINPUT103), .A3(new_n577_), .A4(new_n579_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(G1324gat));
  OR3_X1    g383(.A1(new_n569_), .A2(new_n493_), .A3(new_n373_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n398_), .A2(new_n396_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n366_), .A2(new_n395_), .ZN(new_n587_));
  AOI22_X1  g386(.A1(new_n336_), .A2(new_n366_), .B1(new_n570_), .B2(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n586_), .B1(new_n588_), .B2(new_n393_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n589_), .A2(new_n575_), .A3(new_n572_), .A4(new_n395_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT104), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(G8gat), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT39), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n590_), .A2(new_n591_), .ZN(new_n596_));
  AND3_X1   g395(.A1(new_n594_), .A2(new_n595_), .A3(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n595_), .B1(new_n594_), .B2(new_n596_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n585_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT40), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  OAI211_X1 g400(.A(KEYINPUT40), .B(new_n585_), .C1(new_n597_), .C2(new_n598_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(G1325gat));
  OAI21_X1  g402(.A(G15gat), .B1(new_n576_), .B2(new_n394_), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n604_), .B(KEYINPUT41), .Z(new_n605_));
  NAND2_X1  g404(.A1(new_n393_), .A2(new_n380_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n605_), .B1(new_n569_), .B2(new_n606_), .ZN(G1326gat));
  OAI21_X1  g406(.A(G22gat), .B1(new_n576_), .B2(new_n366_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT42), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n366_), .A2(G22gat), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n609_), .B1(new_n569_), .B2(new_n610_), .ZN(G1327gat));
  NAND3_X1  g410(.A1(new_n489_), .A2(new_n567_), .A3(new_n522_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT105), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n613_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT43), .ZN(new_n617_));
  AND3_X1   g416(.A1(new_n589_), .A2(new_n617_), .A3(new_n547_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n617_), .B1(new_n589_), .B2(new_n547_), .ZN(new_n619_));
  OAI211_X1 g418(.A(KEYINPUT44), .B(new_n616_), .C1(new_n618_), .C2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(G29gat), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n570_), .A2(new_n621_), .ZN(new_n622_));
  OR2_X1    g421(.A1(new_n545_), .A2(new_n546_), .ZN(new_n623_));
  OAI21_X1  g422(.A(KEYINPUT43), .B1(new_n399_), .B2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n589_), .A2(new_n617_), .A3(new_n547_), .ZN(new_n625_));
  AOI22_X1  g424(.A1(new_n624_), .A2(new_n625_), .B1(new_n615_), .B2(new_n614_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(KEYINPUT106), .B(KEYINPUT44), .ZN(new_n627_));
  OAI211_X1 g426(.A(new_n620_), .B(new_n622_), .C1(new_n626_), .C2(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n572_), .A2(new_n566_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n524_), .A2(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n621_), .B1(new_n630_), .B2(new_n570_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n628_), .A2(new_n631_), .ZN(G1328gat));
  OAI211_X1 g431(.A(new_n620_), .B(new_n395_), .C1(new_n626_), .C2(new_n627_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(G36gat), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n373_), .A2(G36gat), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n524_), .A2(new_n629_), .A3(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT45), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n634_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT46), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n634_), .A2(KEYINPUT46), .A3(new_n637_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(G1329gat));
  OAI21_X1  g441(.A(new_n385_), .B1(new_n630_), .B2(new_n394_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n620_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n393_), .A2(G43gat), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n643_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g446(.A(G50gat), .B1(new_n644_), .B2(new_n366_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n366_), .A2(G50gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT107), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n648_), .B1(new_n630_), .B2(new_n650_), .ZN(G1331gat));
  NAND2_X1  g450(.A1(new_n566_), .A2(new_n521_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n489_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n574_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(G57gat), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n654_), .A2(new_n655_), .A3(new_n570_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n489_), .A2(new_n522_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n589_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(new_n568_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n570_), .B1(new_n659_), .B2(KEYINPUT108), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n660_), .B1(KEYINPUT108), .B2(new_n659_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n656_), .B1(new_n661_), .B2(new_n655_), .ZN(G1332gat));
  OAI21_X1  g461(.A(G64gat), .B1(new_n654_), .B2(new_n373_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT48), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n373_), .A2(G64gat), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n664_), .B1(new_n659_), .B2(new_n665_), .ZN(G1333gat));
  OAI21_X1  g465(.A(G71gat), .B1(new_n654_), .B2(new_n394_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT49), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n394_), .A2(G71gat), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n668_), .B1(new_n659_), .B2(new_n669_), .ZN(G1334gat));
  OAI21_X1  g469(.A(G78gat), .B1(new_n654_), .B2(new_n366_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT50), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n365_), .A2(new_n406_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n672_), .B1(new_n659_), .B2(new_n673_), .ZN(G1335gat));
  AND2_X1   g473(.A1(new_n658_), .A2(new_n629_), .ZN(new_n675_));
  AOI21_X1  g474(.A(G85gat), .B1(new_n675_), .B2(new_n397_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n489_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n677_), .A2(new_n567_), .A3(new_n521_), .ZN(new_n678_));
  OAI21_X1  g477(.A(KEYINPUT109), .B1(new_n618_), .B2(new_n619_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT109), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n624_), .A2(new_n680_), .A3(new_n625_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n678_), .B1(new_n679_), .B2(new_n681_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n570_), .A2(new_n414_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n676_), .B1(new_n682_), .B2(new_n683_), .ZN(G1336gat));
  NAND3_X1  g483(.A1(new_n675_), .A2(new_n415_), .A3(new_n395_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n682_), .A2(new_n395_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n685_), .B1(new_n686_), .B2(new_n415_), .ZN(G1337gat));
  INV_X1    g486(.A(KEYINPUT51), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n675_), .A2(new_n430_), .A3(new_n393_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n682_), .A2(new_n393_), .ZN(new_n690_));
  OAI211_X1 g489(.A(new_n688_), .B(new_n689_), .C1(new_n690_), .C2(new_n442_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n442_), .B1(new_n682_), .B2(new_n393_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n689_), .ZN(new_n693_));
  OAI21_X1  g492(.A(KEYINPUT51), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n691_), .A2(new_n694_), .ZN(G1338gat));
  NAND2_X1  g494(.A1(new_n624_), .A2(new_n625_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n678_), .A2(new_n366_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n429_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  OR2_X1    g497(.A1(new_n698_), .A2(KEYINPUT52), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n366_), .A2(G106gat), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n589_), .A2(new_n629_), .A3(new_n657_), .A4(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT110), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n701_), .B(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n703_), .B1(new_n698_), .B2(KEYINPUT52), .ZN(new_n704_));
  XNOR2_X1  g503(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n699_), .A2(new_n704_), .A3(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n705_), .B1(new_n699_), .B2(new_n704_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n706_), .A2(new_n707_), .ZN(G1339gat));
  NAND2_X1  g507(.A1(new_n652_), .A2(KEYINPUT112), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT112), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n566_), .A2(new_n710_), .A3(new_n521_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n709_), .A2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT54), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n623_), .A2(new_n713_), .A3(new_n489_), .A4(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT113), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n547_), .A2(new_n712_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT113), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n717_), .A2(new_n489_), .A3(new_n718_), .A4(new_n714_), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n677_), .A2(new_n547_), .A3(new_n712_), .ZN(new_n720_));
  OAI211_X1 g519(.A(new_n716_), .B(new_n719_), .C1(new_n714_), .C2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT55), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n470_), .A2(new_n722_), .A3(new_n471_), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n440_), .A2(new_n448_), .A3(KEYINPUT69), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n453_), .B1(new_n452_), .B2(new_n454_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n458_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(new_n412_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n457_), .A2(KEYINPUT70), .A3(new_n458_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n410_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n464_), .A2(new_n466_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n473_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n460_), .A2(new_n467_), .A3(KEYINPUT55), .A4(new_n461_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n723_), .A2(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n734_), .A2(KEYINPUT56), .A3(new_n479_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT117), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n479_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT56), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT117), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n734_), .A2(new_n740_), .A3(KEYINPUT56), .A4(new_n479_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n736_), .A2(new_n739_), .A3(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n490_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n510_), .A2(new_n511_), .A3(new_n491_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n743_), .A2(new_n516_), .A3(new_n744_), .ZN(new_n745_));
  AND3_X1   g544(.A1(new_n518_), .A2(new_n745_), .A3(KEYINPUT115), .ZN(new_n746_));
  AOI21_X1  g545(.A(KEYINPUT115), .B1(new_n518_), .B2(new_n745_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n481_), .A2(KEYINPUT73), .ZN(new_n749_));
  OR2_X1    g548(.A1(new_n481_), .A2(KEYINPUT73), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n748_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT58), .ZN(new_n752_));
  AND3_X1   g551(.A1(new_n742_), .A2(new_n751_), .A3(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n742_), .B2(new_n751_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n547_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT114), .ZN(new_n756_));
  AOI21_X1  g555(.A(KEYINPUT56), .B1(new_n734_), .B2(new_n479_), .ZN(new_n757_));
  AOI211_X1 g556(.A(new_n738_), .B(new_n480_), .C1(new_n723_), .C2(new_n733_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n522_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n756_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n521_), .B1(new_n750_), .B2(new_n749_), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n762_), .B(KEYINPUT114), .C1(new_n757_), .C2(new_n758_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n748_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n485_), .A2(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n761_), .A2(new_n763_), .A3(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n766_), .A2(KEYINPUT57), .A3(new_n572_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n762_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n768_));
  AOI22_X1  g567(.A1(new_n768_), .A2(new_n756_), .B1(new_n485_), .B2(new_n764_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n573_), .B1(new_n769_), .B2(new_n763_), .ZN(new_n770_));
  XOR2_X1   g569(.A(KEYINPUT116), .B(KEYINPUT57), .Z(new_n771_));
  OAI211_X1 g570(.A(new_n755_), .B(new_n767_), .C1(new_n770_), .C2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(new_n567_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n721_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT59), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n396_), .A2(new_n397_), .A3(new_n393_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT119), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n774_), .A2(new_n775_), .A3(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n777_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT118), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n772_), .A2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n766_), .A2(new_n572_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n771_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n784_), .A2(KEYINPUT118), .A3(new_n755_), .A4(new_n767_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n781_), .A2(new_n567_), .A3(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n779_), .B1(new_n786_), .B2(new_n721_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n778_), .B1(new_n787_), .B2(new_n775_), .ZN(new_n788_));
  OAI21_X1  g587(.A(G113gat), .B1(new_n788_), .B2(new_n521_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n785_), .A2(new_n567_), .ZN(new_n790_));
  AND2_X1   g589(.A1(new_n755_), .A2(new_n767_), .ZN(new_n791_));
  AOI21_X1  g590(.A(KEYINPUT118), .B1(new_n791_), .B2(new_n784_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n721_), .B1(new_n790_), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(new_n777_), .ZN(new_n794_));
  OR2_X1    g593(.A1(new_n521_), .A2(G113gat), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n789_), .B1(new_n794_), .B2(new_n795_), .ZN(G1340gat));
  OAI21_X1  g595(.A(G120gat), .B1(new_n788_), .B2(new_n489_), .ZN(new_n797_));
  INV_X1    g596(.A(G120gat), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n798_), .B1(new_n489_), .B2(KEYINPUT60), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n799_), .B1(KEYINPUT60), .B2(new_n798_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n797_), .B1(new_n794_), .B2(new_n800_), .ZN(G1341gat));
  INV_X1    g600(.A(G127gat), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n802_), .B1(new_n794_), .B2(new_n567_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n567_), .A2(new_n802_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n803_), .B1(new_n788_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT120), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n803_), .B(KEYINPUT120), .C1(new_n788_), .C2(new_n805_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(G1342gat));
  OAI21_X1  g609(.A(G134gat), .B1(new_n788_), .B2(new_n623_), .ZN(new_n811_));
  OR2_X1    g610(.A1(new_n572_), .A2(G134gat), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n811_), .B1(new_n794_), .B2(new_n812_), .ZN(G1343gat));
  AND4_X1   g612(.A1(new_n397_), .A2(new_n793_), .A3(new_n587_), .A4(new_n394_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n522_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n815_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g615(.A1(new_n814_), .A2(new_n677_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(KEYINPUT121), .B(G148gat), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n817_), .B(new_n818_), .ZN(G1345gat));
  NAND2_X1  g618(.A1(new_n814_), .A2(new_n566_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(KEYINPUT61), .B(G155gat), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n820_), .B(new_n821_), .ZN(G1346gat));
  AOI21_X1  g621(.A(new_n393_), .B1(new_n786_), .B2(new_n721_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n823_), .A2(new_n397_), .A3(new_n587_), .ZN(new_n824_));
  OAI21_X1  g623(.A(G162gat), .B1(new_n824_), .B2(new_n623_), .ZN(new_n825_));
  OR2_X1    g624(.A1(new_n572_), .A2(G162gat), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n825_), .B1(new_n824_), .B2(new_n826_), .ZN(G1347gat));
  INV_X1    g626(.A(G169gat), .ZN(new_n828_));
  NOR3_X1   g627(.A1(new_n397_), .A2(new_n373_), .A3(new_n394_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n522_), .ZN(new_n830_));
  XOR2_X1   g629(.A(new_n830_), .B(KEYINPUT122), .Z(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n366_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n828_), .B1(new_n833_), .B2(new_n774_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n834_), .A2(KEYINPUT123), .A3(KEYINPUT62), .ZN(new_n835_));
  XNOR2_X1  g634(.A(KEYINPUT123), .B(KEYINPUT62), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n774_), .A2(new_n366_), .A3(new_n829_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n838_));
  AND2_X1   g637(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n522_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  OAI221_X1 g639(.A(new_n835_), .B1(new_n834_), .B2(new_n836_), .C1(new_n837_), .C2(new_n840_), .ZN(G1348gat));
  INV_X1    g640(.A(new_n837_), .ZN(new_n842_));
  AOI21_X1  g641(.A(G176gat), .B1(new_n842_), .B2(new_n677_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n365_), .B1(new_n786_), .B2(new_n721_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT124), .ZN(new_n845_));
  OR2_X1    g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n845_), .ZN(new_n847_));
  AND3_X1   g646(.A1(new_n846_), .A2(new_n829_), .A3(new_n847_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n677_), .A2(G176gat), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n843_), .B1(new_n848_), .B2(new_n849_), .ZN(G1349gat));
  NOR3_X1   g649(.A1(new_n837_), .A2(new_n567_), .A3(new_n212_), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n846_), .A2(new_n566_), .A3(new_n829_), .A4(new_n847_), .ZN(new_n852_));
  INV_X1    g651(.A(G183gat), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n851_), .B1(new_n852_), .B2(new_n853_), .ZN(G1350gat));
  OAI21_X1  g653(.A(G190gat), .B1(new_n837_), .B2(new_n623_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n573_), .A2(new_n213_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n855_), .B1(new_n837_), .B2(new_n856_), .ZN(G1351gat));
  NAND3_X1  g656(.A1(new_n570_), .A2(new_n365_), .A3(new_n395_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n793_), .A2(new_n394_), .A3(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(KEYINPUT125), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT125), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n823_), .A2(new_n862_), .A3(new_n859_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(G197gat), .B1(new_n864_), .B2(new_n522_), .ZN(new_n865_));
  AOI211_X1 g664(.A(new_n229_), .B(new_n521_), .C1(new_n861_), .C2(new_n863_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n865_), .A2(new_n866_), .ZN(G1352gat));
  NOR2_X1   g666(.A1(new_n860_), .A2(KEYINPUT125), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n862_), .B1(new_n823_), .B2(new_n859_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n677_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(G204gat), .ZN(new_n871_));
  INV_X1    g670(.A(G204gat), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n864_), .A2(new_n872_), .A3(new_n677_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n871_), .A2(new_n873_), .ZN(G1353gat));
  NOR2_X1   g673(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(KEYINPUT126), .ZN(new_n876_));
  NAND2_X1  g675(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n566_), .A2(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n876_), .B1(new_n864_), .B2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n878_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n876_), .ZN(new_n881_));
  AOI211_X1 g680(.A(new_n880_), .B(new_n881_), .C1(new_n861_), .C2(new_n863_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n879_), .A2(new_n882_), .ZN(G1354gat));
  NAND2_X1  g682(.A1(new_n864_), .A2(new_n573_), .ZN(new_n884_));
  XOR2_X1   g683(.A(KEYINPUT127), .B(G218gat), .Z(new_n885_));
  NOR2_X1   g684(.A1(new_n623_), .A2(new_n885_), .ZN(new_n886_));
  AOI22_X1  g685(.A1(new_n884_), .A2(new_n885_), .B1(new_n864_), .B2(new_n886_), .ZN(G1355gat));
endmodule


