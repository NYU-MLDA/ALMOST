//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 1 1 0 0 1 0 1 0 0 1 1 0 1 0 0 1 1 1 0 1 0 0 1 1 0 0 0 0 1 0 0 0 0 1 0 0 0 1 0 0 0 1 0 1 1 0 1 0 1 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n634_, new_n635_, new_n636_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n839_, new_n841_, new_n842_, new_n843_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n850_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n875_, new_n876_, new_n877_, new_n879_, new_n880_, new_n882_,
    new_n883_, new_n884_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n906_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT23), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT23), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n204_), .A2(G183gat), .A3(G190gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n206_), .B1(G183gat), .B2(G190gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT22), .B(G169gat), .ZN(new_n210_));
  INV_X1    g009(.A(G176gat), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n209_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n207_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G190gat), .ZN(new_n214_));
  OR3_X1    g013(.A1(new_n214_), .A2(KEYINPUT76), .A3(KEYINPUT26), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT25), .B(G183gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT26), .B1(new_n214_), .B2(KEYINPUT76), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT24), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220_));
  AOI22_X1  g019(.A1(new_n203_), .A2(new_n205_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n220_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n222_), .A2(KEYINPUT24), .A3(new_n208_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n218_), .A2(new_n221_), .A3(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n213_), .A2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(KEYINPUT30), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G71gat), .B(G99gat), .ZN(new_n227_));
  INV_X1    g026(.A(G43gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n227_), .B(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G227gat), .A2(G233gat), .ZN(new_n230_));
  INV_X1    g029(.A(G15gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n230_), .B(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n229_), .B(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n226_), .B(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT31), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G127gat), .B(G134gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G113gat), .B(G120gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n235_), .B(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G225gat), .A2(G233gat), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G141gat), .A2(G148gat), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT77), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT2), .ZN(new_n246_));
  NAND3_X1  g045(.A1(KEYINPUT77), .A2(G141gat), .A3(G148gat), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n245_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT79), .ZN(new_n249_));
  INV_X1    g048(.A(G141gat), .ZN(new_n250_));
  INV_X1    g049(.A(G148gat), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n249_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(KEYINPUT3), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT3), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n249_), .A2(new_n254_), .A3(new_n250_), .A4(new_n251_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n248_), .A2(new_n253_), .A3(new_n255_), .A4(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G155gat), .A2(G162gat), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(G155gat), .A2(G162gat), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n257_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n250_), .A2(new_n251_), .ZN(new_n263_));
  AND3_X1   g062(.A1(new_n245_), .A2(new_n263_), .A3(new_n247_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT78), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n258_), .A2(new_n265_), .A3(KEYINPUT1), .ZN(new_n266_));
  INV_X1    g065(.A(new_n260_), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n266_), .B(new_n267_), .C1(KEYINPUT1), .C2(new_n258_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n265_), .B1(new_n258_), .B2(KEYINPUT1), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n264_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n262_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT80), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n262_), .A2(KEYINPUT80), .A3(new_n270_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n273_), .A2(new_n239_), .A3(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(KEYINPUT86), .B1(new_n271_), .B2(new_n239_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n273_), .A2(KEYINPUT86), .A3(new_n239_), .A4(new_n274_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n242_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  AND3_X1   g078(.A1(new_n262_), .A2(KEYINPUT80), .A3(new_n270_), .ZN(new_n280_));
  AOI21_X1  g079(.A(KEYINPUT80), .B1(new_n262_), .B2(new_n270_), .ZN(new_n281_));
  NOR3_X1   g080(.A1(new_n280_), .A2(new_n281_), .A3(new_n238_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n276_), .ZN(new_n283_));
  OAI211_X1 g082(.A(KEYINPUT4), .B(new_n278_), .C1(new_n282_), .C2(new_n283_), .ZN(new_n284_));
  OR2_X1    g083(.A1(new_n275_), .A2(KEYINPUT4), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n279_), .B1(new_n286_), .B2(new_n242_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G1gat), .B(G29gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT0), .ZN(new_n289_));
  INV_X1    g088(.A(G57gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(G85gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n287_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n293_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n241_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n295_), .B1(new_n296_), .B2(new_n279_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n294_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G226gat), .A2(G233gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT19), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT26), .B(G190gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n216_), .A2(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n303_), .A2(new_n221_), .A3(new_n223_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT84), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n303_), .A2(new_n221_), .A3(KEYINPUT84), .A4(new_n223_), .ZN(new_n307_));
  AOI22_X1  g106(.A1(new_n306_), .A2(new_n307_), .B1(new_n207_), .B2(new_n212_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G197gat), .B(G204gat), .ZN(new_n309_));
  XOR2_X1   g108(.A(G211gat), .B(G218gat), .Z(new_n310_));
  INV_X1    g109(.A(KEYINPUT21), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n309_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G211gat), .B(G218gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT21), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n313_), .A2(new_n309_), .A3(KEYINPUT21), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n308_), .A2(new_n318_), .ZN(new_n319_));
  OAI21_X1  g118(.A(KEYINPUT20), .B1(new_n317_), .B2(new_n225_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n301_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n308_), .A2(new_n318_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n301_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n317_), .A2(new_n225_), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n322_), .A2(KEYINPUT20), .A3(new_n323_), .A4(new_n324_), .ZN(new_n325_));
  XOR2_X1   g124(.A(G8gat), .B(G36gat), .Z(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT18), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G64gat), .B(G92gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n321_), .A2(new_n325_), .A3(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT27), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n324_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n213_), .A2(new_n304_), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT20), .B1(new_n317_), .B2(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n301_), .B1(new_n334_), .B2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n320_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n338_), .B1(new_n318_), .B2(new_n308_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n337_), .B1(new_n339_), .B2(new_n301_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n329_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n321_), .A2(new_n325_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(new_n341_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(new_n330_), .ZN(new_n345_));
  AOI22_X1  g144(.A1(new_n333_), .A2(new_n342_), .B1(new_n345_), .B2(new_n332_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n299_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT29), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n348_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n349_));
  XOR2_X1   g148(.A(G22gat), .B(G50gat), .Z(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n269_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT1), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n260_), .B1(new_n259_), .B2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n353_), .A2(new_n355_), .A3(new_n266_), .ZN(new_n356_));
  AOI22_X1  g155(.A1(new_n257_), .A2(new_n261_), .B1(new_n356_), .B2(new_n264_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n317_), .B1(new_n357_), .B2(new_n348_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G228gat), .A2(G233gat), .ZN(new_n359_));
  XOR2_X1   g158(.A(new_n359_), .B(KEYINPUT82), .Z(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n358_), .A2(new_n361_), .ZN(new_n362_));
  NOR3_X1   g161(.A1(new_n280_), .A2(new_n281_), .A3(new_n348_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n317_), .A2(new_n360_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n362_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G78gat), .B(G106gat), .ZN(new_n366_));
  XOR2_X1   g165(.A(new_n366_), .B(KEYINPUT83), .Z(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n365_), .A2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n273_), .A2(KEYINPUT29), .A3(new_n274_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n370_), .A2(new_n317_), .A3(new_n360_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n371_), .A2(new_n367_), .A3(new_n362_), .ZN(new_n372_));
  XOR2_X1   g171(.A(KEYINPUT81), .B(KEYINPUT28), .Z(new_n373_));
  AND3_X1   g172(.A1(new_n369_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n373_), .B1(new_n369_), .B2(new_n372_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n352_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n373_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n365_), .A2(new_n368_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n367_), .B1(new_n371_), .B2(new_n362_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n377_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n369_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n380_), .A2(new_n351_), .A3(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n376_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n240_), .B1(new_n347_), .B2(new_n384_), .ZN(new_n385_));
  OAI211_X1 g184(.A(KEYINPUT33), .B(new_n295_), .C1(new_n296_), .C2(new_n279_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n242_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n241_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n293_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT85), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n329_), .B1(new_n321_), .B2(new_n325_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n390_), .B1(new_n331_), .B2(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n344_), .A2(KEYINPUT85), .A3(new_n330_), .ZN(new_n393_));
  AND4_X1   g192(.A1(new_n386_), .A2(new_n389_), .A3(new_n392_), .A4(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT87), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT33), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n395_), .B1(new_n297_), .B2(new_n396_), .ZN(new_n397_));
  AND3_X1   g196(.A1(new_n297_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n394_), .B(KEYINPUT88), .C1(new_n397_), .C2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT89), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n329_), .A2(KEYINPUT32), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n337_), .ZN(new_n403_));
  NOR3_X1   g202(.A1(new_n319_), .A2(new_n301_), .A3(new_n320_), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n400_), .B(new_n402_), .C1(new_n403_), .C2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n321_), .A2(new_n325_), .A3(new_n401_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n400_), .B1(new_n340_), .B2(new_n402_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n287_), .A2(new_n293_), .ZN(new_n410_));
  NOR3_X1   g209(.A1(new_n296_), .A2(new_n295_), .A3(new_n279_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n409_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n412_), .A2(new_n383_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n399_), .A2(new_n413_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n386_), .A2(new_n389_), .A3(new_n392_), .A4(new_n393_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n297_), .A2(new_n396_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT87), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n297_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n415_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n419_), .A2(KEYINPUT88), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n385_), .B1(new_n414_), .B2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n333_), .A2(new_n342_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n345_), .A2(new_n332_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT90), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n346_), .A2(KEYINPUT90), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n428_), .A2(new_n383_), .A3(new_n299_), .A4(new_n240_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n421_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT37), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G232gat), .A2(G233gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT34), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT35), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT6), .ZN(new_n435_));
  INV_X1    g234(.A(G99gat), .ZN(new_n436_));
  INV_X1    g235(.A(G106gat), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n435_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT7), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n439_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n441_));
  OAI21_X1  g240(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n438_), .A2(new_n440_), .A3(new_n441_), .A4(new_n442_), .ZN(new_n443_));
  XOR2_X1   g242(.A(G85gat), .B(G92gat), .Z(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT8), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT8), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n443_), .A2(new_n447_), .A3(new_n444_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n444_), .A2(KEYINPUT9), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n438_), .A2(new_n441_), .ZN(new_n451_));
  INV_X1    g250(.A(G92gat), .ZN(new_n452_));
  NOR3_X1   g251(.A1(new_n292_), .A2(new_n452_), .A3(KEYINPUT9), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n451_), .A2(new_n453_), .ZN(new_n454_));
  AND2_X1   g253(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n455_));
  NOR2_X1   g254(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  AND3_X1   g256(.A1(new_n457_), .A2(KEYINPUT64), .A3(new_n437_), .ZN(new_n458_));
  AOI21_X1  g257(.A(KEYINPUT64), .B1(new_n457_), .B2(new_n437_), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n450_), .B(new_n454_), .C1(new_n458_), .C2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n449_), .A2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G29gat), .B(G36gat), .ZN(new_n462_));
  OR2_X1    g261(.A1(new_n462_), .A2(KEYINPUT68), .ZN(new_n463_));
  INV_X1    g262(.A(G36gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(G29gat), .ZN(new_n465_));
  INV_X1    g264(.A(G29gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(G36gat), .ZN(new_n467_));
  AND3_X1   g266(.A1(new_n465_), .A2(new_n467_), .A3(KEYINPUT68), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  XOR2_X1   g268(.A(G43gat), .B(G50gat), .Z(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n463_), .A2(new_n469_), .A3(new_n471_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n462_), .A2(KEYINPUT68), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n470_), .B1(new_n473_), .B2(new_n468_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n461_), .A2(new_n475_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n433_), .A2(KEYINPUT35), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n434_), .B1(new_n478_), .B2(KEYINPUT70), .ZN(new_n479_));
  AND3_X1   g278(.A1(new_n443_), .A2(new_n447_), .A3(new_n444_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n447_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n481_));
  OAI21_X1  g280(.A(KEYINPUT67), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT67), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n446_), .A2(new_n483_), .A3(new_n448_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n482_), .A2(new_n484_), .A3(new_n460_), .ZN(new_n485_));
  XOR2_X1   g284(.A(KEYINPUT69), .B(KEYINPUT15), .Z(new_n486_));
  NOR2_X1   g285(.A1(new_n475_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n486_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n488_), .B1(new_n472_), .B2(new_n474_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n485_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n478_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n479_), .A2(new_n491_), .ZN(new_n492_));
  OAI211_X1 g291(.A(new_n478_), .B(new_n490_), .C1(KEYINPUT70), .C2(new_n434_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G190gat), .B(G218gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G134gat), .B(G162gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  XOR2_X1   g296(.A(new_n497_), .B(KEYINPUT36), .Z(new_n498_));
  XOR2_X1   g297(.A(new_n498_), .B(KEYINPUT71), .Z(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n494_), .A2(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n497_), .A2(KEYINPUT36), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n492_), .A2(new_n502_), .A3(new_n493_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n431_), .B1(new_n501_), .B2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n494_), .A2(new_n498_), .ZN(new_n505_));
  AND2_X1   g304(.A1(new_n505_), .A2(new_n503_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n504_), .B1(new_n431_), .B2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(KEYINPUT72), .B(G15gat), .ZN(new_n508_));
  INV_X1    g307(.A(G22gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G1gat), .A2(G8gat), .ZN(new_n510_));
  AOI22_X1  g309(.A1(new_n508_), .A2(new_n509_), .B1(KEYINPUT14), .B2(new_n510_), .ZN(new_n511_));
  XOR2_X1   g310(.A(KEYINPUT72), .B(G15gat), .Z(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(G22gat), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  XOR2_X1   g313(.A(G1gat), .B(G8gat), .Z(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n514_), .A2(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n511_), .A2(new_n513_), .A3(new_n515_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G231gat), .A2(G233gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G57gat), .B(G64gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G71gat), .B(G78gat), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n522_), .A2(new_n523_), .A3(KEYINPUT11), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(KEYINPUT11), .ZN(new_n525_));
  INV_X1    g324(.A(new_n523_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n522_), .A2(KEYINPUT11), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n524_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n521_), .B(new_n529_), .ZN(new_n530_));
  XOR2_X1   g329(.A(G127gat), .B(G155gat), .Z(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT16), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G183gat), .B(G211gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT17), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  AND2_X1   g335(.A1(new_n534_), .A2(new_n535_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n530_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n538_), .B1(new_n536_), .B2(new_n530_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT73), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT73), .ZN(new_n541_));
  OAI211_X1 g340(.A(new_n538_), .B(new_n541_), .C1(new_n536_), .C2(new_n530_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n507_), .A2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G120gat), .B(G148gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT5), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G176gat), .B(G204gat), .ZN(new_n547_));
  XOR2_X1   g346(.A(new_n546_), .B(new_n547_), .Z(new_n548_));
  OAI211_X1 g347(.A(new_n460_), .B(new_n529_), .C1(new_n481_), .C2(new_n480_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT65), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n529_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n461_), .A2(new_n552_), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n449_), .A2(KEYINPUT65), .A3(new_n460_), .A4(new_n529_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n551_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT66), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G230gat), .A2(G233gat), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n555_), .A2(new_n556_), .A3(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n549_), .A2(KEYINPUT12), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(new_n553_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n485_), .A2(KEYINPUT12), .A3(new_n552_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n561_), .A2(new_n562_), .A3(new_n557_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n559_), .A2(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n556_), .B1(new_n555_), .B2(new_n558_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n548_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n565_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n548_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n567_), .A2(new_n559_), .A3(new_n563_), .A4(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n566_), .A2(new_n569_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n570_), .A2(KEYINPUT13), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n570_), .A2(KEYINPUT13), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n518_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n515_), .B1(new_n511_), .B2(new_n513_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n475_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n517_), .A2(new_n472_), .A3(new_n518_), .A4(new_n474_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT74), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n576_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G229gat), .A2(G233gat), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n519_), .A2(KEYINPUT74), .A3(new_n475_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n579_), .A2(new_n581_), .A3(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT75), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n579_), .A2(KEYINPUT75), .A3(new_n581_), .A4(new_n582_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n519_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n587_), .A2(new_n580_), .A3(new_n577_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n585_), .A2(new_n586_), .A3(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G113gat), .B(G141gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G169gat), .B(G197gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n589_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n592_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n585_), .A2(new_n588_), .A3(new_n586_), .A4(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n573_), .A2(new_n597_), .ZN(new_n598_));
  AND3_X1   g397(.A1(new_n430_), .A2(new_n544_), .A3(new_n598_), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n599_), .A2(KEYINPUT91), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(KEYINPUT91), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n299_), .A2(G1gat), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n600_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT92), .ZN(new_n604_));
  OR2_X1    g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n603_), .A2(new_n604_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT38), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n605_), .A2(KEYINPUT38), .A3(new_n606_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n506_), .B1(new_n421_), .B2(new_n429_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n543_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n598_), .B(KEYINPUT93), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n611_), .A2(new_n612_), .A3(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(G1gat), .B1(new_n614_), .B2(new_n299_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT94), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n609_), .A2(new_n610_), .A3(new_n616_), .ZN(G1324gat));
  OAI21_X1  g416(.A(G8gat), .B1(new_n614_), .B2(new_n428_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(KEYINPUT95), .B(KEYINPUT39), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n428_), .A2(G8gat), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n600_), .A2(new_n601_), .A3(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n618_), .A2(new_n619_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n620_), .A2(new_n622_), .A3(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(KEYINPUT96), .B(KEYINPUT40), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(G1325gat));
  XNOR2_X1  g425(.A(new_n235_), .B(new_n238_), .ZN(new_n627_));
  OAI21_X1  g426(.A(G15gat), .B1(new_n614_), .B2(new_n627_), .ZN(new_n628_));
  XOR2_X1   g427(.A(KEYINPUT97), .B(KEYINPUT41), .Z(new_n629_));
  OR2_X1    g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(new_n629_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n599_), .A2(new_n231_), .A3(new_n240_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n630_), .A2(new_n631_), .A3(new_n632_), .ZN(G1326gat));
  OAI21_X1  g432(.A(G22gat), .B1(new_n614_), .B2(new_n383_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT42), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n599_), .A2(new_n509_), .A3(new_n384_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(G1327gat));
  NAND2_X1  g436(.A1(new_n505_), .A2(new_n503_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n612_), .A2(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n424_), .A2(new_n298_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n627_), .B1(new_n640_), .B2(new_n383_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n412_), .A2(new_n383_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n642_), .B1(new_n419_), .B2(KEYINPUT88), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT88), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n398_), .A2(new_n397_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n644_), .B1(new_n645_), .B2(new_n415_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n641_), .B1(new_n643_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n429_), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n598_), .B(new_n639_), .C1(new_n647_), .C2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(KEYINPUT99), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT99), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n430_), .A2(new_n651_), .A3(new_n598_), .A4(new_n639_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(G29gat), .B1(new_n654_), .B2(new_n298_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n613_), .A2(new_n543_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n504_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n505_), .A2(new_n431_), .A3(new_n503_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n657_), .A2(KEYINPUT98), .A3(new_n658_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n659_), .A2(KEYINPUT43), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n661_), .B1(new_n430_), .B2(new_n507_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n657_), .A2(new_n658_), .ZN(new_n663_));
  AOI211_X1 g462(.A(new_n663_), .B(new_n660_), .C1(new_n421_), .C2(new_n429_), .ZN(new_n664_));
  OAI211_X1 g463(.A(new_n656_), .B(KEYINPUT44), .C1(new_n662_), .C2(new_n664_), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n665_), .A2(G29gat), .A3(new_n298_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n656_), .B1(new_n662_), .B2(new_n664_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT44), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n655_), .B1(new_n666_), .B2(new_n669_), .ZN(G1328gat));
  INV_X1    g469(.A(new_n428_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n669_), .A2(new_n671_), .A3(new_n665_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n428_), .A2(G36gat), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n650_), .A2(new_n652_), .A3(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(KEYINPUT101), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT101), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n650_), .A2(new_n652_), .A3(new_n676_), .A4(new_n673_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(new_n678_));
  XOR2_X1   g477(.A(KEYINPUT100), .B(KEYINPUT45), .Z(new_n679_));
  AOI22_X1  g478(.A1(new_n672_), .A2(G36gat), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n679_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n675_), .A2(new_n677_), .A3(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT102), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n683_), .A2(KEYINPUT46), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n682_), .A2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n683_), .A2(KEYINPUT46), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n680_), .A2(new_n685_), .A3(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n686_), .B1(new_n680_), .B2(new_n685_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1329gat));
  NAND4_X1  g488(.A1(new_n669_), .A2(G43gat), .A3(new_n240_), .A4(new_n665_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n228_), .B1(new_n653_), .B2(new_n627_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  XOR2_X1   g491(.A(KEYINPUT103), .B(KEYINPUT47), .Z(new_n693_));
  XNOR2_X1  g492(.A(new_n692_), .B(new_n693_), .ZN(G1330gat));
  AND3_X1   g493(.A1(new_n669_), .A2(new_n384_), .A3(new_n665_), .ZN(new_n695_));
  INV_X1    g494(.A(G50gat), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n384_), .A2(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT104), .ZN(new_n698_));
  OAI22_X1  g497(.A1(new_n695_), .A2(new_n696_), .B1(new_n653_), .B2(new_n698_), .ZN(G1331gat));
  INV_X1    g498(.A(new_n573_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n700_), .A2(new_n596_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n611_), .A2(new_n612_), .A3(new_n701_), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n702_), .A2(new_n290_), .A3(new_n299_), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT105), .Z(new_n704_));
  AND2_X1   g503(.A1(new_n430_), .A2(new_n701_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n705_), .A2(new_n544_), .ZN(new_n706_));
  AOI21_X1  g505(.A(G57gat), .B1(new_n706_), .B2(new_n298_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n704_), .A2(new_n707_), .ZN(G1332gat));
  OAI21_X1  g507(.A(G64gat), .B1(new_n702_), .B2(new_n428_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT48), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n428_), .A2(G64gat), .ZN(new_n711_));
  XOR2_X1   g510(.A(new_n711_), .B(KEYINPUT106), .Z(new_n712_));
  NAND2_X1  g511(.A1(new_n706_), .A2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n710_), .A2(new_n713_), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT107), .Z(G1333gat));
  OAI21_X1  g514(.A(G71gat), .B1(new_n702_), .B2(new_n627_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT49), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n627_), .A2(G71gat), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT108), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n706_), .A2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n717_), .A2(new_n720_), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT109), .Z(G1334gat));
  OAI21_X1  g521(.A(G78gat), .B1(new_n702_), .B2(new_n383_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT50), .ZN(new_n724_));
  INV_X1    g523(.A(G78gat), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n706_), .A2(new_n725_), .A3(new_n384_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(G1335gat));
  AND2_X1   g526(.A1(new_n705_), .A2(new_n639_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n728_), .A2(new_n292_), .A3(new_n298_), .ZN(new_n729_));
  NOR3_X1   g528(.A1(new_n700_), .A2(new_n612_), .A3(new_n596_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n730_), .B1(new_n662_), .B2(new_n664_), .ZN(new_n731_));
  OR2_X1    g530(.A1(new_n731_), .A2(KEYINPUT110), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(KEYINPUT110), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n299_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n729_), .B1(new_n734_), .B2(new_n292_), .ZN(G1336gat));
  NAND3_X1  g534(.A1(new_n728_), .A2(new_n452_), .A3(new_n671_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n428_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n736_), .B1(new_n737_), .B2(new_n452_), .ZN(G1337gat));
  NAND3_X1  g537(.A1(new_n728_), .A2(new_n457_), .A3(new_n240_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n627_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n739_), .B1(new_n740_), .B2(new_n436_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT111), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n741_), .A2(new_n742_), .A3(KEYINPUT51), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(KEYINPUT51), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n739_), .B(new_n744_), .C1(new_n740_), .C2(new_n436_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1338gat));
  OAI211_X1 g545(.A(new_n384_), .B(new_n730_), .C1(new_n662_), .C2(new_n664_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT52), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n747_), .A2(new_n748_), .A3(G106gat), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT112), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n747_), .A2(KEYINPUT112), .A3(new_n748_), .A4(G106gat), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n747_), .A2(G106gat), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(KEYINPUT52), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n751_), .A2(new_n752_), .A3(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n728_), .A2(new_n437_), .A3(new_n384_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(KEYINPUT53), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT53), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n755_), .A2(new_n759_), .A3(new_n756_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(G1339gat));
  INV_X1    g560(.A(KEYINPUT55), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n563_), .A2(new_n762_), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n561_), .A2(new_n562_), .A3(KEYINPUT55), .A4(new_n557_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n561_), .A2(new_n562_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(new_n558_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n763_), .A2(new_n764_), .A3(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(new_n548_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT56), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n767_), .A2(KEYINPUT56), .A3(new_n548_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n587_), .A2(new_n581_), .A3(new_n577_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n579_), .A2(new_n580_), .A3(new_n582_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n773_), .A2(new_n774_), .A3(new_n592_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n595_), .A2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(KEYINPUT113), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT113), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n595_), .A2(new_n778_), .A3(new_n775_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n772_), .A2(KEYINPUT114), .A3(new_n569_), .A4(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(KEYINPUT58), .B1(new_n781_), .B2(KEYINPUT115), .ZN(new_n782_));
  INV_X1    g581(.A(new_n569_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n783_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(KEYINPUT115), .A2(KEYINPUT58), .ZN(new_n785_));
  AOI22_X1  g584(.A1(new_n784_), .A2(new_n780_), .B1(KEYINPUT114), .B2(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n507_), .B1(new_n782_), .B2(new_n786_), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n767_), .A2(KEYINPUT56), .A3(new_n548_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT56), .B1(new_n767_), .B2(new_n548_), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n596_), .B(new_n569_), .C1(new_n788_), .C2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n779_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n778_), .B1(new_n595_), .B2(new_n775_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n570_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n790_), .A2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(KEYINPUT57), .B1(new_n794_), .B2(new_n638_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT57), .ZN(new_n796_));
  AOI211_X1 g595(.A(new_n796_), .B(new_n506_), .C1(new_n790_), .C2(new_n793_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n795_), .A2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n612_), .B1(new_n787_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT54), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n663_), .A2(new_n612_), .A3(new_n597_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n800_), .B1(new_n801_), .B2(new_n573_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n544_), .A2(KEYINPUT54), .A3(new_n597_), .A4(new_n700_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n799_), .A2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n428_), .A2(new_n298_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n240_), .A2(new_n383_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n805_), .A2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(G113gat), .B1(new_n810_), .B2(new_n596_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT59), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n812_), .B(new_n808_), .C1(new_n799_), .C2(new_n804_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT116), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n813_), .B(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(KEYINPUT59), .B1(new_n805_), .B2(new_n809_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  XOR2_X1   g617(.A(KEYINPUT117), .B(G113gat), .Z(new_n819_));
  NOR2_X1   g618(.A1(new_n597_), .A2(new_n819_), .ZN(new_n820_));
  XOR2_X1   g619(.A(new_n820_), .B(KEYINPUT118), .Z(new_n821_));
  AOI21_X1  g620(.A(new_n811_), .B1(new_n818_), .B2(new_n821_), .ZN(G1340gat));
  INV_X1    g621(.A(KEYINPUT60), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(new_n700_), .B2(G120gat), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n810_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n823_), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n813_), .A2(new_n814_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n813_), .A2(new_n814_), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n573_), .B(new_n816_), .C1(new_n828_), .C2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT119), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n815_), .A2(KEYINPUT119), .A3(new_n573_), .A4(new_n816_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n826_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(G120gat), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n827_), .B1(new_n834_), .B2(new_n835_), .ZN(G1341gat));
  NAND3_X1  g635(.A1(new_n818_), .A2(G127gat), .A3(new_n612_), .ZN(new_n837_));
  AOI21_X1  g636(.A(G127gat), .B1(new_n810_), .B2(new_n612_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(KEYINPUT120), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n837_), .A2(new_n839_), .ZN(G1342gat));
  OAI21_X1  g639(.A(G134gat), .B1(new_n817_), .B2(new_n663_), .ZN(new_n841_));
  INV_X1    g640(.A(G134gat), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n810_), .A2(new_n842_), .A3(new_n506_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n843_), .ZN(G1343gat));
  NOR3_X1   g643(.A1(new_n805_), .A2(new_n383_), .A3(new_n240_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n806_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n847_), .A2(new_n597_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n848_), .B(new_n250_), .ZN(G1344gat));
  NOR2_X1   g648(.A1(new_n847_), .A2(new_n700_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(new_n251_), .ZN(G1345gat));
  INV_X1    g650(.A(KEYINPUT121), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n852_), .B1(new_n847_), .B2(new_n543_), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n845_), .A2(KEYINPUT121), .A3(new_n612_), .A4(new_n846_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(KEYINPUT61), .B(G155gat), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n855_), .B(new_n856_), .ZN(G1346gat));
  OAI21_X1  g656(.A(G162gat), .B1(new_n847_), .B2(new_n663_), .ZN(new_n858_));
  OR2_X1    g657(.A1(new_n638_), .A2(G162gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n847_), .B2(new_n859_), .ZN(G1347gat));
  INV_X1    g659(.A(G169gat), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n428_), .A2(new_n298_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n863_), .A2(new_n807_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n805_), .A2(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n861_), .B1(new_n866_), .B2(new_n596_), .ZN(new_n867_));
  XOR2_X1   g666(.A(new_n867_), .B(KEYINPUT62), .Z(new_n868_));
  NAND2_X1  g667(.A1(new_n866_), .A2(KEYINPUT122), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT122), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n870_), .B1(new_n805_), .B2(new_n865_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n871_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n872_), .A2(new_n596_), .A3(new_n210_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n868_), .A2(new_n873_), .ZN(G1348gat));
  NAND3_X1  g673(.A1(new_n866_), .A2(G176gat), .A3(new_n573_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n700_), .B1(new_n869_), .B2(new_n871_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(new_n876_), .B2(G176gat), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(KEYINPUT123), .ZN(G1349gat));
  AOI21_X1  g677(.A(G183gat), .B1(new_n866_), .B2(new_n612_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n543_), .A2(new_n216_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n879_), .B1(new_n872_), .B2(new_n880_), .ZN(G1350gat));
  INV_X1    g680(.A(new_n872_), .ZN(new_n882_));
  OAI21_X1  g681(.A(G190gat), .B1(new_n882_), .B2(new_n663_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n872_), .A2(new_n506_), .A3(new_n302_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(G1351gat));
  NOR2_X1   g684(.A1(new_n240_), .A2(new_n383_), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n886_), .B(new_n862_), .C1(new_n799_), .C2(new_n804_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(KEYINPUT124), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n888_), .A2(new_n597_), .ZN(new_n889_));
  OAI21_X1  g688(.A(KEYINPUT125), .B1(new_n889_), .B2(G197gat), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT125), .ZN(new_n891_));
  INV_X1    g690(.A(G197gat), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n891_), .B(new_n892_), .C1(new_n888_), .C2(new_n597_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n889_), .A2(G197gat), .ZN(new_n894_));
  AND3_X1   g693(.A1(new_n890_), .A2(new_n893_), .A3(new_n894_), .ZN(G1352gat));
  INV_X1    g694(.A(new_n888_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n573_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g697(.A1(new_n888_), .A2(new_n543_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n900_));
  AND2_X1   g699(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n899_), .B1(new_n900_), .B2(new_n901_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n902_), .B1(new_n899_), .B2(new_n900_), .ZN(G1354gat));
  XOR2_X1   g702(.A(KEYINPUT126), .B(G218gat), .Z(new_n904_));
  NOR3_X1   g703(.A1(new_n888_), .A2(new_n663_), .A3(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n896_), .A2(new_n506_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n905_), .B1(new_n906_), .B2(new_n904_), .ZN(G1355gat));
endmodule


