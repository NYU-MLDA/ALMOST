//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 1 1 1 0 0 0 0 1 0 1 1 0 1 0 0 1 0 1 1 0 1 0 1 0 0 0 0 0 0 1 0 1 1 1 0 1 1 0 0 0 0 0 0 1 0 0 1 0 0 1 1 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n619_, new_n620_, new_n621_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n701_, new_n702_, new_n703_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n722_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n868_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n906_,
    new_n907_, new_n909_, new_n910_, new_n911_, new_n912_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_, new_n924_;
  AND2_X1   g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G85gat), .A2(G92gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  NOR2_X1   g003(.A1(G85gat), .A2(G92gat), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  OR3_X1    g005(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT6), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n208_), .B1(G99gat), .B2(G106gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n210_), .A2(KEYINPUT6), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n207_), .B1(new_n209_), .B2(new_n211_), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT66), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT66), .ZN(new_n215_));
  OAI211_X1 g014(.A(new_n215_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n206_), .B1(new_n212_), .B2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT8), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n210_), .A2(KEYINPUT6), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n208_), .A2(G99gat), .A3(G106gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n222_), .A2(new_n207_), .A3(new_n214_), .A4(new_n216_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT8), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n223_), .A2(new_n224_), .A3(new_n206_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n205_), .B1(new_n204_), .B2(KEYINPUT9), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT9), .ZN(new_n227_));
  AND3_X1   g026(.A1(new_n203_), .A2(KEYINPUT65), .A3(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(KEYINPUT65), .B1(new_n203_), .B2(new_n227_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n226_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  OR2_X1    g029(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT64), .ZN(new_n232_));
  NAND2_X1  g031(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n231_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  AND2_X1   g033(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n235_));
  NOR2_X1   g034(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT64), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n234_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(G106gat), .ZN(new_n239_));
  AOI22_X1  g038(.A1(new_n238_), .A2(new_n239_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n240_));
  AOI22_X1  g039(.A1(new_n219_), .A2(new_n225_), .B1(new_n230_), .B2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G57gat), .B(G64gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT11), .ZN(new_n243_));
  XOR2_X1   g042(.A(G71gat), .B(G78gat), .Z(new_n244_));
  OR2_X1    g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n244_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n242_), .A2(KEYINPUT11), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n245_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n241_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n241_), .A2(new_n248_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n202_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT12), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n253_), .B1(new_n241_), .B2(new_n248_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n202_), .B1(new_n241_), .B2(new_n248_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT67), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n223_), .A2(new_n224_), .A3(new_n206_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n224_), .B1(new_n223_), .B2(new_n206_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n256_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n219_), .A2(KEYINPUT67), .A3(new_n225_), .ZN(new_n260_));
  AOI22_X1  g059(.A1(new_n259_), .A2(new_n260_), .B1(new_n230_), .B2(new_n240_), .ZN(new_n261_));
  OR2_X1    g060(.A1(new_n248_), .A2(new_n253_), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n254_), .B(new_n255_), .C1(new_n261_), .C2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n252_), .A2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G120gat), .B(G148gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT5), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G176gat), .B(G204gat), .ZN(new_n267_));
  XOR2_X1   g066(.A(new_n266_), .B(new_n267_), .Z(new_n268_));
  NAND2_X1  g067(.A1(new_n264_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n268_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n252_), .A2(new_n263_), .A3(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT13), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT13), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n272_), .A2(new_n275_), .ZN(new_n276_));
  AND2_X1   g075(.A1(new_n274_), .A2(new_n276_), .ZN(new_n277_));
  OR2_X1    g076(.A1(new_n277_), .A2(KEYINPUT68), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(KEYINPUT68), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G113gat), .B(G141gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G169gat), .B(G197gat), .ZN(new_n282_));
  XOR2_X1   g081(.A(new_n281_), .B(new_n282_), .Z(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(KEYINPUT74), .B(G1gat), .ZN(new_n285_));
  INV_X1    g084(.A(G8gat), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT14), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G15gat), .B(G22gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT75), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G1gat), .B(G8gat), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n290_), .B(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G43gat), .B(G50gat), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(G36gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(G29gat), .ZN(new_n297_));
  INV_X1    g096(.A(G29gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(G36gat), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n297_), .A2(new_n299_), .A3(KEYINPUT69), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(KEYINPUT69), .B1(new_n297_), .B2(new_n299_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n295_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n297_), .A2(new_n299_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT69), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n306_), .A2(new_n300_), .A3(new_n294_), .ZN(new_n307_));
  AND3_X1   g106(.A1(new_n303_), .A2(new_n307_), .A3(KEYINPUT15), .ZN(new_n308_));
  AOI21_X1  g107(.A(KEYINPUT15), .B1(new_n303_), .B2(new_n307_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n293_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n290_), .B(new_n291_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n303_), .A2(new_n307_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT78), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n311_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G229gat), .A2(G233gat), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n310_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n293_), .A2(new_n313_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n316_), .B1(new_n315_), .B2(new_n319_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n284_), .B1(new_n318_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n320_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n322_), .A2(new_n317_), .A3(new_n283_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n321_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n280_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT33), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G225gat), .A2(G233gat), .ZN(new_n327_));
  XOR2_X1   g126(.A(new_n327_), .B(KEYINPUT91), .Z(new_n328_));
  XOR2_X1   g127(.A(new_n328_), .B(KEYINPUT92), .Z(new_n329_));
  XOR2_X1   g128(.A(G127gat), .B(G134gat), .Z(new_n330_));
  XOR2_X1   g129(.A(G113gat), .B(G120gat), .Z(new_n331_));
  XOR2_X1   g130(.A(new_n330_), .B(new_n331_), .Z(new_n332_));
  INV_X1    g131(.A(KEYINPUT2), .ZN(new_n333_));
  INV_X1    g132(.A(G141gat), .ZN(new_n334_));
  INV_X1    g133(.A(G148gat), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n333_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT3), .ZN(new_n338_));
  NOR2_X1   g137(.A1(G141gat), .A2(G148gat), .ZN(new_n339_));
  OAI211_X1 g138(.A(new_n336_), .B(new_n337_), .C1(new_n338_), .C2(new_n339_), .ZN(new_n340_));
  NOR3_X1   g139(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n341_));
  OR2_X1    g140(.A1(new_n341_), .A2(KEYINPUT83), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(KEYINPUT83), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n340_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G155gat), .A2(G162gat), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(G155gat), .A2(G162gat), .ZN(new_n347_));
  NOR3_X1   g146(.A1(new_n344_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n348_));
  AND2_X1   g147(.A1(new_n345_), .A2(KEYINPUT1), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n345_), .A2(KEYINPUT1), .ZN(new_n350_));
  NOR3_X1   g149(.A1(new_n349_), .A2(new_n350_), .A3(new_n347_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n334_), .A2(new_n335_), .ZN(new_n352_));
  NOR3_X1   g151(.A1(new_n351_), .A2(new_n339_), .A3(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n332_), .B1(new_n348_), .B2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n329_), .B1(new_n354_), .B2(KEYINPUT4), .ZN(new_n355_));
  OR3_X1    g154(.A1(new_n344_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n332_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n353_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n356_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n359_), .A2(KEYINPUT4), .A3(new_n354_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT90), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n359_), .A2(new_n354_), .A3(KEYINPUT90), .A4(KEYINPUT4), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n355_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n359_), .A2(new_n354_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n328_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n364_), .A2(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G1gat), .B(G29gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(G85gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT0), .B(G57gat), .ZN(new_n372_));
  XOR2_X1   g171(.A(new_n371_), .B(new_n372_), .Z(new_n373_));
  AOI21_X1  g172(.A(new_n326_), .B1(new_n369_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n373_), .ZN(new_n375_));
  NOR4_X1   g174(.A1(new_n364_), .A2(new_n368_), .A3(KEYINPUT33), .A4(new_n375_), .ZN(new_n376_));
  XOR2_X1   g175(.A(G8gat), .B(G36gat), .Z(new_n377_));
  XNOR2_X1  g176(.A(G64gat), .B(G92gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT88), .B(KEYINPUT18), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G183gat), .A2(G190gat), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n383_), .A2(KEYINPUT23), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT79), .B(KEYINPUT23), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n384_), .B1(new_n385_), .B2(new_n383_), .ZN(new_n386_));
  OR2_X1    g185(.A1(G169gat), .A2(G176gat), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n387_), .A2(KEYINPUT24), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  OR2_X1    g188(.A1(new_n389_), .A2(KEYINPUT80), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(KEYINPUT80), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT25), .B(G183gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT26), .B(G190gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G169gat), .A2(G176gat), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n394_), .A2(KEYINPUT24), .ZN(new_n395_));
  AOI22_X1  g194(.A1(new_n392_), .A2(new_n393_), .B1(new_n395_), .B2(new_n387_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n390_), .A2(new_n391_), .A3(new_n396_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(G169gat), .ZN(new_n399_));
  INV_X1    g198(.A(new_n383_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n385_), .A2(new_n400_), .ZN(new_n401_));
  OR2_X1    g200(.A1(new_n400_), .A2(KEYINPUT23), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(G183gat), .A2(G190gat), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n399_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n397_), .A2(new_n405_), .ZN(new_n406_));
  XOR2_X1   g205(.A(G197gat), .B(G204gat), .Z(new_n407_));
  OR2_X1    g206(.A1(new_n407_), .A2(KEYINPUT21), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(KEYINPUT21), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G211gat), .B(G218gat), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n408_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n411_));
  OR2_X1    g210(.A1(new_n409_), .A2(new_n410_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n406_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G226gat), .A2(G233gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT19), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  OR3_X1    g216(.A1(new_n403_), .A2(KEYINPUT86), .A3(new_n388_), .ZN(new_n418_));
  OAI21_X1  g217(.A(KEYINPUT86), .B1(new_n403_), .B2(new_n388_), .ZN(new_n419_));
  OR2_X1    g218(.A1(new_n396_), .A2(KEYINPUT85), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n396_), .A2(KEYINPUT85), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n418_), .A2(new_n419_), .A3(new_n420_), .A4(new_n421_), .ZN(new_n422_));
  XOR2_X1   g221(.A(KEYINPUT22), .B(G169gat), .Z(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT87), .ZN(new_n424_));
  OAI221_X1 g223(.A(new_n394_), .B1(new_n386_), .B2(new_n404_), .C1(new_n424_), .C2(G176gat), .ZN(new_n425_));
  INV_X1    g224(.A(new_n413_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n422_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n414_), .A2(KEYINPUT20), .A3(new_n417_), .A4(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT20), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n422_), .A2(new_n425_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n429_), .B1(new_n430_), .B2(new_n413_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n397_), .A2(new_n426_), .A3(new_n405_), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n382_), .B(new_n428_), .C1(new_n433_), .C2(new_n417_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n428_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n417_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n381_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n434_), .A2(new_n437_), .ZN(new_n438_));
  OAI22_X1  g237(.A1(new_n374_), .A2(new_n376_), .B1(new_n438_), .B2(KEYINPUT89), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(KEYINPUT89), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n362_), .A2(new_n363_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n354_), .A2(KEYINPUT4), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n442_), .A2(new_n328_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n441_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(KEYINPUT93), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT93), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n441_), .A2(new_n446_), .A3(new_n443_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n373_), .B1(new_n365_), .B2(new_n329_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n445_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n440_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n364_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n451_), .A2(new_n367_), .A3(new_n373_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n375_), .B1(new_n364_), .B2(new_n368_), .ZN(new_n453_));
  AND2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n433_), .A2(new_n417_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n414_), .A2(KEYINPUT20), .A3(new_n427_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(new_n416_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n435_), .A2(new_n436_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n382_), .A2(KEYINPUT32), .ZN(new_n460_));
  MUX2_X1   g259(.A(new_n458_), .B(new_n459_), .S(new_n460_), .Z(new_n461_));
  OAI22_X1  g260(.A1(new_n439_), .A2(new_n450_), .B1(new_n454_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT84), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT29), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n356_), .A2(new_n464_), .A3(new_n358_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT28), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n348_), .A2(new_n353_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT28), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n467_), .A2(new_n468_), .A3(new_n464_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G22gat), .B(G50gat), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n466_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n470_), .B1(new_n466_), .B2(new_n469_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n463_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n413_), .B1(new_n467_), .B2(new_n464_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G228gat), .A2(G233gat), .ZN(new_n476_));
  INV_X1    g275(.A(G78gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(G106gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n475_), .B(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n466_), .A2(new_n469_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n470_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n484_), .A2(KEYINPUT84), .A3(new_n471_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n474_), .A2(new_n481_), .A3(new_n485_), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n480_), .A2(KEYINPUT84), .A3(new_n471_), .A4(new_n484_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n462_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n458_), .A2(new_n381_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT94), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n490_), .A2(new_n491_), .A3(KEYINPUT27), .A4(new_n434_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT27), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n438_), .A2(new_n493_), .ZN(new_n494_));
  AND2_X1   g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT95), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n434_), .A2(KEYINPUT27), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n382_), .B1(new_n455_), .B2(new_n457_), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT94), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  AND4_X1   g298(.A1(new_n453_), .A2(new_n486_), .A3(new_n452_), .A4(new_n487_), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n495_), .A2(new_n496_), .A3(new_n499_), .A4(new_n500_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n500_), .A2(new_n499_), .A3(new_n492_), .A4(new_n494_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT95), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n489_), .A2(new_n501_), .A3(new_n503_), .ZN(new_n504_));
  XOR2_X1   g303(.A(KEYINPUT82), .B(G15gat), .Z(new_n505_));
  NAND2_X1  g304(.A1(G227gat), .A2(G233gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(KEYINPUT81), .B(G43gat), .ZN(new_n508_));
  XOR2_X1   g307(.A(new_n507_), .B(new_n508_), .Z(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(new_n332_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  XOR2_X1   g310(.A(new_n406_), .B(KEYINPUT30), .Z(new_n512_));
  XNOR2_X1  g311(.A(G71gat), .B(G99gat), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n406_), .B(KEYINPUT30), .ZN(new_n515_));
  INV_X1    g314(.A(new_n513_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT31), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n514_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n518_), .B1(new_n514_), .B2(new_n517_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n511_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n521_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n523_), .A2(new_n519_), .A3(new_n510_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n504_), .A2(new_n525_), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n492_), .A2(new_n499_), .A3(new_n494_), .A4(new_n488_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT96), .ZN(new_n528_));
  OR2_X1    g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n525_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n529_), .A2(new_n530_), .A3(new_n454_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n325_), .B1(new_n526_), .B2(new_n531_), .ZN(new_n532_));
  XOR2_X1   g331(.A(G127gat), .B(G155gat), .Z(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G183gat), .B(G211gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G231gat), .A2(G233gat), .ZN(new_n538_));
  XOR2_X1   g337(.A(new_n248_), .B(new_n538_), .Z(new_n539_));
  XNOR2_X1  g338(.A(new_n293_), .B(new_n539_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n537_), .B1(new_n540_), .B2(KEYINPUT17), .ZN(new_n541_));
  OR2_X1    g340(.A1(new_n537_), .A2(KEYINPUT17), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n540_), .A2(KEYINPUT77), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G232gat), .A2(G233gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT34), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT35), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n308_), .A2(new_n309_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n259_), .A2(new_n260_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n240_), .A2(new_n230_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n551_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n553_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n555_));
  OAI22_X1  g354(.A1(new_n555_), .A2(new_n312_), .B1(KEYINPUT35), .B2(new_n547_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n550_), .B1(new_n554_), .B2(new_n556_), .ZN(new_n557_));
  XOR2_X1   g356(.A(G190gat), .B(G218gat), .Z(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT70), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G134gat), .B(G162gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT36), .ZN(new_n562_));
  AND2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n312_), .ZN(new_n564_));
  AOI22_X1  g363(.A1(new_n241_), .A2(new_n564_), .B1(new_n549_), .B2(new_n548_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n550_), .ZN(new_n566_));
  OAI211_X1 g365(.A(new_n565_), .B(new_n566_), .C1(new_n261_), .C2(new_n551_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n557_), .A2(new_n563_), .A3(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(KEYINPUT71), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT71), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n557_), .A2(new_n570_), .A3(new_n563_), .A4(new_n567_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT37), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n557_), .A2(new_n567_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n561_), .B(KEYINPUT36), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n572_), .A2(new_n573_), .A3(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT73), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n575_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n580_), .B1(new_n557_), .B2(new_n567_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n581_), .B1(new_n569_), .B2(new_n571_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n582_), .A2(KEYINPUT73), .A3(new_n573_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n579_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n576_), .A2(KEYINPUT72), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT72), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n581_), .A2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n572_), .A2(new_n585_), .A3(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n588_), .A2(KEYINPUT37), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n545_), .B1(new_n584_), .B2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n532_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT97), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n532_), .A2(KEYINPUT97), .A3(new_n590_), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n454_), .B(KEYINPUT98), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n595_), .A2(new_n285_), .A3(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT38), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n582_), .B1(new_n526_), .B2(new_n531_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n325_), .A2(new_n545_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(G1gat), .B1(new_n603_), .B2(new_n454_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n598_), .A2(new_n599_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n600_), .A2(new_n604_), .A3(new_n605_), .ZN(G1324gat));
  NAND2_X1  g405(.A1(new_n495_), .A2(new_n499_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n595_), .A2(new_n286_), .A3(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n601_), .A2(new_n607_), .A3(new_n602_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(KEYINPUT99), .A2(KEYINPUT39), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n286_), .B1(KEYINPUT99), .B2(KEYINPUT39), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n609_), .A2(new_n610_), .A3(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n610_), .B1(new_n609_), .B2(new_n611_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n608_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n615_), .B(new_n617_), .ZN(G1325gat));
  OAI21_X1  g417(.A(G15gat), .B1(new_n603_), .B2(new_n525_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT41), .ZN(new_n620_));
  NOR3_X1   g419(.A1(new_n591_), .A2(G15gat), .A3(new_n525_), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n620_), .A2(new_n621_), .ZN(G1326gat));
  OAI21_X1  g421(.A(G22gat), .B1(new_n603_), .B2(new_n488_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(KEYINPUT101), .B(KEYINPUT42), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n488_), .A2(G22gat), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n625_), .B1(new_n591_), .B2(new_n626_), .ZN(G1327gat));
  XOR2_X1   g426(.A(new_n543_), .B(new_n544_), .Z(new_n628_));
  INV_X1    g427(.A(new_n582_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n532_), .A2(new_n630_), .ZN(new_n631_));
  OR3_X1    g430(.A1(new_n631_), .A2(G29gat), .A3(new_n454_), .ZN(new_n632_));
  AND4_X1   g431(.A1(KEYINPUT73), .A2(new_n572_), .A3(new_n573_), .A4(new_n576_), .ZN(new_n633_));
  AOI21_X1  g432(.A(KEYINPUT73), .B1(new_n582_), .B2(new_n573_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n589_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n525_), .ZN(new_n637_));
  AOI22_X1  g436(.A1(new_n462_), .A2(new_n488_), .B1(new_n502_), .B2(KEYINPUT95), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n637_), .B1(new_n638_), .B2(new_n501_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n531_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n636_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(KEYINPUT43), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n526_), .A2(new_n531_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT43), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n643_), .A2(new_n644_), .A3(new_n636_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n642_), .A2(new_n645_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n325_), .A2(new_n628_), .ZN(new_n647_));
  AOI21_X1  g446(.A(KEYINPUT44), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT44), .ZN(new_n649_));
  INV_X1    g448(.A(new_n647_), .ZN(new_n650_));
  AOI211_X1 g449(.A(new_n649_), .B(new_n650_), .C1(new_n642_), .C2(new_n645_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n648_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n652_), .A2(KEYINPUT102), .A3(new_n597_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(G29gat), .ZN(new_n654_));
  AOI21_X1  g453(.A(KEYINPUT102), .B1(new_n652_), .B2(new_n597_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n632_), .B1(new_n654_), .B2(new_n655_), .ZN(G1328gat));
  INV_X1    g455(.A(KEYINPUT46), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n296_), .B1(new_n652_), .B2(new_n607_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n607_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n659_), .A2(G36gat), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  OR3_X1    g460(.A1(new_n631_), .A2(KEYINPUT45), .A3(new_n661_), .ZN(new_n662_));
  OAI21_X1  g461(.A(KEYINPUT45), .B1(new_n631_), .B2(new_n661_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n657_), .B1(new_n658_), .B2(new_n665_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n648_), .A2(new_n651_), .A3(new_n659_), .ZN(new_n667_));
  OAI211_X1 g466(.A(KEYINPUT46), .B(new_n664_), .C1(new_n667_), .C2(new_n296_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(G1329gat));
  NAND2_X1  g468(.A1(new_n637_), .A2(G43gat), .ZN(new_n670_));
  NOR3_X1   g469(.A1(new_n648_), .A2(new_n651_), .A3(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n631_), .ZN(new_n672_));
  AOI21_X1  g471(.A(G43gat), .B1(new_n672_), .B2(new_n637_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(KEYINPUT103), .B(KEYINPUT47), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  OR3_X1    g474(.A1(new_n671_), .A2(new_n673_), .A3(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n675_), .B1(new_n671_), .B2(new_n673_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(G1330gat));
  NOR3_X1   g477(.A1(new_n648_), .A2(new_n651_), .A3(new_n488_), .ZN(new_n679_));
  INV_X1    g478(.A(G50gat), .ZN(new_n680_));
  INV_X1    g479(.A(new_n488_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(new_n680_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT104), .ZN(new_n683_));
  OAI22_X1  g482(.A1(new_n679_), .A2(new_n680_), .B1(new_n631_), .B2(new_n683_), .ZN(G1331gat));
  NOR2_X1   g483(.A1(new_n280_), .A2(new_n324_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n686_), .A2(new_n545_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n601_), .A2(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(G57gat), .B1(new_n688_), .B2(new_n454_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n643_), .A2(new_n590_), .A3(new_n685_), .ZN(new_n690_));
  OR2_X1    g489(.A1(new_n596_), .A2(G57gat), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n689_), .B1(new_n690_), .B2(new_n691_), .ZN(G1332gat));
  OR3_X1    g491(.A1(new_n690_), .A2(G64gat), .A3(new_n659_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n601_), .A2(new_n687_), .A3(new_n607_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT48), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n694_), .A2(new_n695_), .A3(G64gat), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n695_), .B1(new_n694_), .B2(G64gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n693_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT105), .ZN(G1333gat));
  OAI21_X1  g499(.A(G71gat), .B1(new_n688_), .B2(new_n525_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT49), .ZN(new_n702_));
  OR2_X1    g501(.A1(new_n525_), .A2(G71gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n702_), .B1(new_n690_), .B2(new_n703_), .ZN(G1334gat));
  OAI21_X1  g503(.A(G78gat), .B1(new_n688_), .B2(new_n488_), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n705_), .A2(KEYINPUT107), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(KEYINPUT107), .ZN(new_n707_));
  XOR2_X1   g506(.A(KEYINPUT106), .B(KEYINPUT50), .Z(new_n708_));
  AND3_X1   g507(.A1(new_n706_), .A2(new_n707_), .A3(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n708_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n681_), .A2(new_n477_), .ZN(new_n711_));
  OAI22_X1  g510(.A1(new_n709_), .A2(new_n710_), .B1(new_n690_), .B2(new_n711_), .ZN(G1335gat));
  NAND3_X1  g511(.A1(new_n643_), .A2(new_n630_), .A3(new_n685_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(G85gat), .B1(new_n714_), .B2(new_n597_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n686_), .A2(new_n628_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n646_), .A2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(G85gat), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n454_), .A2(new_n718_), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT108), .Z(new_n720_));
  AOI21_X1  g519(.A(new_n715_), .B1(new_n717_), .B2(new_n720_), .ZN(G1336gat));
  INV_X1    g520(.A(G92gat), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n714_), .A2(new_n722_), .A3(new_n607_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n717_), .A2(new_n607_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n723_), .B1(new_n724_), .B2(new_n722_), .ZN(G1337gat));
  INV_X1    g524(.A(KEYINPUT109), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n637_), .A2(new_n238_), .ZN(new_n727_));
  OR3_X1    g526(.A1(new_n713_), .A2(new_n726_), .A3(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n726_), .B1(new_n713_), .B2(new_n727_), .ZN(new_n729_));
  AOI22_X1  g528(.A1(new_n728_), .A2(new_n729_), .B1(KEYINPUT110), .B2(KEYINPUT51), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n646_), .A2(new_n637_), .A3(new_n716_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(G99gat), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n730_), .A2(new_n732_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n733_), .B(new_n734_), .Z(G1338gat));
  XNOR2_X1  g534(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n681_), .A2(new_n239_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n713_), .A2(new_n738_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT111), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n646_), .A2(new_n681_), .A3(new_n716_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n741_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(KEYINPUT52), .B1(new_n741_), .B2(G106gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n737_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n744_), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n746_), .A2(new_n742_), .A3(new_n740_), .A4(new_n736_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n745_), .A2(new_n747_), .ZN(G1339gat));
  AND3_X1   g547(.A1(new_n529_), .A2(new_n597_), .A3(new_n530_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n321_), .A2(new_n323_), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n750_), .A2(new_n274_), .A3(new_n276_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n635_), .A2(new_n628_), .A3(new_n751_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n752_), .A2(KEYINPUT113), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT114), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n752_), .A2(KEYINPUT113), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT54), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n755_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  AOI211_X1 g557(.A(KEYINPUT114), .B(KEYINPUT54), .C1(new_n752_), .C2(KEYINPUT113), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n754_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT113), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n761_), .B1(new_n590_), .B2(new_n751_), .ZN(new_n762_));
  OAI21_X1  g561(.A(KEYINPUT114), .B1(new_n762_), .B2(KEYINPUT54), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n756_), .A2(new_n755_), .A3(new_n757_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n763_), .A2(new_n753_), .A3(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n760_), .A2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT58), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT56), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n254_), .B(new_n249_), .C1(new_n261_), .C2(new_n262_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n263_), .A2(KEYINPUT55), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n257_), .A2(new_n258_), .A3(new_n256_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT67), .B1(new_n219_), .B2(new_n225_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n553_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n262_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT55), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n775_), .A2(new_n776_), .A3(new_n254_), .A4(new_n255_), .ZN(new_n777_));
  AOI221_X4 g576(.A(KEYINPUT115), .B1(new_n202_), .B2(new_n769_), .C1(new_n770_), .C2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT115), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n770_), .A2(new_n777_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n769_), .A2(new_n202_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n779_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n268_), .B1(new_n778_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n780_), .A2(new_n781_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT115), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n780_), .A2(new_n779_), .A3(new_n781_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n270_), .A2(new_n768_), .ZN(new_n788_));
  AOI22_X1  g587(.A1(new_n768_), .A2(new_n783_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n315_), .A2(new_n319_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(new_n316_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n310_), .A2(G229gat), .A3(new_n315_), .A4(G233gat), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(new_n284_), .A3(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n323_), .A2(new_n793_), .A3(new_n271_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n767_), .B1(new_n789_), .B2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n794_), .ZN(new_n796_));
  AOI21_X1  g595(.A(KEYINPUT56), .B1(new_n787_), .B2(new_n268_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n788_), .B1(new_n778_), .B2(new_n782_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  OAI211_X1 g598(.A(KEYINPUT58), .B(new_n796_), .C1(new_n797_), .C2(new_n799_), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n795_), .A2(new_n636_), .A3(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n323_), .A2(new_n793_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n802_), .A2(new_n273_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n783_), .A2(new_n768_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n798_), .A2(KEYINPUT116), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT116), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n806_), .B(new_n788_), .C1(new_n778_), .C2(new_n782_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n804_), .A2(new_n805_), .A3(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n324_), .A2(new_n271_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n803_), .B1(new_n808_), .B2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n629_), .A2(KEYINPUT57), .ZN(new_n812_));
  OAI21_X1  g611(.A(KEYINPUT119), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT119), .ZN(new_n814_));
  INV_X1    g613(.A(new_n812_), .ZN(new_n815_));
  AOI22_X1  g614(.A1(KEYINPUT116), .A2(new_n798_), .B1(new_n783_), .B2(new_n768_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n809_), .B1(new_n816_), .B2(new_n807_), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n814_), .B(new_n815_), .C1(new_n817_), .C2(new_n803_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n801_), .B1(new_n813_), .B2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(KEYINPUT117), .B1(new_n811_), .B2(new_n582_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT117), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n821_), .B(new_n629_), .C1(new_n817_), .C2(new_n803_), .ZN(new_n822_));
  XOR2_X1   g621(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n823_));
  NAND3_X1  g622(.A1(new_n820_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n628_), .B1(new_n819_), .B2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n749_), .B1(new_n766_), .B2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(KEYINPUT120), .ZN(new_n827_));
  INV_X1    g626(.A(G113gat), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT120), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n829_), .B(new_n749_), .C1(new_n766_), .C2(new_n825_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n827_), .A2(new_n828_), .A3(new_n324_), .A4(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT59), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n826_), .A2(new_n832_), .ZN(new_n833_));
  OAI211_X1 g632(.A(KEYINPUT59), .B(new_n749_), .C1(new_n766_), .C2(new_n825_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n750_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n831_), .B1(new_n835_), .B2(new_n828_), .ZN(G1340gat));
  INV_X1    g635(.A(new_n280_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT60), .ZN(new_n838_));
  AOI21_X1  g637(.A(G120gat), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n839_), .B1(new_n838_), .B2(G120gat), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n827_), .A2(new_n830_), .A3(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n280_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n842_));
  INV_X1    g641(.A(G120gat), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n841_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(KEYINPUT121), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT121), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n846_), .B(new_n841_), .C1(new_n842_), .C2(new_n843_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(G1341gat));
  INV_X1    g647(.A(G127gat), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n827_), .A2(new_n849_), .A3(new_n628_), .A4(new_n830_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n545_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n850_), .B1(new_n851_), .B2(new_n849_), .ZN(G1342gat));
  INV_X1    g651(.A(G134gat), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n827_), .A2(new_n853_), .A3(new_n582_), .A4(new_n830_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n635_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n855_), .B2(new_n853_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(KEYINPUT122), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT122), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n858_), .B(new_n854_), .C1(new_n855_), .C2(new_n853_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n859_), .ZN(G1343gat));
  OR2_X1    g659(.A1(new_n766_), .A2(new_n825_), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n659_), .A2(new_n597_), .A3(new_n681_), .A4(new_n525_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(KEYINPUT123), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n324_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g666(.A1(new_n865_), .A2(new_n837_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g668(.A1(new_n865_), .A2(new_n628_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(KEYINPUT61), .B(G155gat), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n870_), .B(new_n871_), .ZN(G1346gat));
  NAND3_X1  g671(.A1(new_n865_), .A2(G162gat), .A3(new_n636_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(G162gat), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n875_), .B1(new_n864_), .B2(new_n629_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT124), .ZN(new_n877_));
  OR2_X1    g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n877_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n874_), .B1(new_n878_), .B2(new_n879_), .ZN(G1347gat));
  NOR3_X1   g679(.A1(new_n659_), .A2(new_n597_), .A3(new_n525_), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n881_), .A2(new_n324_), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n488_), .B(new_n882_), .C1(new_n766_), .C2(new_n825_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(G169gat), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n884_), .B(KEYINPUT62), .C1(new_n424_), .C2(new_n883_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT62), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n883_), .A2(new_n886_), .A3(G169gat), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n885_), .A2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(KEYINPUT125), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT125), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n885_), .A2(new_n890_), .A3(new_n887_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n891_), .ZN(G1348gat));
  XNOR2_X1  g691(.A(KEYINPUT126), .B(G176gat), .ZN(new_n893_));
  AND2_X1   g692(.A1(new_n861_), .A2(new_n488_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n881_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n893_), .B1(new_n895_), .B2(new_n280_), .ZN(new_n896_));
  OR2_X1    g695(.A1(KEYINPUT126), .A2(G176gat), .ZN(new_n897_));
  NAND4_X1  g696(.A1(new_n894_), .A2(new_n837_), .A3(new_n881_), .A4(new_n897_), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n896_), .A2(new_n898_), .ZN(G1349gat));
  OAI22_X1  g698(.A1(new_n895_), .A2(new_n545_), .B1(KEYINPUT127), .B2(G183gat), .ZN(new_n900_));
  INV_X1    g699(.A(new_n392_), .ZN(new_n901_));
  INV_X1    g700(.A(G183gat), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n901_), .B1(KEYINPUT127), .B2(new_n902_), .ZN(new_n903_));
  NAND4_X1  g702(.A1(new_n894_), .A2(new_n628_), .A3(new_n881_), .A4(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n900_), .A2(new_n904_), .ZN(G1350gat));
  OAI21_X1  g704(.A(G190gat), .B1(new_n895_), .B2(new_n635_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n582_), .A2(new_n393_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n895_), .B2(new_n907_), .ZN(G1351gat));
  AND3_X1   g707(.A1(new_n607_), .A2(new_n525_), .A3(new_n500_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n861_), .A2(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n324_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g712(.A1(new_n911_), .A2(new_n837_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g714(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n916_));
  AND2_X1   g715(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n917_));
  NOR4_X1   g716(.A1(new_n910_), .A2(new_n545_), .A3(new_n916_), .A4(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n911_), .A2(new_n628_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n918_), .B1(new_n919_), .B2(new_n916_), .ZN(G1354gat));
  INV_X1    g719(.A(G218gat), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n911_), .A2(new_n921_), .A3(new_n582_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n911_), .A2(new_n636_), .ZN(new_n923_));
  INV_X1    g722(.A(new_n923_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n922_), .B1(new_n924_), .B2(new_n921_), .ZN(G1355gat));
endmodule


