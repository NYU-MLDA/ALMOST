//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 0 0 1 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 1 1 1 0 1 1 0 0 0 1 1 1 0 1 1 1 0 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n672_,
    new_n673_, new_n674_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n747_, new_n748_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n783_, new_n784_,
    new_n785_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n883_, new_n885_,
    new_n886_, new_n888_, new_n889_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n902_, new_n903_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n910_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n938_, new_n939_, new_n940_, new_n942_, new_n943_,
    new_n945_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n953_, new_n954_;
  INV_X1    g000(.A(G120gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G127gat), .A2(G134gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  NOR2_X1   g003(.A1(G127gat), .A2(G134gat), .ZN(new_n205_));
  NOR3_X1   g004(.A1(new_n204_), .A2(new_n205_), .A3(G113gat), .ZN(new_n206_));
  INV_X1    g005(.A(G113gat), .ZN(new_n207_));
  INV_X1    g006(.A(G127gat), .ZN(new_n208_));
  INV_X1    g007(.A(G134gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n207_), .B1(new_n210_), .B2(new_n203_), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n202_), .B1(new_n206_), .B2(new_n211_), .ZN(new_n212_));
  OAI21_X1  g011(.A(G113gat), .B1(new_n204_), .B2(new_n205_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n210_), .A2(new_n207_), .A3(new_n203_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n213_), .A2(new_n214_), .A3(G120gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n212_), .A2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT31), .ZN(new_n217_));
  XOR2_X1   g016(.A(G15gat), .B(G43gat), .Z(new_n218_));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT78), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT78), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(G183gat), .A3(G190gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n220_), .A2(new_n222_), .A3(KEYINPUT23), .ZN(new_n223_));
  INV_X1    g022(.A(G183gat), .ZN(new_n224_));
  AND2_X1   g023(.A1(KEYINPUT77), .A2(G190gat), .ZN(new_n225_));
  NOR2_X1   g024(.A1(KEYINPUT77), .A2(G190gat), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n224_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT23), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n219_), .A2(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n223_), .A2(new_n227_), .A3(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT81), .ZN(new_n231_));
  AND2_X1   g030(.A1(KEYINPUT79), .A2(KEYINPUT22), .ZN(new_n232_));
  NOR2_X1   g031(.A1(KEYINPUT79), .A2(KEYINPUT22), .ZN(new_n233_));
  OAI21_X1  g032(.A(G169gat), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT80), .ZN(new_n235_));
  INV_X1    g034(.A(G176gat), .ZN(new_n236_));
  INV_X1    g035(.A(G169gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT22), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT80), .ZN(new_n239_));
  OAI211_X1 g038(.A(new_n239_), .B(G169gat), .C1(new_n232_), .C2(new_n233_), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n235_), .A2(new_n236_), .A3(new_n238_), .A4(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G169gat), .A2(G176gat), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT81), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n223_), .A2(new_n227_), .A3(new_n243_), .A4(new_n229_), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n231_), .A2(new_n241_), .A3(new_n242_), .A4(new_n244_), .ZN(new_n245_));
  XOR2_X1   g044(.A(KEYINPUT25), .B(G183gat), .Z(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT76), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT76), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT25), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n248_), .B1(new_n249_), .B2(G183gat), .ZN(new_n250_));
  OAI21_X1  g049(.A(KEYINPUT26), .B1(new_n225_), .B2(new_n226_), .ZN(new_n251_));
  INV_X1    g050(.A(G190gat), .ZN(new_n252_));
  OR2_X1    g051(.A1(new_n252_), .A2(KEYINPUT26), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n247_), .A2(new_n250_), .A3(new_n251_), .A4(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n237_), .A2(new_n236_), .ZN(new_n255_));
  OR2_X1    g054(.A1(new_n255_), .A2(KEYINPUT24), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n255_), .A2(KEYINPUT24), .A3(new_n242_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n220_), .A2(new_n222_), .A3(new_n228_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n219_), .A2(KEYINPUT23), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n254_), .A2(new_n256_), .A3(new_n257_), .A4(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G227gat), .A2(G233gat), .ZN(new_n262_));
  XOR2_X1   g061(.A(new_n262_), .B(KEYINPUT30), .Z(new_n263_));
  NAND3_X1  g062(.A1(new_n245_), .A2(new_n261_), .A3(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n263_), .B1(new_n245_), .B2(new_n261_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n218_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n245_), .A2(new_n261_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n263_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n218_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n270_), .A2(new_n271_), .A3(new_n264_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G71gat), .B(G99gat), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n267_), .A2(new_n272_), .A3(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n273_), .B1(new_n267_), .B2(new_n272_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n217_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT83), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT83), .ZN(new_n279_));
  OAI211_X1 g078(.A(new_n279_), .B(new_n217_), .C1(new_n275_), .C2(new_n276_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n276_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n217_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n282_), .A2(new_n283_), .A3(new_n274_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT82), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n282_), .A2(KEYINPUT82), .A3(new_n283_), .A4(new_n274_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  AND2_X1   g087(.A1(new_n281_), .A2(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NOR3_X1   g090(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  AND3_X1   g092(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n294_));
  AOI21_X1  g093(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(KEYINPUT84), .B1(G155gat), .B2(G162gat), .ZN(new_n297_));
  NOR2_X1   g096(.A1(G155gat), .A2(G162gat), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT84), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  AOI22_X1  g099(.A1(new_n293_), .A2(new_n296_), .B1(new_n297_), .B2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G155gat), .A2(G162gat), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT85), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(KEYINPUT85), .A2(G155gat), .A3(G162gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  AND3_X1   g105(.A1(KEYINPUT85), .A2(G155gat), .A3(G162gat), .ZN(new_n307_));
  AOI21_X1  g106(.A(KEYINPUT85), .B1(G155gat), .B2(G162gat), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT1), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n300_), .A2(new_n297_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT1), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n304_), .A2(new_n311_), .A3(new_n305_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n309_), .A2(new_n310_), .A3(new_n312_), .ZN(new_n313_));
  XOR2_X1   g112(.A(G141gat), .B(G148gat), .Z(new_n314_));
  AOI22_X1  g113(.A1(new_n301_), .A2(new_n306_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT29), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G22gat), .B(G50gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT28), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n317_), .B(new_n319_), .ZN(new_n320_));
  XOR2_X1   g119(.A(G78gat), .B(G106gat), .Z(new_n321_));
  XOR2_X1   g120(.A(G211gat), .B(G218gat), .Z(new_n322_));
  INV_X1    g121(.A(G197gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(G204gat), .ZN(new_n324_));
  INV_X1    g123(.A(G204gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(G197gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n324_), .A2(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT87), .B1(new_n327_), .B2(KEYINPUT21), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G197gat), .B(G204gat), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT87), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT21), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n329_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n322_), .B1(new_n328_), .B2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n323_), .A2(KEYINPUT86), .A3(G204gat), .ZN(new_n334_));
  OAI211_X1 g133(.A(KEYINPUT21), .B(new_n334_), .C1(new_n327_), .C2(KEYINPUT86), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n329_), .A2(new_n331_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(new_n322_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G228gat), .A2(G233gat), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n339_), .B(new_n340_), .C1(new_n316_), .C2(new_n315_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n293_), .A2(new_n296_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n342_), .A2(new_n310_), .A3(new_n306_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n313_), .A2(new_n314_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n316_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  AOI22_X1  g144(.A1(new_n333_), .A2(new_n335_), .B1(new_n322_), .B2(new_n337_), .ZN(new_n346_));
  OAI211_X1 g145(.A(G228gat), .B(G233gat), .C1(new_n345_), .C2(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n321_), .B1(new_n341_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT88), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n320_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n341_), .A2(new_n347_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n321_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n341_), .A2(new_n347_), .A3(new_n321_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n350_), .A2(new_n355_), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n353_), .A2(new_n320_), .A3(new_n349_), .A4(new_n354_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT33), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G225gat), .A2(G233gat), .ZN(new_n360_));
  XOR2_X1   g159(.A(new_n360_), .B(KEYINPUT92), .Z(new_n361_));
  NAND2_X1  g160(.A1(new_n343_), .A2(new_n344_), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n362_), .A2(KEYINPUT93), .A3(KEYINPUT4), .A4(new_n216_), .ZN(new_n363_));
  AND2_X1   g162(.A1(new_n212_), .A2(new_n215_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT93), .ZN(new_n365_));
  NOR3_X1   g164(.A1(new_n315_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT4), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n367_), .B1(new_n315_), .B2(new_n364_), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n361_), .B(new_n363_), .C1(new_n366_), .C2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n361_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n362_), .A2(new_n216_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n315_), .A2(new_n364_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n370_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n369_), .A2(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT0), .B(G57gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(G85gat), .ZN(new_n376_));
  XOR2_X1   g175(.A(G1gat), .B(G29gat), .Z(new_n377_));
  XOR2_X1   g176(.A(new_n376_), .B(new_n377_), .Z(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n374_), .A2(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n359_), .B1(new_n380_), .B2(KEYINPUT94), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n378_), .B1(new_n369_), .B2(new_n373_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT94), .ZN(new_n383_));
  NOR3_X1   g182(.A1(new_n382_), .A2(new_n383_), .A3(KEYINPUT33), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n381_), .A2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n346_), .A2(new_n245_), .A3(new_n261_), .ZN(new_n386_));
  XOR2_X1   g185(.A(KEYINPUT26), .B(G190gat), .Z(new_n387_));
  NOR2_X1   g186(.A1(new_n246_), .A2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT89), .B(KEYINPUT24), .ZN(new_n389_));
  AND3_X1   g188(.A1(new_n389_), .A2(new_n255_), .A3(new_n242_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n223_), .A2(new_n229_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n389_), .A2(new_n255_), .ZN(new_n392_));
  NOR4_X1   g191(.A1(new_n388_), .A2(new_n390_), .A3(new_n391_), .A4(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT91), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT22), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(G169gat), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n238_), .A2(new_n396_), .A3(new_n236_), .ZN(new_n397_));
  AND3_X1   g196(.A1(new_n397_), .A2(KEYINPUT90), .A3(new_n242_), .ZN(new_n398_));
  AOI21_X1  g197(.A(KEYINPUT90), .B1(new_n397_), .B2(new_n242_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n224_), .A2(new_n252_), .ZN(new_n401_));
  AND2_X1   g200(.A1(new_n260_), .A2(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n394_), .B1(new_n400_), .B2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n260_), .A2(new_n401_), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n404_), .B(KEYINPUT91), .C1(new_n399_), .C2(new_n398_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n393_), .B1(new_n403_), .B2(new_n405_), .ZN(new_n406_));
  OAI211_X1 g205(.A(KEYINPUT20), .B(new_n386_), .C1(new_n406_), .C2(new_n346_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G226gat), .A2(G233gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT19), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(KEYINPUT18), .B(G64gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(G92gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G8gat), .B(G36gat), .ZN(new_n413_));
  XOR2_X1   g212(.A(new_n412_), .B(new_n413_), .Z(new_n414_));
  NAND2_X1  g213(.A1(new_n406_), .A2(new_n346_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n409_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n268_), .A2(new_n339_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n415_), .A2(KEYINPUT20), .A3(new_n416_), .A4(new_n417_), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n410_), .A2(new_n414_), .A3(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n414_), .B1(new_n410_), .B2(new_n418_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  OR3_X1    g220(.A1(new_n371_), .A2(new_n372_), .A3(new_n370_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n366_), .A2(new_n368_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n423_), .B1(KEYINPUT4), .B2(new_n366_), .ZN(new_n424_));
  OAI211_X1 g223(.A(new_n378_), .B(new_n422_), .C1(new_n424_), .C2(new_n361_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n385_), .A2(new_n421_), .A3(new_n425_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n374_), .A2(new_n379_), .ZN(new_n427_));
  OR2_X1    g226(.A1(new_n427_), .A2(new_n382_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n414_), .A2(KEYINPUT32), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n410_), .A2(new_n418_), .A3(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n400_), .A2(new_n402_), .ZN(new_n431_));
  NOR3_X1   g230(.A1(new_n339_), .A2(new_n431_), .A3(new_n393_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n346_), .B1(new_n245_), .B2(new_n261_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n416_), .B1(new_n434_), .B2(KEYINPUT20), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n407_), .A2(new_n409_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  OAI211_X1 g236(.A(new_n428_), .B(new_n430_), .C1(new_n437_), .C2(new_n429_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n358_), .B1(new_n426_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n428_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT27), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n441_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n414_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n443_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n410_), .A2(new_n414_), .A3(new_n418_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n444_), .A2(KEYINPUT27), .A3(new_n445_), .ZN(new_n446_));
  AND4_X1   g245(.A1(new_n440_), .A2(new_n442_), .A3(new_n446_), .A4(new_n358_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n289_), .B1(new_n439_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n358_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n449_), .A2(new_n442_), .A3(new_n446_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT95), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n281_), .A2(new_n288_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT95), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n449_), .A2(new_n442_), .A3(new_n446_), .A4(new_n453_), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n451_), .A2(new_n452_), .A3(new_n440_), .A4(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n448_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT75), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT15), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G29gat), .B(G36gat), .ZN(new_n459_));
  OR2_X1    g258(.A1(new_n459_), .A2(G43gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(G43gat), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n460_), .A2(G50gat), .A3(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(G50gat), .B1(new_n460_), .B2(new_n461_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n458_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n460_), .A2(new_n461_), .ZN(new_n466_));
  INV_X1    g265(.A(G50gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n468_), .A2(KEYINPUT15), .A3(new_n462_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n465_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(G8gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(KEYINPUT73), .B(G1gat), .ZN(new_n472_));
  OAI21_X1  g271(.A(KEYINPUT14), .B1(new_n472_), .B2(new_n471_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G15gat), .B(G22gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(G1gat), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n475_), .A2(G1gat), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n471_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  OR2_X1    g278(.A1(new_n475_), .A2(G1gat), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n480_), .A2(G8gat), .A3(new_n476_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n470_), .A2(new_n479_), .A3(new_n481_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n463_), .A2(new_n464_), .ZN(new_n483_));
  NOR3_X1   g282(.A1(new_n477_), .A2(new_n478_), .A3(new_n471_), .ZN(new_n484_));
  AOI21_X1  g283(.A(G8gat), .B1(new_n480_), .B2(new_n476_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n483_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G229gat), .A2(G233gat), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n482_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n483_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n479_), .A2(new_n490_), .A3(new_n481_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n487_), .B1(new_n486_), .B2(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n457_), .B1(new_n489_), .B2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G113gat), .B(G141gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(new_n237_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(new_n323_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n493_), .A2(new_n497_), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n457_), .B(new_n496_), .C1(new_n489_), .C2(new_n492_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n456_), .A2(new_n500_), .ZN(new_n501_));
  AND2_X1   g300(.A1(new_n501_), .A2(KEYINPUT96), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n501_), .A2(KEYINPUT96), .ZN(new_n503_));
  OR2_X1    g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  AND2_X1   g303(.A1(G85gat), .A2(G92gat), .ZN(new_n505_));
  NOR2_X1   g304(.A1(G85gat), .A2(G92gat), .ZN(new_n506_));
  OAI21_X1  g305(.A(KEYINPUT9), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT65), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n507_), .B(new_n508_), .C1(KEYINPUT9), .C2(new_n505_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT66), .ZN(new_n510_));
  NAND3_X1  g309(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n510_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G99gat), .A2(G106gat), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT6), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n517_), .A2(KEYINPUT66), .A3(new_n511_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n514_), .A2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n505_), .A2(KEYINPUT65), .A3(KEYINPUT9), .ZN(new_n520_));
  XOR2_X1   g319(.A(KEYINPUT10), .B(G99gat), .Z(new_n521_));
  INV_X1    g320(.A(G106gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n509_), .A2(new_n519_), .A3(new_n520_), .A4(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT67), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT7), .ZN(new_n526_));
  INV_X1    g325(.A(G99gat), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n526_), .A2(new_n527_), .A3(new_n522_), .ZN(new_n528_));
  OAI21_X1  g327(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n519_), .A2(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n505_), .A2(new_n506_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT8), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n532_), .A2(new_n536_), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n528_), .A2(new_n517_), .A3(new_n511_), .A4(new_n529_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(new_n533_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT8), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n525_), .B1(new_n537_), .B2(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n530_), .B1(new_n514_), .B2(new_n518_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n542_), .A2(new_n535_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n534_), .B1(new_n538_), .B2(new_n533_), .ZN(new_n544_));
  NOR3_X1   g343(.A1(new_n543_), .A2(KEYINPUT67), .A3(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n524_), .B1(new_n541_), .B2(new_n545_), .ZN(new_n546_));
  XOR2_X1   g345(.A(G57gat), .B(G64gat), .Z(new_n547_));
  INV_X1    g346(.A(KEYINPUT11), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G57gat), .B(G64gat), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(KEYINPUT11), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G71gat), .B(G78gat), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n549_), .A2(new_n551_), .A3(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n550_), .A2(new_n552_), .A3(KEYINPUT11), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT12), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n546_), .A2(new_n558_), .ZN(new_n559_));
  OAI211_X1 g358(.A(new_n556_), .B(new_n524_), .C1(new_n543_), .C2(new_n544_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n540_), .B1(new_n542_), .B2(new_n535_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(new_n524_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n556_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n561_), .B1(new_n565_), .B2(new_n557_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G230gat), .A2(G233gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT64), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n559_), .A2(new_n566_), .A3(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n568_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n556_), .B1(new_n562_), .B2(new_n524_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n570_), .B1(new_n561_), .B2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n569_), .A2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G120gat), .B(G148gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(new_n325_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT5), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(new_n236_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n573_), .A2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n569_), .A2(new_n572_), .A3(new_n577_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n581_), .B1(KEYINPUT68), .B2(KEYINPUT13), .ZN(new_n582_));
  NOR2_X1   g381(.A1(KEYINPUT68), .A2(KEYINPUT13), .ZN(new_n583_));
  AND2_X1   g382(.A1(KEYINPUT68), .A2(KEYINPUT13), .ZN(new_n584_));
  OAI211_X1 g383(.A(new_n579_), .B(new_n580_), .C1(new_n583_), .C2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n582_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n479_), .A2(new_n481_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(G231gat), .A2(G233gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n556_), .B(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n587_), .B(new_n589_), .Z(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(KEYINPUT16), .B(G183gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(G211gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G127gat), .B(G155gat), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n593_), .B(new_n594_), .Z(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NOR3_X1   g395(.A1(new_n591_), .A2(KEYINPUT17), .A3(new_n596_), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n590_), .A2(KEYINPUT74), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n596_), .A2(KEYINPUT17), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n599_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n597_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT37), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT71), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n483_), .A2(new_n562_), .A3(new_n524_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n465_), .A2(new_n469_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n524_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n537_), .A2(new_n525_), .A3(new_n540_), .ZN(new_n608_));
  OAI21_X1  g407(.A(KEYINPUT67), .B1(new_n543_), .B2(new_n544_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n607_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n605_), .B1(new_n606_), .B2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(G232gat), .A2(G233gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT34), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n613_), .A2(KEYINPUT35), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(KEYINPUT35), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n604_), .B1(new_n611_), .B2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n546_), .A2(new_n470_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n614_), .A2(new_n615_), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n618_), .A2(KEYINPUT71), .A3(new_n605_), .A4(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n617_), .A2(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(KEYINPUT70), .B(G134gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(G162gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G190gat), .B(G218gat), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n623_), .B(new_n624_), .Z(new_n625_));
  NOR2_X1   g424(.A1(new_n625_), .A2(KEYINPUT36), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n611_), .A2(KEYINPUT69), .A3(new_n614_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(KEYINPUT69), .B1(new_n611_), .B2(new_n614_), .ZN(new_n629_));
  OAI211_X1 g428(.A(new_n621_), .B(new_n626_), .C1(new_n628_), .C2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT72), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n603_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n629_), .ZN(new_n633_));
  AOI22_X1  g432(.A1(new_n633_), .A2(new_n627_), .B1(new_n617_), .B2(new_n620_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n625_), .B(KEYINPUT36), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n630_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n632_), .A2(new_n636_), .ZN(new_n637_));
  OAI221_X1 g436(.A(new_n630_), .B1(new_n631_), .B2(new_n603_), .C1(new_n634_), .C2(new_n635_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n602_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n504_), .A2(new_n586_), .A3(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n641_), .A2(new_n428_), .A3(new_n472_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT38), .ZN(new_n643_));
  AND3_X1   g442(.A1(new_n586_), .A2(KEYINPUT97), .A3(new_n500_), .ZN(new_n644_));
  AOI21_X1  g443(.A(KEYINPUT97), .B1(new_n586_), .B2(new_n500_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n636_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n602_), .A2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n646_), .A2(new_n456_), .A3(new_n648_), .ZN(new_n649_));
  OAI21_X1  g448(.A(G1gat), .B1(new_n649_), .B2(new_n440_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n643_), .A2(new_n650_), .ZN(G1324gat));
  NAND2_X1  g450(.A1(new_n442_), .A2(new_n446_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(new_n471_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT39), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n646_), .A2(new_n456_), .A3(new_n652_), .A4(new_n648_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n654_), .B1(new_n655_), .B2(G8gat), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n655_), .A2(new_n654_), .A3(G8gat), .ZN(new_n657_));
  OAI22_X1  g456(.A1(new_n640_), .A2(new_n653_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(KEYINPUT98), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT98), .ZN(new_n660_));
  OAI221_X1 g459(.A(new_n660_), .B1(new_n657_), .B2(new_n656_), .C1(new_n640_), .C2(new_n653_), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n659_), .A2(new_n661_), .A3(KEYINPUT40), .ZN(new_n662_));
  AOI21_X1  g461(.A(KEYINPUT40), .B1(new_n659_), .B2(new_n661_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1325gat));
  OR3_X1    g463(.A1(new_n640_), .A2(G15gat), .A3(new_n289_), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n665_), .A2(KEYINPUT100), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(KEYINPUT100), .ZN(new_n667_));
  OAI21_X1  g466(.A(G15gat), .B1(new_n649_), .B2(new_n289_), .ZN(new_n668_));
  XOR2_X1   g467(.A(KEYINPUT99), .B(KEYINPUT41), .Z(new_n669_));
  XNOR2_X1  g468(.A(new_n668_), .B(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n666_), .A2(new_n667_), .A3(new_n670_), .ZN(G1326gat));
  OAI21_X1  g470(.A(G22gat), .B1(new_n649_), .B2(new_n449_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT42), .ZN(new_n673_));
  OR2_X1    g472(.A1(new_n449_), .A2(G22gat), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n673_), .B1(new_n640_), .B2(new_n674_), .ZN(G1327gat));
  INV_X1    g474(.A(new_n602_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n586_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n504_), .A2(new_n647_), .A3(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(G29gat), .B1(new_n680_), .B2(new_n428_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n646_), .A2(new_n602_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT43), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT101), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n448_), .A2(new_n686_), .A3(new_n455_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n686_), .B1(new_n448_), .B2(new_n455_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n637_), .A2(new_n638_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n685_), .B1(new_n689_), .B2(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n456_), .A2(new_n685_), .A3(new_n691_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT102), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(KEYINPUT43), .B1(new_n448_), .B2(new_n455_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n696_), .A2(KEYINPUT102), .A3(new_n691_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(new_n698_));
  OAI211_X1 g497(.A(new_n682_), .B(new_n684_), .C1(new_n692_), .C2(new_n698_), .ZN(new_n699_));
  XOR2_X1   g498(.A(KEYINPUT104), .B(KEYINPUT44), .Z(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n701_), .A2(KEYINPUT103), .ZN(new_n702_));
  AND4_X1   g501(.A1(KEYINPUT102), .A2(new_n456_), .A3(new_n685_), .A4(new_n691_), .ZN(new_n703_));
  AOI21_X1  g502(.A(KEYINPUT102), .B1(new_n696_), .B2(new_n691_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n456_), .A2(KEYINPUT101), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n448_), .A2(new_n455_), .A3(new_n686_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n706_), .A2(new_n691_), .A3(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(KEYINPUT43), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n683_), .B1(new_n705_), .B2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT103), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n701_), .A2(new_n711_), .ZN(new_n712_));
  OAI22_X1  g511(.A1(new_n699_), .A2(new_n702_), .B1(new_n710_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n714_), .A2(new_n440_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n681_), .B1(new_n715_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g515(.A(new_n652_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n717_), .A2(G36gat), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(KEYINPUT45), .B1(new_n679_), .B2(new_n719_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n502_), .A2(new_n503_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n721_), .A2(new_n636_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT45), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n722_), .A2(new_n723_), .A3(new_n678_), .A4(new_n718_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n720_), .A2(new_n724_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n692_), .A2(new_n698_), .ZN(new_n726_));
  OAI22_X1  g525(.A1(new_n726_), .A2(new_n683_), .B1(new_n711_), .B2(new_n701_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n702_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n710_), .A2(new_n682_), .A3(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n717_), .B1(new_n727_), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(G36gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n725_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT105), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n733_), .A2(KEYINPUT46), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(new_n735_));
  OAI221_X1 g534(.A(new_n725_), .B1(new_n733_), .B2(KEYINPUT46), .C1(new_n730_), .C2(new_n731_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(G1329gat));
  INV_X1    g536(.A(G43gat), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n738_), .B1(new_n713_), .B2(new_n452_), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n679_), .A2(G43gat), .A3(new_n289_), .ZN(new_n740_));
  OAI21_X1  g539(.A(KEYINPUT47), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n740_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT47), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n289_), .B1(new_n727_), .B2(new_n729_), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n742_), .B(new_n743_), .C1(new_n744_), .C2(new_n738_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n741_), .A2(new_n745_), .ZN(G1330gat));
  AOI21_X1  g545(.A(G50gat), .B1(new_n680_), .B2(new_n358_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n714_), .A2(new_n449_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n748_), .B2(G50gat), .ZN(G1331gat));
  AOI211_X1 g548(.A(new_n500_), .B(new_n586_), .C1(new_n448_), .C2(new_n455_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(new_n639_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT106), .ZN(new_n752_));
  AOI21_X1  g551(.A(G57gat), .B1(new_n752_), .B2(new_n428_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n750_), .A2(new_n648_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n754_), .A2(new_n428_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n753_), .B1(G57gat), .B2(new_n755_), .ZN(G1332gat));
  INV_X1    g555(.A(G64gat), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n757_), .B1(new_n754_), .B2(new_n652_), .ZN(new_n758_));
  XOR2_X1   g557(.A(new_n758_), .B(KEYINPUT48), .Z(new_n759_));
  NAND3_X1  g558(.A1(new_n752_), .A2(new_n757_), .A3(new_n652_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(G1333gat));
  INV_X1    g560(.A(G71gat), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n762_), .B1(new_n754_), .B2(new_n452_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT107), .ZN(new_n764_));
  XOR2_X1   g563(.A(new_n764_), .B(KEYINPUT49), .Z(new_n765_));
  NAND3_X1  g564(.A1(new_n752_), .A2(new_n762_), .A3(new_n452_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(G1334gat));
  INV_X1    g566(.A(G78gat), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n768_), .B1(new_n754_), .B2(new_n358_), .ZN(new_n769_));
  XOR2_X1   g568(.A(new_n769_), .B(KEYINPUT50), .Z(new_n770_));
  NAND3_X1  g569(.A1(new_n752_), .A2(new_n768_), .A3(new_n358_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(G1335gat));
  NOR3_X1   g571(.A1(new_n676_), .A2(new_n500_), .A3(new_n586_), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n456_), .A2(new_n647_), .A3(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(G85gat), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n774_), .A2(new_n775_), .A3(new_n428_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n705_), .A2(new_n709_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n777_), .A2(new_n773_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(new_n428_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n776_), .B1(new_n779_), .B2(G85gat), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT108), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n780_), .B(new_n781_), .ZN(G1336gat));
  AOI21_X1  g581(.A(G92gat), .B1(new_n774_), .B2(new_n652_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n652_), .A2(G92gat), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT109), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n783_), .B1(new_n778_), .B2(new_n785_), .ZN(G1337gat));
  AND2_X1   g585(.A1(new_n452_), .A2(new_n521_), .ZN(new_n787_));
  AOI21_X1  g586(.A(KEYINPUT110), .B1(new_n774_), .B2(new_n787_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n778_), .A2(new_n452_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n788_), .B1(new_n789_), .B2(new_n527_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT51), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n792_), .B(new_n788_), .C1(new_n789_), .C2(new_n527_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n791_), .A2(new_n793_), .ZN(G1338gat));
  NAND3_X1  g593(.A1(new_n777_), .A2(new_n358_), .A3(new_n773_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(G106gat), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT111), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n796_), .A2(new_n797_), .A3(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n774_), .A2(new_n522_), .A3(new_n358_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n797_), .A2(new_n798_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(KEYINPUT111), .A2(KEYINPUT52), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n795_), .A2(G106gat), .A3(new_n801_), .A4(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n799_), .A2(new_n800_), .A3(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(KEYINPUT53), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n799_), .A2(new_n806_), .A3(new_n800_), .A4(new_n803_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n805_), .A2(new_n807_), .ZN(G1339gat));
  INV_X1    g607(.A(new_n558_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n608_), .A2(new_n609_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n809_), .B1(new_n810_), .B2(new_n524_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n560_), .B1(new_n571_), .B2(KEYINPUT12), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n570_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n569_), .A2(new_n813_), .A3(KEYINPUT55), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT55), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n559_), .A2(new_n566_), .A3(new_n815_), .A4(new_n568_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n814_), .A2(new_n578_), .A3(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(KEYINPUT56), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT56), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n814_), .A2(new_n819_), .A3(new_n578_), .A4(new_n816_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n818_), .A2(new_n820_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n821_), .A2(KEYINPUT114), .A3(new_n500_), .A4(new_n580_), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n489_), .A2(new_n492_), .A3(new_n496_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n482_), .A2(new_n486_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n487_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n486_), .A2(new_n487_), .A3(new_n491_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n497_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n823_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT115), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n829_), .A2(new_n581_), .A3(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n830_), .B1(new_n829_), .B2(new_n581_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n500_), .A2(new_n818_), .A3(new_n580_), .A4(new_n820_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT114), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n822_), .A2(new_n834_), .A3(new_n837_), .ZN(new_n838_));
  AND3_X1   g637(.A1(new_n838_), .A2(KEYINPUT57), .A3(new_n636_), .ZN(new_n839_));
  AOI21_X1  g638(.A(KEYINPUT57), .B1(new_n838_), .B2(new_n636_), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n818_), .A2(new_n580_), .A3(new_n820_), .A4(new_n829_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT58), .ZN(new_n842_));
  AND3_X1   g641(.A1(new_n841_), .A2(KEYINPUT116), .A3(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n842_), .B1(new_n841_), .B2(KEYINPUT116), .ZN(new_n844_));
  NOR3_X1   g643(.A1(new_n843_), .A2(new_n690_), .A3(new_n844_), .ZN(new_n845_));
  NOR3_X1   g644(.A1(new_n839_), .A2(new_n840_), .A3(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(KEYINPUT119), .B1(new_n846_), .B2(new_n676_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n848_));
  INV_X1    g647(.A(new_n500_), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n639_), .A2(new_n848_), .A3(new_n849_), .A4(new_n586_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n850_), .A2(KEYINPUT112), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n850_), .A2(KEYINPUT112), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n690_), .A2(new_n849_), .A3(new_n676_), .A4(new_n586_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT113), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n853_), .A2(new_n854_), .A3(KEYINPUT54), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n854_), .B1(new_n853_), .B2(KEYINPUT54), .ZN(new_n856_));
  OAI22_X1  g655(.A1(new_n851_), .A2(new_n852_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n838_), .A2(new_n636_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT57), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n845_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n838_), .A2(KEYINPUT57), .A3(new_n636_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n860_), .A2(new_n861_), .A3(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT119), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n863_), .A2(new_n864_), .A3(new_n602_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n847_), .A2(new_n857_), .A3(new_n865_), .ZN(new_n866_));
  XOR2_X1   g665(.A(KEYINPUT117), .B(KEYINPUT59), .Z(new_n867_));
  AND4_X1   g666(.A1(new_n428_), .A2(new_n451_), .A3(new_n452_), .A4(new_n454_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(KEYINPUT118), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n866_), .A2(new_n867_), .A3(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n863_), .A2(new_n602_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n857_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n868_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(KEYINPUT59), .ZN(new_n874_));
  OAI21_X1  g673(.A(G113gat), .B1(new_n849_), .B2(KEYINPUT120), .ZN(new_n875_));
  OR2_X1    g674(.A1(KEYINPUT120), .A2(G113gat), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n870_), .A2(new_n874_), .A3(new_n875_), .A4(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n207_), .B1(new_n873_), .B2(new_n849_), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n877_), .A2(new_n878_), .ZN(G1340gat));
  INV_X1    g678(.A(new_n873_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n202_), .B1(new_n586_), .B2(KEYINPUT60), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n880_), .B(new_n881_), .C1(KEYINPUT60), .C2(new_n202_), .ZN(new_n882_));
  AND3_X1   g681(.A1(new_n870_), .A2(new_n677_), .A3(new_n874_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n883_), .B2(new_n202_), .ZN(G1341gat));
  NAND4_X1  g683(.A1(new_n870_), .A2(new_n874_), .A3(G127gat), .A4(new_n676_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n208_), .B1(new_n873_), .B2(new_n602_), .ZN(new_n886_));
  AND2_X1   g685(.A1(new_n885_), .A2(new_n886_), .ZN(G1342gat));
  NAND4_X1  g686(.A1(new_n870_), .A2(new_n874_), .A3(G134gat), .A4(new_n691_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n209_), .B1(new_n873_), .B2(new_n636_), .ZN(new_n889_));
  AND2_X1   g688(.A1(new_n888_), .A2(new_n889_), .ZN(G1343gat));
  NOR2_X1   g689(.A1(new_n452_), .A2(new_n449_), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n872_), .A2(new_n428_), .A3(new_n717_), .A4(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT121), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n891_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n895_), .B1(new_n871_), .B2(new_n857_), .ZN(new_n896_));
  NAND4_X1  g695(.A1(new_n896_), .A2(KEYINPUT121), .A3(new_n428_), .A4(new_n717_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n849_), .B1(new_n894_), .B2(new_n897_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(KEYINPUT122), .B(G141gat), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n898_), .B(new_n899_), .ZN(G1344gat));
  AOI21_X1  g699(.A(new_n586_), .B1(new_n894_), .B2(new_n897_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(KEYINPUT123), .B(G148gat), .ZN(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n901_), .B(new_n903_), .ZN(G1345gat));
  AOI21_X1  g703(.A(new_n602_), .B1(new_n894_), .B2(new_n897_), .ZN(new_n905_));
  XOR2_X1   g704(.A(KEYINPUT61), .B(G155gat), .Z(new_n906_));
  XNOR2_X1  g705(.A(KEYINPUT124), .B(KEYINPUT125), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n906_), .B(new_n907_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n905_), .B(new_n908_), .ZN(G1346gat));
  NAND2_X1  g708(.A1(new_n894_), .A2(new_n897_), .ZN(new_n910_));
  AND3_X1   g709(.A1(new_n910_), .A2(G162gat), .A3(new_n691_), .ZN(new_n911_));
  AOI21_X1  g710(.A(G162gat), .B1(new_n910_), .B2(new_n647_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n911_), .A2(new_n912_), .ZN(G1347gat));
  NOR2_X1   g712(.A1(new_n717_), .A2(new_n428_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n914_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n915_), .A2(new_n289_), .ZN(new_n916_));
  NAND4_X1  g715(.A1(new_n866_), .A2(new_n500_), .A3(new_n449_), .A4(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(G169gat), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT62), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n917_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n238_), .A2(new_n396_), .ZN(new_n922_));
  OAI211_X1 g721(.A(new_n920_), .B(new_n921_), .C1(new_n922_), .C2(new_n917_), .ZN(G1348gat));
  NAND4_X1  g722(.A1(new_n866_), .A2(new_n677_), .A3(new_n449_), .A4(new_n916_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(new_n236_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n358_), .B1(new_n871_), .B2(new_n857_), .ZN(new_n926_));
  NAND4_X1  g725(.A1(new_n926_), .A2(G176gat), .A3(new_n677_), .A4(new_n916_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n925_), .A2(new_n927_), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT126), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n925_), .A2(KEYINPUT126), .A3(new_n927_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(G1349gat));
  NOR3_X1   g731(.A1(new_n915_), .A2(new_n289_), .A3(new_n602_), .ZN(new_n933_));
  AOI21_X1  g732(.A(G183gat), .B1(new_n926_), .B2(new_n933_), .ZN(new_n934_));
  AND2_X1   g733(.A1(new_n866_), .A2(new_n449_), .ZN(new_n935_));
  AND2_X1   g734(.A1(new_n933_), .A2(new_n246_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n934_), .B1(new_n935_), .B2(new_n936_), .ZN(G1350gat));
  NOR2_X1   g736(.A1(new_n636_), .A2(new_n387_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n935_), .A2(new_n916_), .A3(new_n938_), .ZN(new_n939_));
  AND3_X1   g738(.A1(new_n935_), .A2(new_n691_), .A3(new_n916_), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n939_), .B1(new_n940_), .B2(new_n252_), .ZN(G1351gat));
  NAND2_X1  g740(.A1(new_n896_), .A2(new_n914_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n942_), .A2(new_n849_), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n943_), .B(new_n323_), .ZN(G1352gat));
  NOR2_X1   g743(.A1(new_n942_), .A2(new_n586_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(new_n945_), .B(new_n325_), .ZN(G1353gat));
  NOR2_X1   g745(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n947_));
  AND2_X1   g746(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n948_));
  NOR4_X1   g747(.A1(new_n942_), .A2(new_n602_), .A3(new_n947_), .A4(new_n948_), .ZN(new_n949_));
  INV_X1    g748(.A(new_n942_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n950_), .A2(new_n676_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n949_), .B1(new_n951_), .B2(new_n947_), .ZN(G1354gat));
  AND3_X1   g751(.A1(new_n950_), .A2(G218gat), .A3(new_n691_), .ZN(new_n953_));
  AOI21_X1  g752(.A(G218gat), .B1(new_n950_), .B2(new_n647_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n953_), .A2(new_n954_), .ZN(G1355gat));
endmodule


