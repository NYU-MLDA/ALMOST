//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 1 0 0 1 0 0 0 0 0 0 1 0 1 0 0 1 0 1 1 1 0 0 0 1 1 0 1 0 0 0 0 0 1 0 0 1 0 0 0 1 1 1 1 1 1 1 0 1 0 1 0 1 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n594_, new_n595_, new_n596_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n641_, new_n642_, new_n643_, new_n645_, new_n646_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n694_,
    new_n695_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n804_, new_n805_, new_n806_, new_n808_, new_n810_, new_n811_,
    new_n813_, new_n814_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n839_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n848_, new_n849_, new_n850_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n871_, new_n872_;
  NOR2_X1   g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT86), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT1), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n204_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G141gat), .ZN(new_n209_));
  INV_X1    g008(.A(G148gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G141gat), .A2(G148gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n208_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n212_), .B(KEYINPUT2), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT87), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n211_), .B1(new_n215_), .B2(KEYINPUT3), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT3), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n217_), .A2(new_n209_), .A3(new_n210_), .A4(KEYINPUT87), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n214_), .A2(new_n216_), .A3(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n219_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n220_));
  AND2_X1   g019(.A1(new_n213_), .A2(new_n220_), .ZN(new_n221_));
  XOR2_X1   g020(.A(G127gat), .B(G134gat), .Z(new_n222_));
  XOR2_X1   g021(.A(G113gat), .B(G120gat), .Z(new_n223_));
  XOR2_X1   g022(.A(new_n222_), .B(new_n223_), .Z(new_n224_));
  XNOR2_X1  g023(.A(new_n221_), .B(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT4), .ZN(new_n226_));
  INV_X1    g025(.A(new_n224_), .ZN(new_n227_));
  OR3_X1    g026(.A1(new_n221_), .A2(KEYINPUT4), .A3(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G225gat), .A2(G233gat), .ZN(new_n229_));
  XOR2_X1   g028(.A(new_n229_), .B(KEYINPUT95), .Z(new_n230_));
  NAND3_X1  g029(.A1(new_n226_), .A2(new_n228_), .A3(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n225_), .A2(new_n229_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G1gat), .B(G29gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(G85gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT0), .B(G57gat), .ZN(new_n235_));
  XOR2_X1   g034(.A(new_n234_), .B(new_n235_), .Z(new_n236_));
  NAND3_X1  g035(.A1(new_n231_), .A2(new_n232_), .A3(new_n236_), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n237_), .A2(KEYINPUT98), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(KEYINPUT98), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n231_), .A2(new_n232_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n236_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n238_), .A2(new_n239_), .A3(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT99), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n238_), .A2(KEYINPUT99), .A3(new_n239_), .A4(new_n242_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G227gat), .A2(G233gat), .ZN(new_n248_));
  INV_X1    g047(.A(G15gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT30), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT31), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G71gat), .B(G99gat), .ZN(new_n254_));
  INV_X1    g053(.A(G43gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G183gat), .A2(G190gat), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n258_), .A2(KEYINPUT23), .ZN(new_n259_));
  XOR2_X1   g058(.A(KEYINPUT83), .B(KEYINPUT23), .Z(new_n260_));
  AOI21_X1  g059(.A(new_n259_), .B1(new_n260_), .B2(new_n258_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT24), .ZN(new_n262_));
  NOR2_X1   g061(.A1(G169gat), .A2(G176gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT81), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n261_), .B1(new_n262_), .B2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT84), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G169gat), .A2(G176gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(KEYINPUT24), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n264_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT82), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT25), .B(G183gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(KEYINPUT26), .B(G190gat), .ZN(new_n272_));
  AOI22_X1  g071(.A1(new_n269_), .A2(new_n270_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n266_), .B(new_n273_), .C1(new_n270_), .C2(new_n269_), .ZN(new_n274_));
  AOI21_X1  g073(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n275_));
  AND2_X1   g074(.A1(G183gat), .A2(G190gat), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n275_), .B1(new_n260_), .B2(new_n276_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n277_), .B1(G183gat), .B2(G190gat), .ZN(new_n278_));
  INV_X1    g077(.A(G176gat), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT22), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT85), .B1(new_n280_), .B2(G169gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT22), .B(G169gat), .ZN(new_n282_));
  OAI211_X1 g081(.A(new_n279_), .B(new_n281_), .C1(new_n282_), .C2(KEYINPUT85), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n278_), .A2(new_n267_), .A3(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n257_), .B1(new_n274_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n274_), .A2(new_n284_), .A3(new_n257_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n227_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n287_), .ZN(new_n289_));
  NOR3_X1   g088(.A1(new_n289_), .A2(new_n224_), .A3(new_n285_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n253_), .B1(new_n288_), .B2(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n224_), .B1(new_n289_), .B2(new_n285_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n286_), .A2(new_n227_), .A3(new_n287_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n292_), .A2(new_n293_), .A3(new_n252_), .ZN(new_n294_));
  AND2_X1   g093(.A1(new_n291_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G78gat), .B(G106gat), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  XOR2_X1   g096(.A(G22gat), .B(G50gat), .Z(new_n298_));
  INV_X1    g097(.A(KEYINPUT29), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n221_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT28), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT88), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT28), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n221_), .A2(new_n303_), .A3(new_n299_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n301_), .A2(new_n302_), .A3(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n302_), .B1(new_n301_), .B2(new_n304_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n298_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n307_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n298_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n309_), .A2(new_n310_), .A3(new_n305_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n297_), .B1(new_n308_), .B2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n296_), .A2(KEYINPUT93), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n308_), .A2(new_n311_), .A3(new_n314_), .ZN(new_n315_));
  XOR2_X1   g114(.A(G211gat), .B(G218gat), .Z(new_n316_));
  INV_X1    g115(.A(G204gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(G197gat), .ZN(new_n318_));
  INV_X1    g117(.A(G197gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(G204gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n316_), .B1(KEYINPUT21), .B2(new_n321_), .ZN(new_n322_));
  OR2_X1    g121(.A1(new_n318_), .A2(KEYINPUT89), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n318_), .A2(KEYINPUT89), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n323_), .A2(new_n324_), .A3(new_n320_), .ZN(new_n325_));
  XOR2_X1   g124(.A(KEYINPUT90), .B(KEYINPUT21), .Z(new_n326_));
  OAI21_X1  g125(.A(new_n322_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  XOR2_X1   g126(.A(new_n327_), .B(KEYINPUT91), .Z(new_n328_));
  NAND3_X1  g127(.A1(new_n325_), .A2(KEYINPUT21), .A3(new_n316_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n330_), .B1(new_n299_), .B2(new_n221_), .ZN(new_n331_));
  AND3_X1   g130(.A1(KEYINPUT92), .A2(G228gat), .A3(G233gat), .ZN(new_n332_));
  OR2_X1    g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(KEYINPUT92), .B1(G228gat), .B2(G233gat), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n331_), .B1(new_n334_), .B2(new_n332_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  AND3_X1   g135(.A1(new_n313_), .A2(new_n315_), .A3(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n336_), .B1(new_n313_), .B2(new_n315_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n295_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n315_), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n335_), .B(new_n333_), .C1(new_n340_), .C2(new_n312_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n291_), .A2(new_n294_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n313_), .A2(new_n315_), .A3(new_n336_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n341_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n247_), .B1(new_n339_), .B2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT20), .ZN(new_n346_));
  NOR2_X1   g145(.A1(G183gat), .A2(G190gat), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n261_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n282_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n267_), .B1(new_n349_), .B2(G176gat), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n269_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n264_), .A2(new_n262_), .ZN(new_n353_));
  AND3_X1   g152(.A1(new_n352_), .A2(new_n277_), .A3(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n271_), .B(KEYINPUT94), .ZN(new_n355_));
  INV_X1    g154(.A(new_n272_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n351_), .B1(new_n354_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n346_), .B1(new_n330_), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n274_), .A2(new_n284_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n361_), .B1(new_n362_), .B2(new_n330_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G226gat), .A2(G233gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT19), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT20), .B1(new_n330_), .B2(new_n360_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n362_), .A2(new_n330_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n365_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n368_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G8gat), .B(G36gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT18), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G64gat), .B(G92gat), .ZN(new_n374_));
  XOR2_X1   g173(.A(new_n373_), .B(new_n374_), .Z(new_n375_));
  NAND3_X1  g174(.A1(new_n366_), .A2(new_n371_), .A3(new_n375_), .ZN(new_n376_));
  OR2_X1    g175(.A1(new_n376_), .A2(KEYINPUT100), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(KEYINPUT100), .ZN(new_n378_));
  INV_X1    g177(.A(new_n330_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n379_), .B1(new_n284_), .B2(new_n274_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n365_), .B1(new_n380_), .B2(new_n367_), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n361_), .B(new_n370_), .C1(new_n362_), .C2(new_n330_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n375_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n377_), .A2(KEYINPUT27), .A3(new_n378_), .A4(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n366_), .A2(new_n371_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(new_n384_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(new_n376_), .ZN(new_n389_));
  XOR2_X1   g188(.A(KEYINPUT101), .B(KEYINPUT27), .Z(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  AND2_X1   g190(.A1(new_n386_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n237_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n226_), .A2(new_n229_), .A3(new_n228_), .ZN(new_n394_));
  XOR2_X1   g193(.A(new_n394_), .B(KEYINPUT96), .Z(new_n395_));
  AOI21_X1  g194(.A(new_n236_), .B1(new_n225_), .B2(new_n230_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n393_), .B1(new_n397_), .B2(KEYINPUT33), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n393_), .A2(KEYINPUT33), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n388_), .A2(new_n376_), .A3(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n375_), .A2(KEYINPUT32), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n381_), .A2(new_n382_), .A3(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n366_), .A2(new_n371_), .A3(KEYINPUT97), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT97), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n366_), .A2(new_n371_), .A3(new_n405_), .ZN(new_n406_));
  AOI22_X1  g205(.A1(new_n403_), .A2(new_n404_), .B1(new_n406_), .B2(new_n401_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n243_), .ZN(new_n408_));
  OAI22_X1  g207(.A1(new_n398_), .A2(new_n400_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n295_), .B1(new_n341_), .B2(new_n343_), .ZN(new_n410_));
  AOI22_X1  g209(.A1(new_n345_), .A2(new_n392_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G230gat), .A2(G233gat), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G99gat), .A2(G106gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT6), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT6), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n416_), .A2(G99gat), .A3(G106gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n415_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT66), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT7), .ZN(new_n421_));
  INV_X1    g220(.A(G99gat), .ZN(new_n422_));
  INV_X1    g221(.A(G106gat), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n421_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n415_), .A2(new_n417_), .A3(KEYINPUT66), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n420_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  XOR2_X1   g228(.A(G85gat), .B(G92gat), .Z(new_n430_));
  INV_X1    g229(.A(KEYINPUT8), .ZN(new_n431_));
  AND2_X1   g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n429_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT67), .ZN(new_n434_));
  AND2_X1   g233(.A1(new_n415_), .A2(new_n417_), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n434_), .B(new_n430_), .C1(new_n435_), .C2(new_n426_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT8), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n418_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n434_), .B1(new_n438_), .B2(new_n430_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n433_), .B1(new_n437_), .B2(new_n439_), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n420_), .A2(new_n428_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(KEYINPUT65), .B(G85gat), .ZN(new_n442_));
  INV_X1    g241(.A(G92gat), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n443_), .A2(KEYINPUT9), .ZN(new_n444_));
  AOI22_X1  g243(.A1(new_n430_), .A2(KEYINPUT9), .B1(new_n442_), .B2(new_n444_), .ZN(new_n445_));
  XOR2_X1   g244(.A(KEYINPUT10), .B(G99gat), .Z(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(KEYINPUT64), .ZN(new_n447_));
  OAI211_X1 g246(.A(new_n441_), .B(new_n445_), .C1(new_n447_), .C2(G106gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n440_), .A2(new_n448_), .ZN(new_n449_));
  OR2_X1    g248(.A1(KEYINPUT68), .A2(G71gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(KEYINPUT68), .A2(G71gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(G78gat), .ZN(new_n453_));
  INV_X1    g252(.A(G78gat), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n450_), .A2(new_n454_), .A3(new_n451_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G57gat), .B(G64gat), .ZN(new_n456_));
  AOI22_X1  g255(.A1(new_n453_), .A2(new_n455_), .B1(KEYINPUT11), .B2(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(KEYINPUT11), .ZN(new_n458_));
  AND2_X1   g257(.A1(new_n453_), .A2(new_n455_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n457_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n449_), .A2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n440_), .A2(new_n460_), .A3(new_n448_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n462_), .A2(KEYINPUT12), .A3(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n460_), .B1(new_n440_), .B2(new_n448_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT12), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n413_), .B1(new_n464_), .B2(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n412_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G120gat), .B(G148gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n470_), .B(KEYINPUT5), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G176gat), .B(G204gat), .ZN(new_n472_));
  XOR2_X1   g271(.A(new_n471_), .B(new_n472_), .Z(new_n473_));
  OR3_X1    g272(.A1(new_n468_), .A2(new_n469_), .A3(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n473_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n475_));
  AND2_X1   g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  OR2_X1    g275(.A1(new_n476_), .A2(KEYINPUT13), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(KEYINPUT13), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(KEYINPUT74), .B(G15gat), .ZN(new_n481_));
  INV_X1    g280(.A(G22gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n481_), .B(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT75), .B(G1gat), .ZN(new_n484_));
  INV_X1    g283(.A(G8gat), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT14), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n483_), .A2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G1gat), .B(G8gat), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n483_), .A2(new_n486_), .A3(new_n488_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  XOR2_X1   g291(.A(G29gat), .B(G36gat), .Z(new_n493_));
  XOR2_X1   g292(.A(G43gat), .B(G50gat), .Z(new_n494_));
  XOR2_X1   g293(.A(new_n493_), .B(new_n494_), .Z(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n492_), .B(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n497_), .A2(G229gat), .A3(G233gat), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT15), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n495_), .B(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n500_), .A2(new_n491_), .A3(new_n490_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n492_), .A2(new_n496_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G229gat), .A2(G233gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT79), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n501_), .A2(new_n502_), .A3(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n498_), .A2(new_n505_), .ZN(new_n506_));
  XOR2_X1   g305(.A(G113gat), .B(G141gat), .Z(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT80), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G169gat), .B(G197gat), .ZN(new_n509_));
  XOR2_X1   g308(.A(new_n508_), .B(new_n509_), .Z(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n506_), .A2(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n498_), .A2(new_n505_), .A3(new_n510_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n480_), .A2(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n411_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT71), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n500_), .A2(new_n449_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G232gat), .A2(G233gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  OR2_X1    g320(.A1(new_n521_), .A2(KEYINPUT35), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n440_), .A2(new_n448_), .A3(new_n496_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n518_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n524_), .A2(KEYINPUT35), .A3(new_n521_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n521_), .A2(KEYINPUT35), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n518_), .A2(new_n526_), .A3(new_n522_), .A4(new_n523_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n525_), .A2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G190gat), .B(G218gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT70), .ZN(new_n530_));
  XOR2_X1   g329(.A(G134gat), .B(G162gat), .Z(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n532_), .A2(KEYINPUT36), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n517_), .B1(new_n528_), .B2(new_n534_), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n525_), .A2(KEYINPUT71), .A3(new_n533_), .A4(new_n527_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n532_), .B(KEYINPUT36), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n528_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n537_), .A2(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n541_), .A2(KEYINPUT37), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT72), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n537_), .A2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n538_), .B(KEYINPUT73), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n528_), .A2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n535_), .A2(KEYINPUT72), .A3(new_n536_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n544_), .A2(new_n546_), .A3(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n542_), .B1(KEYINPUT37), .B2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G231gat), .A2(G233gat), .ZN(new_n550_));
  XOR2_X1   g349(.A(new_n550_), .B(KEYINPUT76), .Z(new_n551_));
  XNOR2_X1  g350(.A(new_n492_), .B(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(new_n461_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT17), .ZN(new_n554_));
  XOR2_X1   g353(.A(G127gat), .B(G155gat), .Z(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT78), .ZN(new_n556_));
  XOR2_X1   g355(.A(G183gat), .B(G211gat), .Z(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  XOR2_X1   g357(.A(KEYINPUT77), .B(KEYINPUT16), .Z(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  OR3_X1    g359(.A1(new_n553_), .A2(new_n554_), .A3(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(KEYINPUT17), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(new_n553_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n549_), .A2(new_n564_), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n516_), .A2(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n566_), .A2(new_n484_), .A3(new_n247_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT38), .ZN(new_n568_));
  OR2_X1    g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n568_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n541_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n411_), .A2(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n515_), .A2(new_n564_), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n245_), .A2(new_n246_), .ZN(new_n576_));
  OAI21_X1  g375(.A(G1gat), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n569_), .A2(new_n570_), .A3(new_n577_), .ZN(G1324gat));
  XNOR2_X1  g377(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n485_), .B1(KEYINPUT103), .B2(KEYINPUT39), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n581_), .B1(new_n575_), .B2(new_n392_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(KEYINPUT103), .A2(KEYINPUT39), .ZN(new_n583_));
  OR2_X1    g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n582_), .A2(new_n583_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n386_), .A2(new_n391_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n566_), .A2(new_n485_), .A3(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT102), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n580_), .B1(new_n586_), .B2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n589_), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n591_), .A2(new_n584_), .A3(new_n585_), .A4(new_n579_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n590_), .A2(new_n592_), .ZN(G1325gat));
  AOI21_X1  g392(.A(new_n249_), .B1(new_n574_), .B2(new_n295_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT41), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n566_), .A2(new_n249_), .A3(new_n295_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(G1326gat));
  NOR2_X1   g396(.A1(new_n337_), .A2(new_n338_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n482_), .B1(new_n574_), .B2(new_n598_), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n599_), .B(KEYINPUT42), .Z(new_n600_));
  NAND3_X1  g399(.A1(new_n566_), .A2(new_n482_), .A3(new_n598_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(G1327gat));
  INV_X1    g401(.A(new_n564_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n603_), .A2(new_n541_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n516_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(G29gat), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n605_), .A2(new_n606_), .A3(new_n247_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n549_), .ZN(new_n608_));
  OAI21_X1  g407(.A(KEYINPUT43), .B1(new_n411_), .B2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n409_), .A2(new_n410_), .ZN(new_n610_));
  AND3_X1   g409(.A1(new_n341_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n342_), .B1(new_n341_), .B2(new_n343_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n576_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n610_), .B1(new_n613_), .B2(new_n587_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT43), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n614_), .A2(new_n615_), .A3(new_n549_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n609_), .A2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n480_), .A2(new_n564_), .A3(new_n514_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(KEYINPUT44), .B1(new_n617_), .B2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT44), .ZN(new_n621_));
  AOI211_X1 g420(.A(new_n621_), .B(new_n618_), .C1(new_n609_), .C2(new_n616_), .ZN(new_n622_));
  NOR3_X1   g421(.A1(new_n620_), .A2(new_n622_), .A3(new_n576_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n607_), .B1(new_n623_), .B2(new_n606_), .ZN(G1328gat));
  INV_X1    g423(.A(G36gat), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n605_), .A2(new_n625_), .A3(new_n587_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT45), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n617_), .A2(new_n619_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(new_n621_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT105), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n617_), .A2(KEYINPUT44), .A3(new_n619_), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n629_), .A2(new_n630_), .A3(new_n587_), .A4(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(G36gat), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n620_), .A2(new_n622_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n630_), .B1(new_n634_), .B2(new_n587_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n627_), .B1(new_n633_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT46), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  OAI211_X1 g437(.A(KEYINPUT46), .B(new_n627_), .C1(new_n633_), .C2(new_n635_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(G1329gat));
  NAND3_X1  g439(.A1(new_n605_), .A2(new_n255_), .A3(new_n295_), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n620_), .A2(new_n622_), .A3(new_n342_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n641_), .B1(new_n642_), .B2(new_n255_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g443(.A(G50gat), .B1(new_n605_), .B2(new_n598_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n598_), .A2(G50gat), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n645_), .B1(new_n634_), .B2(new_n646_), .ZN(G1331gat));
  NOR2_X1   g446(.A1(new_n564_), .A2(new_n514_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n479_), .A2(new_n648_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n572_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(G57gat), .B1(new_n651_), .B2(new_n576_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n411_), .A2(new_n514_), .ZN(new_n653_));
  AND3_X1   g452(.A1(new_n653_), .A2(new_n565_), .A3(new_n479_), .ZN(new_n654_));
  INV_X1    g453(.A(G57gat), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n654_), .A2(new_n655_), .A3(new_n247_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n652_), .A2(new_n656_), .ZN(G1332gat));
  INV_X1    g456(.A(G64gat), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n654_), .A2(new_n658_), .A3(new_n587_), .ZN(new_n659_));
  OAI21_X1  g458(.A(G64gat), .B1(new_n651_), .B2(new_n392_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n660_), .A2(KEYINPUT48), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n660_), .A2(KEYINPUT48), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n659_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT106), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  OAI211_X1 g464(.A(KEYINPUT106), .B(new_n659_), .C1(new_n661_), .C2(new_n662_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(G1333gat));
  INV_X1    g466(.A(G71gat), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n668_), .B1(new_n650_), .B2(new_n295_), .ZN(new_n669_));
  XOR2_X1   g468(.A(new_n669_), .B(KEYINPUT49), .Z(new_n670_));
  NAND2_X1  g469(.A1(new_n295_), .A2(new_n668_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT107), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n654_), .A2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n670_), .A2(new_n673_), .ZN(G1334gat));
  NAND3_X1  g473(.A1(new_n654_), .A2(new_n454_), .A3(new_n598_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n598_), .ZN(new_n676_));
  OAI21_X1  g475(.A(G78gat), .B1(new_n651_), .B2(new_n676_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n677_), .A2(KEYINPUT50), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n677_), .A2(KEYINPUT50), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n675_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(KEYINPUT108), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT108), .ZN(new_n682_));
  OAI211_X1 g481(.A(new_n682_), .B(new_n675_), .C1(new_n678_), .C2(new_n679_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n681_), .A2(new_n683_), .ZN(G1335gat));
  AND2_X1   g483(.A1(new_n479_), .A2(new_n604_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n653_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(G85gat), .B1(new_n687_), .B2(new_n247_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT109), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n603_), .A2(new_n514_), .ZN(new_n690_));
  AND3_X1   g489(.A1(new_n617_), .A2(new_n479_), .A3(new_n690_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n247_), .A2(new_n442_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n689_), .B1(new_n691_), .B2(new_n692_), .ZN(G1336gat));
  NAND3_X1  g492(.A1(new_n687_), .A2(new_n443_), .A3(new_n587_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n691_), .A2(new_n587_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n694_), .B1(new_n695_), .B2(new_n443_), .ZN(G1337gat));
  OR3_X1    g495(.A1(new_n686_), .A2(new_n447_), .A3(new_n342_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n691_), .A2(new_n295_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n697_), .B1(new_n698_), .B2(new_n422_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g499(.A1(new_n617_), .A2(new_n598_), .A3(new_n479_), .A4(new_n690_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(G106gat), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n702_), .A2(KEYINPUT52), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT52), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n704_), .B1(new_n701_), .B2(G106gat), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n598_), .A2(new_n423_), .ZN(new_n706_));
  OAI22_X1  g505(.A1(new_n703_), .A2(new_n705_), .B1(new_n686_), .B2(new_n706_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(KEYINPUT110), .B(KEYINPUT53), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n707_), .B(new_n708_), .ZN(G1339gat));
  INV_X1    g508(.A(KEYINPUT57), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(KEYINPUT114), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n514_), .A2(new_n474_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT55), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n713_), .B1(new_n413_), .B2(KEYINPUT112), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n464_), .B2(new_n467_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n464_), .A2(new_n467_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n714_), .B1(new_n717_), .B2(new_n412_), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n440_), .A2(new_n460_), .A3(new_n448_), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n719_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n467_), .ZN(new_n721_));
  OAI21_X1  g520(.A(KEYINPUT55), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  AOI211_X1 g521(.A(KEYINPUT113), .B(new_n716_), .C1(new_n718_), .C2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT113), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n412_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n725_), .A2(new_n722_), .A3(new_n715_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n716_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n724_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n473_), .B1(new_n723_), .B2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT56), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  OAI211_X1 g530(.A(KEYINPUT56), .B(new_n473_), .C1(new_n723_), .C2(new_n728_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n712_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n497_), .A2(new_n504_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n504_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n501_), .A2(new_n502_), .A3(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n734_), .A2(new_n511_), .A3(new_n736_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n513_), .A2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n476_), .A2(new_n739_), .ZN(new_n740_));
  OAI211_X1 g539(.A(new_n541_), .B(new_n711_), .C1(new_n733_), .C2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n738_), .A2(new_n474_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n742_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n549_), .B1(new_n743_), .B2(KEYINPUT58), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT58), .ZN(new_n745_));
  AOI211_X1 g544(.A(new_n745_), .B(new_n742_), .C1(new_n731_), .C2(new_n732_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n741_), .B1(new_n744_), .B2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n712_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n713_), .B1(new_n464_), .B2(new_n467_), .ZN(new_n749_));
  NOR3_X1   g548(.A1(new_n468_), .A2(new_n749_), .A3(new_n714_), .ZN(new_n750_));
  OAI21_X1  g549(.A(KEYINPUT113), .B1(new_n750_), .B2(new_n716_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n726_), .A2(new_n724_), .A3(new_n727_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(KEYINPUT56), .B1(new_n753_), .B2(new_n473_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n732_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n748_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n740_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n711_), .B1(new_n758_), .B2(new_n541_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n564_), .B1(new_n747_), .B2(new_n759_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n477_), .A2(new_n478_), .A3(new_n648_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT111), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n761_), .A2(new_n762_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n608_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT54), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT54), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n767_), .B(new_n608_), .C1(new_n763_), .C2(new_n764_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n760_), .A2(new_n769_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n587_), .A2(new_n576_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n612_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT115), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n770_), .A2(new_n773_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT59), .ZN(new_n775_));
  INV_X1    g574(.A(new_n514_), .ZN(new_n776_));
  OAI21_X1  g575(.A(G113gat), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n774_), .A2(KEYINPUT116), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT116), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n770_), .A2(new_n779_), .A3(new_n773_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(G113gat), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n781_), .A2(new_n782_), .A3(new_n514_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n777_), .A2(new_n783_), .ZN(G1340gat));
  INV_X1    g583(.A(G120gat), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n785_), .B1(new_n480_), .B2(KEYINPUT60), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n781_), .B(new_n786_), .C1(KEYINPUT60), .C2(new_n785_), .ZN(new_n787_));
  OAI21_X1  g586(.A(G120gat), .B1(new_n775_), .B2(new_n480_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(G1341gat));
  AOI21_X1  g588(.A(G127gat), .B1(new_n781_), .B2(new_n603_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n775_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n603_), .A2(G127gat), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n792_), .B(KEYINPUT117), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n790_), .B1(new_n791_), .B2(new_n793_), .ZN(G1342gat));
  NAND3_X1  g593(.A1(new_n778_), .A2(new_n571_), .A3(new_n780_), .ZN(new_n795_));
  INV_X1    g594(.A(G134gat), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT118), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT118), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n795_), .A2(new_n799_), .A3(new_n796_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n549_), .A2(G134gat), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n801_), .B(KEYINPUT119), .ZN(new_n802_));
  AOI22_X1  g601(.A1(new_n798_), .A2(new_n800_), .B1(new_n791_), .B2(new_n802_), .ZN(G1343gat));
  AOI21_X1  g602(.A(new_n344_), .B1(new_n760_), .B2(new_n769_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n771_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n805_), .A2(new_n776_), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n806_), .B(new_n209_), .ZN(G1344gat));
  NOR2_X1   g606(.A1(new_n805_), .A2(new_n480_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(new_n210_), .ZN(G1345gat));
  NOR2_X1   g608(.A1(new_n805_), .A2(new_n564_), .ZN(new_n810_));
  XOR2_X1   g609(.A(KEYINPUT61), .B(G155gat), .Z(new_n811_));
  XNOR2_X1  g610(.A(new_n810_), .B(new_n811_), .ZN(G1346gat));
  OAI21_X1  g611(.A(G162gat), .B1(new_n805_), .B2(new_n608_), .ZN(new_n813_));
  OR2_X1    g612(.A1(new_n541_), .A2(G162gat), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n813_), .B1(new_n805_), .B2(new_n814_), .ZN(G1347gat));
  INV_X1    g614(.A(KEYINPUT121), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n392_), .A2(new_n247_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n612_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n770_), .A2(new_n514_), .A3(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT120), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n818_), .B1(new_n760_), .B2(new_n769_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n823_), .A2(KEYINPUT120), .A3(new_n514_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n822_), .A2(KEYINPUT62), .A3(G169gat), .A4(new_n824_), .ZN(new_n825_));
  AOI211_X1 g624(.A(new_n776_), .B(new_n818_), .C1(new_n760_), .C2(new_n769_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n282_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n825_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(G169gat), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n829_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n830_));
  AOI21_X1  g629(.A(KEYINPUT62), .B1(new_n830_), .B2(new_n824_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n816_), .B1(new_n828_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT62), .ZN(new_n833_));
  OAI21_X1  g632(.A(G169gat), .B1(new_n826_), .B2(KEYINPUT120), .ZN(new_n834_));
  INV_X1    g633(.A(new_n824_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n833_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n836_), .A2(KEYINPUT121), .A3(new_n827_), .A4(new_n825_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n832_), .A2(new_n837_), .ZN(G1348gat));
  NAND2_X1  g637(.A1(new_n823_), .A2(new_n479_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n839_), .B(G176gat), .ZN(G1349gat));
  INV_X1    g639(.A(new_n823_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n841_), .A2(new_n564_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n355_), .ZN(new_n843_));
  OR2_X1    g642(.A1(new_n843_), .A2(KEYINPUT122), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n842_), .A2(G183gat), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(KEYINPUT122), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n844_), .B1(new_n845_), .B2(new_n846_), .ZN(G1350gat));
  OAI21_X1  g646(.A(G190gat), .B1(new_n841_), .B2(new_n608_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n848_), .B(KEYINPUT123), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n823_), .A2(new_n571_), .A3(new_n272_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(G1351gat));
  XNOR2_X1  g650(.A(KEYINPUT124), .B(G197gat), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n319_), .A2(KEYINPUT124), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n804_), .A2(new_n817_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n854_), .A2(new_n776_), .ZN(new_n855_));
  MUX2_X1   g654(.A(new_n852_), .B(new_n853_), .S(new_n855_), .Z(G1352gat));
  INV_X1    g655(.A(new_n854_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n479_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n317_), .A2(KEYINPUT125), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n858_), .B(new_n859_), .ZN(G1353gat));
  NOR2_X1   g659(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n861_), .B1(new_n854_), .B2(new_n564_), .ZN(new_n862_));
  OR2_X1    g661(.A1(new_n862_), .A2(KEYINPUT127), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(KEYINPUT127), .ZN(new_n864_));
  XOR2_X1   g663(.A(KEYINPUT63), .B(G211gat), .Z(new_n865_));
  NAND3_X1  g664(.A1(new_n857_), .A2(new_n603_), .A3(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT126), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n857_), .A2(KEYINPUT126), .A3(new_n603_), .A4(new_n865_), .ZN(new_n869_));
  AOI22_X1  g668(.A1(new_n863_), .A2(new_n864_), .B1(new_n868_), .B2(new_n869_), .ZN(G1354gat));
  OR3_X1    g669(.A1(new_n854_), .A2(G218gat), .A3(new_n541_), .ZN(new_n871_));
  OAI21_X1  g670(.A(G218gat), .B1(new_n854_), .B2(new_n608_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(G1355gat));
endmodule


