//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 1 1 1 0 0 1 1 0 1 1 0 1 0 0 0 0 1 0 0 1 1 1 0 1 0 1 1 0 0 1 1 1 0 0 1 0 1 0 1 0 0 1 0 1 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n693_, new_n694_, new_n695_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n846_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n914_, new_n915_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n923_, new_n924_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G190gat), .B(G218gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G134gat), .B(G162gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n205_), .A2(KEYINPUT36), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT9), .ZN(new_n208_));
  INV_X1    g007(.A(G85gat), .ZN(new_n209_));
  INV_X1    g008(.A(G92gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G85gat), .A2(G92gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT64), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n208_), .B(new_n211_), .C1(new_n213_), .C2(new_n214_), .ZN(new_n215_));
  XOR2_X1   g014(.A(KEYINPUT10), .B(G99gat), .Z(new_n216_));
  INV_X1    g015(.A(G106gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n211_), .A2(KEYINPUT64), .A3(KEYINPUT9), .A4(new_n212_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G99gat), .A2(G106gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT6), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT6), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n222_), .A2(G99gat), .A3(G106gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n221_), .A2(new_n223_), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n215_), .A2(new_n218_), .A3(new_n219_), .A4(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT8), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n226_), .A2(KEYINPUT65), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NOR3_X1   g028(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  AOI211_X1 g030(.A(new_n213_), .B(new_n227_), .C1(new_n231_), .C2(new_n224_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n227_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT7), .ZN(new_n234_));
  INV_X1    g033(.A(G99gat), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n234_), .A2(new_n235_), .A3(new_n217_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n222_), .B1(G99gat), .B2(G106gat), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n220_), .A2(KEYINPUT6), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n228_), .B(new_n236_), .C1(new_n237_), .C2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n213_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n233_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n225_), .B1(new_n232_), .B2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G29gat), .B(G36gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G43gat), .B(G50gat), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n244_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n242_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G232gat), .A2(G233gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT34), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n251_), .A2(KEYINPUT35), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n249_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT68), .B(KEYINPUT15), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n247_), .B(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT69), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n255_), .A2(new_n256_), .A3(new_n242_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n256_), .B1(new_n255_), .B2(new_n242_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n253_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n251_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT35), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n259_), .A2(new_n262_), .ZN(new_n263_));
  OAI221_X1 g062(.A(new_n253_), .B1(new_n261_), .B2(new_n260_), .C1(new_n257_), .C2(new_n258_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT70), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n207_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n263_), .A2(new_n264_), .A3(KEYINPUT70), .A4(new_n206_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n205_), .A2(KEYINPUT36), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n265_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G127gat), .B(G134gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G113gat), .B(G120gat), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n273_), .A2(new_n274_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT80), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n275_), .A2(KEYINPUT80), .A3(new_n276_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT31), .ZN(new_n282_));
  OR2_X1    g081(.A1(new_n282_), .A2(KEYINPUT79), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G227gat), .A2(G233gat), .ZN(new_n284_));
  XOR2_X1   g083(.A(new_n284_), .B(KEYINPUT78), .Z(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(KEYINPUT30), .ZN(new_n286_));
  AND2_X1   g085(.A1(new_n283_), .A2(new_n286_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n283_), .A2(new_n286_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G15gat), .B(G43gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT77), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(G71gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(new_n235_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT76), .B(G176gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT22), .B(G169gat), .ZN(new_n294_));
  AOI22_X1  g093(.A1(new_n293_), .A2(new_n294_), .B1(G169gat), .B2(G176gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT75), .B(KEYINPUT23), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G183gat), .A2(G190gat), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n298_), .A2(KEYINPUT23), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(G183gat), .A2(G190gat), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n295_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n297_), .A2(KEYINPUT23), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n304_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT25), .B(G183gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(KEYINPUT26), .B(G190gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  OR2_X1    g107(.A1(G169gat), .A2(G176gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G169gat), .A2(G176gat), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n309_), .A2(KEYINPUT24), .A3(new_n310_), .ZN(new_n311_));
  OAI211_X1 g110(.A(new_n308_), .B(new_n311_), .C1(KEYINPUT24), .C2(new_n309_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n303_), .B1(new_n305_), .B2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n292_), .B(new_n313_), .ZN(new_n314_));
  OR3_X1    g113(.A1(new_n287_), .A2(new_n288_), .A3(new_n314_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n314_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n316_));
  AND2_X1   g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G78gat), .B(G106gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT87), .ZN(new_n319_));
  XOR2_X1   g118(.A(G22gat), .B(G50gat), .Z(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G155gat), .A2(G162gat), .ZN(new_n323_));
  OR2_X1    g122(.A1(new_n323_), .A2(KEYINPUT1), .ZN(new_n324_));
  NOR2_X1   g123(.A1(G155gat), .A2(G162gat), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n323_), .A2(KEYINPUT1), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n324_), .A2(new_n326_), .A3(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G141gat), .A2(G148gat), .ZN(new_n329_));
  NOR2_X1   g128(.A1(G141gat), .A2(G148gat), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  AND3_X1   g130(.A1(new_n328_), .A2(new_n329_), .A3(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n326_), .A2(new_n323_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT2), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n329_), .A2(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n335_), .B1(new_n337_), .B2(KEYINPUT81), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n330_), .A2(KEYINPUT3), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT3), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n340_), .B1(G141gat), .B2(G148gat), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT81), .ZN(new_n342_));
  AOI22_X1  g141(.A1(new_n339_), .A2(new_n341_), .B1(new_n336_), .B2(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n333_), .B1(new_n338_), .B2(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(KEYINPUT82), .B1(new_n332_), .B2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n338_), .A2(new_n343_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n333_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT82), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n328_), .A2(new_n329_), .A3(new_n331_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n348_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(KEYINPUT29), .B1(new_n345_), .B2(new_n351_), .ZN(new_n352_));
  XOR2_X1   g151(.A(KEYINPUT83), .B(KEYINPUT28), .Z(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  AOI211_X1 g154(.A(KEYINPUT29), .B(new_n353_), .C1(new_n345_), .C2(new_n351_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G228gat), .A2(G233gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT85), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n345_), .A2(new_n351_), .A3(KEYINPUT29), .ZN(new_n361_));
  OR2_X1    g160(.A1(new_n361_), .A2(KEYINPUT84), .ZN(new_n362_));
  INV_X1    g161(.A(G197gat), .ZN(new_n363_));
  INV_X1    g162(.A(G204gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G197gat), .A2(G204gat), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n365_), .A2(KEYINPUT21), .A3(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G211gat), .B(G218gat), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT86), .ZN(new_n369_));
  OR3_X1    g168(.A1(new_n367_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n369_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n371_));
  AND2_X1   g170(.A1(new_n365_), .A2(new_n366_), .ZN(new_n372_));
  OR2_X1    g171(.A1(new_n372_), .A2(KEYINPUT21), .ZN(new_n373_));
  AND2_X1   g172(.A1(new_n367_), .A2(new_n368_), .ZN(new_n374_));
  AOI22_X1  g173(.A1(new_n370_), .A2(new_n371_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n375_), .B1(new_n361_), .B2(KEYINPUT84), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n360_), .B1(new_n362_), .B2(new_n376_), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT29), .B1(new_n332_), .B2(new_n344_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n370_), .A2(new_n371_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n373_), .A2(new_n374_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n378_), .A2(new_n381_), .A3(new_n360_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n357_), .B1(new_n377_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NOR3_X1   g184(.A1(new_n377_), .A2(new_n357_), .A3(new_n383_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n322_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n386_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n388_), .A2(new_n321_), .A3(new_n384_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n387_), .A2(new_n389_), .ZN(new_n390_));
  XOR2_X1   g189(.A(KEYINPUT94), .B(KEYINPUT4), .Z(new_n391_));
  NAND4_X1  g190(.A1(new_n281_), .A2(new_n345_), .A3(new_n351_), .A4(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G225gat), .A2(G233gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(KEYINPUT93), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n392_), .A2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n281_), .A2(new_n345_), .A3(new_n351_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n348_), .A2(new_n350_), .A3(new_n277_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT4), .ZN(new_n399_));
  OAI21_X1  g198(.A(KEYINPUT92), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT92), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n396_), .A2(new_n401_), .A3(KEYINPUT4), .A4(new_n397_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n395_), .B1(new_n400_), .B2(new_n402_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n398_), .A2(new_n394_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G1gat), .B(G29gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(G85gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT0), .B(G57gat), .ZN(new_n407_));
  XOR2_X1   g206(.A(new_n406_), .B(new_n407_), .Z(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NOR3_X1   g208(.A1(new_n403_), .A2(new_n404_), .A3(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT95), .ZN(new_n411_));
  OAI21_X1  g210(.A(KEYINPUT33), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n400_), .A2(new_n402_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n395_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n404_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n415_), .A2(new_n416_), .A3(new_n408_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT33), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n417_), .A2(KEYINPUT95), .A3(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G226gat), .A2(G233gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(KEYINPUT19), .ZN(new_n421_));
  OAI21_X1  g220(.A(KEYINPUT20), .B1(new_n313_), .B2(new_n381_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT88), .B(KEYINPUT24), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n423_), .A2(new_n309_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n424_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n301_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n423_), .A2(new_n310_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n427_), .A2(KEYINPUT89), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n309_), .B1(new_n427_), .B2(KEYINPUT89), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n425_), .B(new_n426_), .C1(new_n428_), .C2(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n295_), .B1(new_n305_), .B2(new_n302_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n375_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n421_), .B1(new_n422_), .B2(new_n432_), .ZN(new_n433_));
  XOR2_X1   g232(.A(G8gat), .B(G36gat), .Z(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(KEYINPUT18), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G64gat), .B(G92gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n421_), .B1(new_n313_), .B2(new_n381_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n430_), .A2(new_n375_), .A3(new_n431_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n438_), .A2(KEYINPUT20), .A3(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n433_), .A2(new_n437_), .A3(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT90), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n433_), .A2(KEYINPUT90), .A3(new_n440_), .A4(new_n437_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n433_), .A2(new_n440_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n437_), .ZN(new_n446_));
  AOI21_X1  g245(.A(KEYINPUT91), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT91), .ZN(new_n448_));
  AOI211_X1 g247(.A(new_n448_), .B(new_n437_), .C1(new_n433_), .C2(new_n440_), .ZN(new_n449_));
  OAI211_X1 g248(.A(new_n443_), .B(new_n444_), .C1(new_n447_), .C2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n394_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n413_), .A2(new_n452_), .A3(new_n392_), .ZN(new_n453_));
  AOI21_X1  g252(.A(KEYINPUT96), .B1(new_n396_), .B2(new_n397_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT96), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n394_), .B1(new_n398_), .B2(new_n455_), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n453_), .B(new_n409_), .C1(new_n454_), .C2(new_n456_), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n412_), .A2(new_n419_), .A3(new_n451_), .A4(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n437_), .A2(KEYINPUT32), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n433_), .A2(new_n459_), .A3(new_n440_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n421_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n439_), .A2(KEYINPUT20), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT97), .ZN(new_n463_));
  AOI22_X1  g262(.A1(new_n462_), .A2(new_n463_), .B1(new_n381_), .B2(new_n313_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n439_), .A2(KEYINPUT97), .A3(KEYINPUT20), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n461_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  NOR3_X1   g265(.A1(new_n422_), .A2(new_n432_), .A3(new_n421_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n408_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n469_));
  OAI221_X1 g268(.A(new_n460_), .B1(new_n468_), .B2(new_n459_), .C1(new_n469_), .C2(new_n410_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n390_), .B1(new_n458_), .B2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT27), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT98), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n472_), .B1(new_n441_), .B2(new_n473_), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n433_), .A2(KEYINPUT98), .A3(new_n440_), .A4(new_n437_), .ZN(new_n475_));
  AND2_X1   g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n446_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n477_));
  AOI22_X1  g276(.A1(new_n450_), .A2(new_n472_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n469_), .A2(new_n410_), .ZN(new_n479_));
  AND3_X1   g278(.A1(new_n478_), .A2(new_n479_), .A3(new_n390_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n317_), .B1(new_n471_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n478_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n482_), .A2(new_n390_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n479_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n317_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n272_), .B1(new_n481_), .B2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G1gat), .B(G8gat), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT72), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n488_), .B(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(G15gat), .ZN(new_n491_));
  INV_X1    g290(.A(G22gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G15gat), .A2(G22gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G1gat), .A2(G8gat), .ZN(new_n495_));
  AOI22_X1  g294(.A1(new_n493_), .A2(new_n494_), .B1(KEYINPUT14), .B2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n490_), .B(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G231gat), .A2(G233gat), .ZN(new_n498_));
  XOR2_X1   g297(.A(new_n498_), .B(KEYINPUT73), .Z(new_n499_));
  XNOR2_X1  g298(.A(new_n497_), .B(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(G71gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(G78gat), .ZN(new_n502_));
  INV_X1    g301(.A(G78gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(G71gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n502_), .A2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G57gat), .B(G64gat), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n505_), .B1(new_n506_), .B2(KEYINPUT11), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT66), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n508_), .B1(new_n506_), .B2(KEYINPUT11), .ZN(new_n509_));
  INV_X1    g308(.A(G64gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(G57gat), .ZN(new_n511_));
  INV_X1    g310(.A(G57gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(G64gat), .ZN(new_n513_));
  AND4_X1   g312(.A1(new_n508_), .A2(new_n511_), .A3(new_n513_), .A4(KEYINPUT11), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n507_), .B1(new_n509_), .B2(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n511_), .A2(new_n513_), .A3(KEYINPUT11), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT66), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n511_), .A2(new_n513_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT11), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n511_), .A2(new_n513_), .A3(new_n508_), .A4(KEYINPUT11), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n517_), .A2(new_n520_), .A3(new_n505_), .A4(new_n521_), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n515_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n500_), .B(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT17), .ZN(new_n525_));
  XOR2_X1   g324(.A(G127gat), .B(G155gat), .Z(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT16), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G183gat), .B(G211gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  OR3_X1    g328(.A1(new_n524_), .A2(new_n525_), .A3(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(KEYINPUT17), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n524_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G229gat), .A2(G233gat), .ZN(new_n535_));
  XOR2_X1   g334(.A(new_n490_), .B(new_n496_), .Z(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(new_n248_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n497_), .A2(new_n247_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n254_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n254_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n248_), .A2(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n535_), .B1(new_n539_), .B2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n537_), .A2(new_n538_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n542_), .B1(new_n535_), .B2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G113gat), .B(G141gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G169gat), .B(G197gat), .ZN(new_n546_));
  XOR2_X1   g345(.A(new_n545_), .B(new_n546_), .Z(new_n547_));
  OR2_X1    g346(.A1(new_n544_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n544_), .A2(new_n547_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G230gat), .A2(G233gat), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n242_), .A2(new_n523_), .ZN(new_n552_));
  AND2_X1   g351(.A1(new_n221_), .A2(new_n223_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n236_), .A2(new_n228_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n240_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(new_n227_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n239_), .A2(new_n240_), .A3(new_n233_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n515_), .A2(new_n522_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n558_), .A2(new_n225_), .A3(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n551_), .B1(new_n552_), .B2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n552_), .A2(new_n560_), .A3(KEYINPUT12), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT12), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n242_), .A2(new_n523_), .A3(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n561_), .B1(new_n565_), .B2(new_n551_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G120gat), .B(G148gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT5), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G176gat), .B(G204gat), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n568_), .B(new_n569_), .Z(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n571_), .A2(KEYINPUT67), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n566_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n566_), .A2(new_n573_), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n576_), .A2(KEYINPUT13), .ZN(new_n577_));
  AND3_X1   g376(.A1(new_n574_), .A2(KEYINPUT13), .A3(new_n575_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  AND4_X1   g378(.A1(new_n487_), .A2(new_n534_), .A3(new_n550_), .A4(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n202_), .B1(new_n580_), .B2(new_n484_), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n581_), .B(KEYINPUT99), .Z(new_n582_));
  XOR2_X1   g381(.A(new_n550_), .B(KEYINPUT74), .Z(new_n583_));
  NAND3_X1  g382(.A1(new_n272_), .A2(KEYINPUT71), .A3(KEYINPUT37), .ZN(new_n584_));
  AOI22_X1  g383(.A1(new_n267_), .A2(new_n268_), .B1(new_n265_), .B2(new_n270_), .ZN(new_n585_));
  OR2_X1    g384(.A1(KEYINPUT71), .A2(KEYINPUT37), .ZN(new_n586_));
  NAND2_X1  g385(.A1(KEYINPUT71), .A2(KEYINPUT37), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n585_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n584_), .A2(new_n579_), .A3(new_n534_), .A4(new_n588_), .ZN(new_n589_));
  AOI211_X1 g388(.A(new_n583_), .B(new_n589_), .C1(new_n481_), .C2(new_n486_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n590_), .A2(new_n202_), .A3(new_n484_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT38), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n591_), .B1(KEYINPUT100), .B2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT100), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n593_), .B1(new_n594_), .B2(KEYINPUT38), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n591_), .A2(KEYINPUT100), .A3(new_n592_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n582_), .A2(new_n595_), .A3(new_n596_), .ZN(G1324gat));
  INV_X1    g396(.A(G8gat), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n590_), .A2(new_n598_), .A3(new_n482_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT39), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n580_), .A2(new_n482_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n600_), .B1(new_n601_), .B2(G8gat), .ZN(new_n602_));
  AOI211_X1 g401(.A(KEYINPUT39), .B(new_n598_), .C1(new_n580_), .C2(new_n482_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n599_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT40), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(G1325gat));
  INV_X1    g405(.A(new_n317_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n580_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(G15gat), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(KEYINPUT101), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT101), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n608_), .A2(new_n611_), .A3(G15gat), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT41), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n590_), .A2(new_n491_), .A3(new_n607_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n610_), .A2(KEYINPUT41), .A3(new_n612_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n615_), .A2(new_n616_), .A3(new_n617_), .ZN(G1326gat));
  XNOR2_X1  g417(.A(new_n390_), .B(KEYINPUT102), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n492_), .B1(new_n580_), .B2(new_n620_), .ZN(new_n621_));
  XOR2_X1   g420(.A(KEYINPUT103), .B(KEYINPUT42), .Z(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n590_), .A2(new_n492_), .A3(new_n620_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(G1327gat));
  AOI21_X1  g424(.A(new_n583_), .B1(new_n481_), .B2(new_n486_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n579_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n272_), .A2(new_n533_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n626_), .A2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT105), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT105), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n626_), .A2(new_n632_), .A3(new_n629_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n631_), .A2(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(G29gat), .B1(new_n634_), .B2(new_n484_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n550_), .ZN(new_n636_));
  NOR3_X1   g435(.A1(new_n627_), .A2(new_n534_), .A3(new_n636_), .ZN(new_n637_));
  AND3_X1   g436(.A1(new_n585_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n587_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT104), .ZN(new_n641_));
  AOI221_X4 g440(.A(new_n640_), .B1(new_n641_), .B2(KEYINPUT43), .C1(new_n481_), .C2(new_n486_), .ZN(new_n642_));
  OAI21_X1  g441(.A(KEYINPUT43), .B1(new_n640_), .B2(new_n641_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n481_), .A2(new_n486_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n584_), .A2(new_n588_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n643_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n637_), .B1(new_n642_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT44), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  OAI211_X1 g448(.A(KEYINPUT44), .B(new_n637_), .C1(new_n642_), .C2(new_n646_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n484_), .A2(G29gat), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n635_), .B1(new_n651_), .B2(new_n652_), .ZN(G1328gat));
  NAND3_X1  g452(.A1(new_n649_), .A2(new_n482_), .A3(new_n650_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(G36gat), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n478_), .A2(G36gat), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n631_), .A2(new_n633_), .A3(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT45), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n655_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT46), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n655_), .A2(new_n658_), .A3(KEYINPUT46), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1329gat));
  NAND4_X1  g462(.A1(new_n649_), .A2(G43gat), .A3(new_n607_), .A4(new_n650_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n631_), .A2(new_n607_), .A3(new_n633_), .ZN(new_n665_));
  INV_X1    g464(.A(G43gat), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n664_), .A2(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g468(.A1(new_n651_), .A2(new_n390_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(G50gat), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n619_), .A2(G50gat), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n672_), .B(KEYINPUT106), .Z(new_n673_));
  NAND2_X1  g472(.A1(new_n634_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n671_), .A2(new_n674_), .ZN(G1331gat));
  AND4_X1   g474(.A1(new_n487_), .A2(new_n534_), .A3(new_n627_), .A4(new_n583_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(KEYINPUT107), .A2(G57gat), .ZN(new_n677_));
  AND2_X1   g476(.A1(KEYINPUT107), .A2(G57gat), .ZN(new_n678_));
  OAI211_X1 g477(.A(new_n676_), .B(new_n484_), .C1(new_n677_), .C2(new_n678_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT108), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n644_), .A2(new_n636_), .A3(new_n627_), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n681_), .A2(new_n533_), .A3(new_n645_), .ZN(new_n682_));
  AOI21_X1  g481(.A(G57gat), .B1(new_n682_), .B2(new_n484_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n680_), .A2(new_n683_), .ZN(G1332gat));
  NAND3_X1  g483(.A1(new_n682_), .A2(new_n510_), .A3(new_n482_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT48), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n676_), .A2(new_n482_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n686_), .B1(new_n687_), .B2(G64gat), .ZN(new_n688_));
  AOI211_X1 g487(.A(KEYINPUT48), .B(new_n510_), .C1(new_n676_), .C2(new_n482_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n685_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT109), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n690_), .B(new_n691_), .ZN(G1333gat));
  AOI21_X1  g491(.A(new_n501_), .B1(new_n676_), .B2(new_n607_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT49), .Z(new_n694_));
  NAND3_X1  g493(.A1(new_n682_), .A2(new_n501_), .A3(new_n607_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(G1334gat));
  AOI21_X1  g495(.A(new_n503_), .B1(new_n676_), .B2(new_n620_), .ZN(new_n697_));
  XOR2_X1   g496(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n698_));
  XNOR2_X1  g497(.A(new_n697_), .B(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n682_), .A2(new_n503_), .A3(new_n620_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1335gat));
  OR2_X1    g500(.A1(new_n642_), .A2(new_n646_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n627_), .A2(new_n533_), .A3(new_n636_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT111), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(G85gat), .B1(new_n705_), .B2(new_n479_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n681_), .A2(new_n628_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n707_), .A2(new_n209_), .A3(new_n484_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n708_), .ZN(G1336gat));
  AOI21_X1  g508(.A(G92gat), .B1(new_n707_), .B2(new_n482_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n705_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n478_), .A2(new_n210_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT112), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n710_), .B1(new_n711_), .B2(new_n713_), .ZN(G1337gat));
  NAND3_X1  g513(.A1(new_n707_), .A2(new_n607_), .A3(new_n216_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n702_), .A2(new_n607_), .A3(new_n704_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n718_), .B2(G99gat), .ZN(new_n719_));
  NOR2_X1   g518(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n719_), .B(new_n720_), .ZN(G1338gat));
  NAND3_X1  g520(.A1(new_n707_), .A2(new_n217_), .A3(new_n390_), .ZN(new_n722_));
  OAI211_X1 g521(.A(new_n390_), .B(new_n704_), .C1(new_n642_), .C2(new_n646_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT52), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n723_), .A2(new_n724_), .A3(G106gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n723_), .B2(G106gat), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n722_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g527(.A1(new_n566_), .A2(new_n571_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n550_), .A2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n551_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n562_), .A2(new_n731_), .A3(new_n564_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT114), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n562_), .A2(KEYINPUT114), .A3(new_n731_), .A4(new_n564_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n565_), .A2(new_n551_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(KEYINPUT55), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT55), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n565_), .A2(new_n738_), .A3(new_n551_), .ZN(new_n739_));
  AOI221_X4 g538(.A(KEYINPUT115), .B1(new_n734_), .B2(new_n735_), .C1(new_n737_), .C2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT115), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n737_), .A2(new_n739_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n734_), .A2(new_n735_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n741_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n570_), .B1(new_n740_), .B2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT56), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n738_), .B1(new_n565_), .B2(new_n551_), .ZN(new_n748_));
  AOI211_X1 g547(.A(KEYINPUT55), .B(new_n731_), .C1(new_n562_), .C2(new_n564_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n743_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT115), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n742_), .A2(new_n741_), .A3(new_n743_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n753_), .A2(KEYINPUT56), .A3(new_n570_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n730_), .B1(new_n747_), .B2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT117), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n543_), .A2(new_n540_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT116), .ZN(new_n758_));
  INV_X1    g557(.A(new_n541_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n757_), .A2(new_n758_), .A3(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(KEYINPUT116), .B1(new_n539_), .B2(new_n541_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n535_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n547_), .B1(new_n543_), .B2(new_n535_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n756_), .B1(new_n762_), .B2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n535_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n758_), .B1(new_n757_), .B2(new_n759_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n539_), .A2(KEYINPUT116), .A3(new_n541_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n766_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n769_), .A2(KEYINPUT117), .A3(new_n763_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n765_), .A2(new_n770_), .A3(new_n549_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n771_), .A2(new_n576_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n585_), .B1(new_n755_), .B2(new_n772_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(KEYINPUT118), .A2(KEYINPUT57), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n774_), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n585_), .B(new_n776_), .C1(new_n755_), .C2(new_n772_), .ZN(new_n777_));
  AND4_X1   g576(.A1(new_n549_), .A2(new_n765_), .A3(new_n770_), .A4(new_n729_), .ZN(new_n778_));
  AOI21_X1  g577(.A(KEYINPUT56), .B1(new_n753_), .B2(new_n570_), .ZN(new_n779_));
  AOI211_X1 g578(.A(new_n746_), .B(new_n571_), .C1(new_n751_), .C2(new_n752_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n778_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT58), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  OAI211_X1 g582(.A(KEYINPUT58), .B(new_n778_), .C1(new_n779_), .C2(new_n780_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n783_), .A2(new_n645_), .A3(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n775_), .A2(new_n777_), .A3(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(new_n533_), .ZN(new_n787_));
  NOR3_X1   g586(.A1(new_n638_), .A2(new_n639_), .A3(new_n533_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT54), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n788_), .A2(new_n789_), .A3(new_n579_), .A4(new_n583_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n550_), .B(KEYINPUT74), .ZN(new_n791_));
  OAI21_X1  g590(.A(KEYINPUT54), .B1(new_n589_), .B2(new_n791_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n790_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n787_), .A2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT59), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n483_), .A2(new_n484_), .A3(new_n607_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n795_), .A2(new_n796_), .A3(new_n798_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(KEYINPUT120), .B(G113gat), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n583_), .A2(new_n800_), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n550_), .A2(new_n729_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n802_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n772_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n272_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n784_), .A2(new_n645_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n747_), .A2(new_n754_), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT58), .B1(new_n807_), .B2(new_n778_), .ZN(new_n808_));
  OAI22_X1  g607(.A1(new_n805_), .A2(new_n776_), .B1(new_n806_), .B2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n777_), .ZN(new_n810_));
  OAI21_X1  g609(.A(KEYINPUT119), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT119), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n775_), .A2(new_n785_), .A3(new_n812_), .A4(new_n777_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n811_), .A2(new_n533_), .A3(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n797_), .B1(new_n814_), .B2(new_n794_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n799_), .B(new_n801_), .C1(new_n815_), .C2(new_n796_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(G113gat), .B1(new_n815_), .B2(new_n550_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n817_), .A2(new_n818_), .ZN(G1340gat));
  INV_X1    g618(.A(KEYINPUT60), .ZN(new_n820_));
  AOI21_X1  g619(.A(G120gat), .B1(new_n627_), .B2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(G120gat), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n823_), .A2(KEYINPUT60), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n822_), .B1(KEYINPUT121), .B2(new_n824_), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n815_), .B(new_n825_), .C1(KEYINPUT121), .C2(new_n822_), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n627_), .B(new_n799_), .C1(new_n815_), .C2(new_n796_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n826_), .B1(new_n828_), .B2(new_n823_), .ZN(G1341gat));
  INV_X1    g628(.A(G127gat), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n815_), .A2(new_n830_), .A3(new_n534_), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n534_), .B(new_n799_), .C1(new_n815_), .C2(new_n796_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n831_), .B1(new_n833_), .B2(new_n830_), .ZN(G1342gat));
  INV_X1    g633(.A(G134gat), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n815_), .A2(new_n835_), .A3(new_n272_), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n645_), .B(new_n799_), .C1(new_n815_), .C2(new_n796_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n836_), .B1(new_n838_), .B2(new_n835_), .ZN(G1343gat));
  INV_X1    g638(.A(new_n390_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n482_), .A2(new_n840_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n841_), .A2(new_n484_), .A3(new_n317_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n842_), .B1(new_n814_), .B2(new_n794_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n550_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n627_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g646(.A(KEYINPUT61), .B(G155gat), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT122), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n850_), .B1(new_n843_), .B2(new_n534_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n534_), .B1(new_n786_), .B2(KEYINPUT119), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n793_), .B1(new_n852_), .B2(new_n813_), .ZN(new_n853_));
  NOR4_X1   g652(.A1(new_n853_), .A2(KEYINPUT122), .A3(new_n533_), .A4(new_n842_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n849_), .B1(new_n851_), .B2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n814_), .A2(new_n794_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n842_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n856_), .A2(new_n534_), .A3(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(KEYINPUT122), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n843_), .A2(new_n850_), .A3(new_n534_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n859_), .A2(new_n860_), .A3(new_n848_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n855_), .A2(new_n861_), .ZN(G1346gat));
  INV_X1    g661(.A(new_n843_), .ZN(new_n863_));
  INV_X1    g662(.A(G162gat), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n863_), .A2(new_n864_), .A3(new_n640_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT123), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n853_), .A2(new_n585_), .A3(new_n842_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n866_), .B1(new_n867_), .B2(G162gat), .ZN(new_n868_));
  OAI211_X1 g667(.A(KEYINPUT123), .B(new_n864_), .C1(new_n863_), .C2(new_n585_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n865_), .B1(new_n868_), .B2(new_n869_), .ZN(G1347gat));
  NAND2_X1  g669(.A1(new_n485_), .A2(new_n482_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n619_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n795_), .A2(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(G169gat), .B1(new_n875_), .B2(new_n636_), .ZN(new_n876_));
  AND2_X1   g675(.A1(new_n876_), .A2(KEYINPUT62), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n876_), .A2(KEYINPUT62), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n550_), .A2(new_n294_), .ZN(new_n879_));
  XOR2_X1   g678(.A(new_n879_), .B(KEYINPUT124), .Z(new_n880_));
  OAI22_X1  g679(.A1(new_n877_), .A2(new_n878_), .B1(new_n875_), .B2(new_n880_), .ZN(G1348gat));
  AOI21_X1  g680(.A(new_n390_), .B1(new_n814_), .B2(new_n794_), .ZN(new_n882_));
  AND3_X1   g681(.A1(new_n872_), .A2(G176gat), .A3(new_n627_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT125), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n882_), .A2(KEYINPUT125), .A3(new_n883_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n873_), .B1(new_n787_), .B2(new_n794_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(new_n627_), .ZN(new_n889_));
  AOI22_X1  g688(.A1(new_n886_), .A2(new_n887_), .B1(new_n293_), .B2(new_n889_), .ZN(G1349gat));
  NOR2_X1   g689(.A1(new_n871_), .A2(new_n533_), .ZN(new_n891_));
  AOI21_X1  g690(.A(G183gat), .B1(new_n882_), .B2(new_n891_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n533_), .A2(new_n306_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n806_), .ZN(new_n894_));
  AOI22_X1  g693(.A1(new_n894_), .A2(new_n783_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n534_), .B1(new_n895_), .B2(new_n777_), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n874_), .B(new_n893_), .C1(new_n896_), .C2(new_n793_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(KEYINPUT126), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT126), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n888_), .A2(new_n899_), .A3(new_n893_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n900_), .ZN(new_n901_));
  OAI21_X1  g700(.A(KEYINPUT127), .B1(new_n892_), .B2(new_n901_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n856_), .A2(new_n840_), .A3(new_n891_), .ZN(new_n903_));
  INV_X1    g702(.A(G183gat), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n899_), .B1(new_n888_), .B2(new_n893_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n793_), .B1(new_n786_), .B2(new_n533_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n893_), .ZN(new_n908_));
  NOR4_X1   g707(.A1(new_n907_), .A2(KEYINPUT126), .A3(new_n873_), .A4(new_n908_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n906_), .A2(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT127), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n905_), .A2(new_n910_), .A3(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n902_), .A2(new_n912_), .ZN(G1350gat));
  OAI21_X1  g712(.A(G190gat), .B1(new_n875_), .B2(new_n640_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n888_), .A2(new_n307_), .A3(new_n272_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(G1351gat));
  NOR4_X1   g715(.A1(new_n607_), .A2(new_n840_), .A3(new_n484_), .A4(new_n478_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n856_), .A2(new_n917_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  AOI21_X1  g718(.A(G197gat), .B1(new_n919_), .B2(new_n550_), .ZN(new_n920_));
  NOR3_X1   g719(.A1(new_n918_), .A2(new_n363_), .A3(new_n636_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n920_), .A2(new_n921_), .ZN(G1352gat));
  NAND3_X1  g721(.A1(new_n919_), .A2(new_n364_), .A3(new_n627_), .ZN(new_n923_));
  OAI21_X1  g722(.A(G204gat), .B1(new_n918_), .B2(new_n579_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(new_n924_), .ZN(G1353gat));
  XNOR2_X1  g724(.A(KEYINPUT63), .B(G211gat), .ZN(new_n926_));
  NOR3_X1   g725(.A1(new_n918_), .A2(new_n533_), .A3(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n919_), .A2(new_n534_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n927_), .B1(new_n928_), .B2(new_n929_), .ZN(G1354gat));
  OR3_X1    g729(.A1(new_n918_), .A2(G218gat), .A3(new_n585_), .ZN(new_n931_));
  OAI21_X1  g730(.A(G218gat), .B1(new_n918_), .B2(new_n640_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(new_n932_), .ZN(G1355gat));
endmodule


