//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 1 1 0 0 1 0 0 0 1 1 0 0 1 1 1 1 1 0 1 0 0 1 1 0 0 0 1 1 1 0 1 0 0 1 0 0 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n703_, new_n704_, new_n705_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n742_,
    new_n743_, new_n744_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n833_, new_n834_, new_n835_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n842_, new_n844_, new_n845_, new_n847_, new_n848_,
    new_n849_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n884_, new_n885_, new_n887_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_, new_n910_,
    new_n911_;
  INV_X1    g000(.A(KEYINPUT100), .ZN(new_n202_));
  XOR2_X1   g001(.A(G197gat), .B(G204gat), .Z(new_n203_));
  INV_X1    g002(.A(KEYINPUT85), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n203_), .A2(new_n204_), .A3(KEYINPUT21), .ZN(new_n205_));
  XOR2_X1   g004(.A(G211gat), .B(G218gat), .Z(new_n206_));
  OR2_X1    g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n206_), .ZN(new_n208_));
  OR2_X1    g007(.A1(new_n203_), .A2(KEYINPUT21), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n207_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n214_), .A2(KEYINPUT23), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n213_), .B(KEYINPUT81), .ZN(new_n216_));
  AOI211_X1 g015(.A(new_n212_), .B(new_n215_), .C1(new_n216_), .C2(KEYINPUT23), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT22), .B(G169gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n219_), .A2(KEYINPUT82), .ZN(new_n220_));
  INV_X1    g019(.A(G176gat), .ZN(new_n221_));
  INV_X1    g020(.A(G169gat), .ZN(new_n222_));
  AND2_X1   g021(.A1(new_n222_), .A2(KEYINPUT22), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT82), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n221_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n218_), .B1(new_n220_), .B2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT23), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n214_), .A2(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n228_), .B1(new_n216_), .B2(new_n227_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT26), .B(G190gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT79), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT25), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n231_), .B1(new_n232_), .B2(G183gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT25), .B(G183gat), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n230_), .B(new_n233_), .C1(new_n234_), .C2(new_n231_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(G169gat), .A2(G176gat), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT80), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(KEYINPUT80), .B1(G169gat), .B2(G176gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT24), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n238_), .A2(KEYINPUT24), .A3(new_n239_), .A4(new_n218_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n235_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  OAI22_X1  g043(.A1(new_n217_), .A2(new_n226_), .B1(new_n229_), .B2(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT20), .B1(new_n211_), .B2(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n215_), .B1(new_n216_), .B2(KEYINPUT23), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n236_), .A2(new_n241_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n230_), .A2(new_n234_), .ZN(new_n249_));
  AND3_X1   g048(.A1(new_n249_), .A2(new_n243_), .A3(KEYINPUT90), .ZN(new_n250_));
  AOI21_X1  g049(.A(KEYINPUT90), .B1(new_n249_), .B2(new_n243_), .ZN(new_n251_));
  OAI211_X1 g050(.A(new_n247_), .B(new_n248_), .C1(new_n250_), .C2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n219_), .A2(new_n221_), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n218_), .B(new_n253_), .C1(new_n229_), .C2(new_n212_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n210_), .B1(new_n252_), .B2(new_n254_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n246_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G226gat), .A2(G233gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT19), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT89), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n256_), .A2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n252_), .A2(new_n210_), .A3(new_n254_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT97), .ZN(new_n263_));
  AND3_X1   g062(.A1(new_n262_), .A2(new_n263_), .A3(KEYINPUT20), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n263_), .B1(new_n262_), .B2(KEYINPUT20), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n211_), .A2(new_n245_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NOR3_X1   g066(.A1(new_n264_), .A2(new_n265_), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n258_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n261_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G8gat), .B(G36gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT18), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G64gat), .B(G92gat), .ZN(new_n274_));
  XOR2_X1   g073(.A(new_n273_), .B(new_n274_), .Z(new_n275_));
  OAI21_X1  g074(.A(new_n202_), .B1(new_n271_), .B2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n275_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n270_), .A2(KEYINPUT100), .A3(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n276_), .A2(new_n278_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n259_), .B1(new_n246_), .B2(new_n255_), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n266_), .A2(KEYINPUT20), .A3(new_n262_), .A4(new_n269_), .ZN(new_n281_));
  AND3_X1   g080(.A1(new_n280_), .A2(new_n281_), .A3(new_n275_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT27), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n275_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n282_), .A2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT101), .B1(new_n286_), .B2(KEYINPUT27), .ZN(new_n287_));
  OR3_X1    g086(.A1(new_n286_), .A2(KEYINPUT101), .A3(KEYINPUT27), .ZN(new_n288_));
  AOI22_X1  g087(.A1(new_n279_), .A2(new_n284_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G15gat), .B(G43gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT83), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(G71gat), .ZN(new_n292_));
  INV_X1    g091(.A(G99gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  OR2_X1    g093(.A1(new_n294_), .A2(new_n245_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G127gat), .B(G134gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G113gat), .B(G120gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n294_), .A2(new_n245_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n295_), .A2(new_n298_), .A3(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G227gat), .A2(G233gat), .ZN(new_n302_));
  XOR2_X1   g101(.A(new_n302_), .B(KEYINPUT84), .Z(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT30), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT31), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n298_), .B1(new_n295_), .B2(new_n299_), .ZN(new_n307_));
  OR3_X1    g106(.A1(new_n301_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n306_), .B1(new_n301_), .B2(new_n307_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G141gat), .A2(G148gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT2), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n313_));
  NOR2_X1   g112(.A1(G141gat), .A2(G148gat), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT3), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n312_), .A2(new_n313_), .A3(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G155gat), .B(G162gat), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(G155gat), .A2(G162gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G155gat), .A2(G162gat), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n321_), .B1(KEYINPUT1), .B2(new_n322_), .ZN(new_n323_));
  OR2_X1    g122(.A1(new_n322_), .A2(KEYINPUT1), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n311_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n326_), .A2(new_n314_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n325_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n320_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT4), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n296_), .A2(new_n297_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n296_), .A2(new_n297_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n329_), .A2(new_n330_), .A3(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G225gat), .A2(G233gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT92), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(new_n336_), .ZN(new_n337_));
  AND2_X1   g136(.A1(new_n325_), .A2(new_n327_), .ZN(new_n338_));
  AND2_X1   g137(.A1(new_n316_), .A2(new_n313_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n318_), .B1(new_n339_), .B2(new_n312_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n333_), .B1(new_n338_), .B2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n320_), .A2(new_n328_), .A3(new_n298_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n341_), .A2(new_n342_), .A3(KEYINPUT91), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT91), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n320_), .A2(new_n344_), .A3(new_n328_), .A4(new_n298_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n337_), .B1(new_n346_), .B2(KEYINPUT4), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT93), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT93), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n330_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n349_), .B1(new_n350_), .B2(new_n337_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n346_), .A2(new_n335_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n348_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n353_));
  XOR2_X1   g152(.A(G1gat), .B(G29gat), .Z(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G57gat), .B(G85gat), .ZN(new_n357_));
  XOR2_X1   g156(.A(new_n356_), .B(new_n357_), .Z(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n353_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT98), .ZN(new_n361_));
  AOI22_X1  g160(.A1(new_n347_), .A2(KEYINPUT93), .B1(new_n346_), .B2(new_n335_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n362_), .A2(new_n358_), .A3(new_n351_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n360_), .A2(new_n361_), .A3(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n353_), .A2(KEYINPUT98), .A3(new_n359_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n310_), .A2(new_n367_), .ZN(new_n368_));
  AND2_X1   g167(.A1(new_n329_), .A2(KEYINPUT29), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n369_), .A2(new_n210_), .ZN(new_n370_));
  INV_X1    g169(.A(G228gat), .ZN(new_n371_));
  INV_X1    g170(.A(G233gat), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n370_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  OAI211_X1 g172(.A(G228gat), .B(G233gat), .C1(new_n369_), .C2(new_n210_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G78gat), .B(G106gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT86), .ZN(new_n378_));
  INV_X1    g177(.A(new_n376_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n373_), .A2(new_n374_), .A3(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n377_), .A2(new_n378_), .A3(new_n380_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n329_), .A2(KEYINPUT29), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT28), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G22gat), .B(G50gat), .ZN(new_n384_));
  AND2_X1   g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n383_), .A2(new_n384_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n381_), .B(new_n388_), .C1(new_n378_), .C2(new_n377_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT88), .ZN(new_n390_));
  OR2_X1    g189(.A1(new_n380_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n380_), .A2(new_n390_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n391_), .A2(new_n392_), .A3(new_n387_), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n373_), .A2(KEYINPUT87), .A3(new_n374_), .ZN(new_n394_));
  AOI21_X1  g193(.A(KEYINPUT87), .B1(new_n373_), .B2(new_n374_), .ZN(new_n395_));
  NOR3_X1   g194(.A1(new_n394_), .A2(new_n395_), .A3(new_n379_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n389_), .B1(new_n393_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n289_), .A2(new_n368_), .A3(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n275_), .A2(KEYINPUT32), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n280_), .A2(new_n281_), .A3(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n400_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n401_), .B1(new_n270_), .B2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n364_), .A2(new_n403_), .A3(new_n365_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(KEYINPUT99), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT99), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n364_), .A2(new_n403_), .A3(new_n406_), .A4(new_n365_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT33), .ZN(new_n408_));
  OR2_X1    g207(.A1(new_n363_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n363_), .A2(new_n408_), .ZN(new_n410_));
  OR2_X1    g209(.A1(new_n346_), .A2(KEYINPUT95), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n346_), .A2(KEYINPUT95), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n411_), .A2(new_n336_), .A3(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n350_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT96), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n334_), .A2(new_n335_), .ZN(new_n416_));
  AND3_X1   g215(.A1(new_n414_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n415_), .B1(new_n414_), .B2(new_n416_), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n413_), .B(new_n359_), .C1(new_n417_), .C2(new_n418_), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n409_), .A2(new_n286_), .A3(new_n410_), .A4(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n405_), .A2(new_n407_), .A3(new_n420_), .ZN(new_n421_));
  AND2_X1   g220(.A1(new_n397_), .A2(new_n366_), .ZN(new_n422_));
  AOI22_X1  g221(.A1(new_n398_), .A2(new_n421_), .B1(new_n422_), .B2(new_n289_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n310_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n399_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT70), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G29gat), .B(G36gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G43gat), .B(G50gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n427_), .B(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(KEYINPUT69), .B(KEYINPUT15), .ZN(new_n430_));
  XOR2_X1   g229(.A(new_n429_), .B(new_n430_), .Z(new_n431_));
  INV_X1    g230(.A(G106gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n293_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT7), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT66), .B1(G99gat), .B2(G106gat), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT7), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NOR3_X1   g236(.A1(KEYINPUT66), .A2(G99gat), .A3(G106gat), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n434_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G99gat), .A2(G106gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(KEYINPUT6), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT6), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n442_), .A2(G99gat), .A3(G106gat), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n441_), .A2(new_n443_), .A3(KEYINPUT65), .ZN(new_n444_));
  AOI21_X1  g243(.A(KEYINPUT65), .B1(new_n441_), .B2(new_n443_), .ZN(new_n445_));
  NOR3_X1   g244(.A1(new_n439_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G85gat), .B(G92gat), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n447_), .A2(KEYINPUT8), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT8), .ZN(new_n450_));
  AOI22_X1  g249(.A1(new_n441_), .A2(new_n443_), .B1(new_n433_), .B2(KEYINPUT7), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT66), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n452_), .A2(new_n293_), .A3(new_n432_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n453_), .A2(new_n436_), .A3(new_n435_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n447_), .B1(new_n451_), .B2(new_n454_), .ZN(new_n455_));
  OAI22_X1  g254(.A1(new_n446_), .A2(new_n449_), .B1(new_n450_), .B2(new_n455_), .ZN(new_n456_));
  OR2_X1    g255(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n457_), .A2(KEYINPUT64), .A3(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(KEYINPUT64), .B1(new_n457_), .B2(new_n458_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n432_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n444_), .A2(new_n445_), .ZN(new_n463_));
  INV_X1    g262(.A(G85gat), .ZN(new_n464_));
  INV_X1    g263(.A(G92gat), .ZN(new_n465_));
  NOR3_X1   g264(.A1(new_n464_), .A2(new_n465_), .A3(KEYINPUT9), .ZN(new_n466_));
  INV_X1    g265(.A(new_n447_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n466_), .B1(new_n467_), .B2(KEYINPUT9), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n462_), .A2(new_n463_), .A3(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n456_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n431_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n441_), .A2(new_n443_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n454_), .A2(new_n472_), .A3(new_n434_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(new_n467_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT65), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n442_), .B1(G99gat), .B2(G106gat), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n440_), .A2(KEYINPUT6), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n475_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n441_), .A2(new_n443_), .A3(KEYINPUT65), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n478_), .A2(new_n479_), .A3(new_n434_), .A4(new_n454_), .ZN(new_n480_));
  AOI22_X1  g279(.A1(KEYINPUT8), .A2(new_n474_), .B1(new_n480_), .B2(new_n448_), .ZN(new_n481_));
  AND3_X1   g280(.A1(new_n462_), .A2(new_n463_), .A3(new_n468_), .ZN(new_n482_));
  OAI21_X1  g281(.A(KEYINPUT67), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT67), .ZN(new_n484_));
  INV_X1    g283(.A(new_n439_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n449_), .B1(new_n463_), .B2(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n450_), .B1(new_n473_), .B2(new_n467_), .ZN(new_n487_));
  OAI211_X1 g286(.A(new_n484_), .B(new_n469_), .C1(new_n486_), .C2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n483_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n429_), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n426_), .B(new_n471_), .C1(new_n489_), .C2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G232gat), .A2(G233gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n488_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n484_), .B1(new_n456_), .B2(new_n469_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  AOI22_X1  g296(.A1(new_n497_), .A2(new_n429_), .B1(new_n431_), .B2(new_n470_), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n491_), .B(new_n494_), .C1(new_n498_), .C2(KEYINPUT35), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G190gat), .B(G218gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G134gat), .B(G162gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n502_), .A2(KEYINPUT36), .ZN(new_n503_));
  OR2_X1    g302(.A1(new_n491_), .A2(new_n494_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n499_), .A2(new_n503_), .A3(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  XOR2_X1   g305(.A(new_n502_), .B(KEYINPUT36), .Z(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT71), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n509_), .B1(new_n499_), .B2(new_n504_), .ZN(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT37), .B1(new_n506_), .B2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n499_), .A2(new_n504_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(new_n507_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(new_n505_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n511_), .B1(KEYINPUT37), .B2(new_n514_), .ZN(new_n515_));
  XOR2_X1   g314(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT75), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G127gat), .B(G155gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G183gat), .B(G211gat), .ZN(new_n520_));
  XOR2_X1   g319(.A(new_n519_), .B(new_n520_), .Z(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT17), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G57gat), .B(G64gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT11), .ZN(new_n524_));
  XOR2_X1   g323(.A(G71gat), .B(G78gat), .Z(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n523_), .A2(KEYINPUT11), .ZN(new_n527_));
  OR2_X1    g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  OR2_X1    g327(.A1(new_n524_), .A2(new_n525_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G231gat), .A2(G233gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(KEYINPUT72), .B(G8gat), .ZN(new_n533_));
  INV_X1    g332(.A(G1gat), .ZN(new_n534_));
  OAI21_X1  g333(.A(KEYINPUT14), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G15gat), .B(G22gat), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT73), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT73), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n535_), .A2(new_n539_), .A3(new_n536_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G1gat), .B(G8gat), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n538_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n541_), .B1(new_n538_), .B2(new_n540_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n532_), .B(new_n545_), .ZN(new_n546_));
  OR2_X1    g345(.A1(new_n522_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n546_), .A2(KEYINPUT17), .A3(new_n521_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n515_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT76), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  XOR2_X1   g352(.A(G113gat), .B(G141gat), .Z(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT78), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G169gat), .B(G197gat), .ZN(new_n556_));
  XOR2_X1   g355(.A(new_n555_), .B(new_n556_), .Z(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n431_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G229gat), .A2(G233gat), .ZN(new_n560_));
  INV_X1    g359(.A(new_n544_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n561_), .A2(new_n542_), .A3(new_n429_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n559_), .A2(new_n560_), .A3(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(KEYINPUT77), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n560_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n429_), .B1(new_n561_), .B2(new_n542_), .ZN(new_n567_));
  NOR3_X1   g366(.A1(new_n543_), .A2(new_n544_), .A3(new_n490_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n566_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT77), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n559_), .A2(new_n570_), .A3(new_n562_), .A4(new_n560_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n558_), .B1(new_n565_), .B2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n564_), .A2(new_n569_), .A3(new_n571_), .A4(new_n557_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n530_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n470_), .A2(new_n579_), .A3(KEYINPUT12), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n530_), .B1(new_n483_), .B2(new_n488_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n580_), .B1(new_n581_), .B2(KEYINPUT12), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n483_), .A2(new_n530_), .A3(new_n488_), .ZN(new_n584_));
  INV_X1    g383(.A(G230gat), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n585_), .A2(new_n372_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n584_), .A2(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n579_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(new_n584_), .ZN(new_n590_));
  AOI22_X1  g389(.A1(new_n583_), .A2(new_n588_), .B1(new_n586_), .B2(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G120gat), .B(G148gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT5), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G176gat), .B(G204gat), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n593_), .B(new_n594_), .Z(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n591_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n591_), .A2(new_n596_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT13), .ZN(new_n600_));
  OAI211_X1 g399(.A(new_n598_), .B(new_n599_), .C1(KEYINPUT68), .C2(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(KEYINPUT68), .B(KEYINPUT13), .Z(new_n602_));
  INV_X1    g401(.A(new_n599_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n602_), .B1(new_n603_), .B2(new_n597_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n601_), .A2(new_n604_), .ZN(new_n605_));
  AND4_X1   g404(.A1(new_n425_), .A2(new_n553_), .A3(new_n578_), .A4(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n606_), .A2(new_n534_), .A3(new_n367_), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n607_), .A2(KEYINPUT102), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(KEYINPUT102), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n608_), .A2(KEYINPUT38), .A3(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n399_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n421_), .A2(new_n398_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n422_), .A2(new_n289_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n611_), .B1(new_n614_), .B2(new_n310_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n514_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n605_), .ZN(new_n618_));
  NOR3_X1   g417(.A1(new_n618_), .A2(new_n577_), .A3(new_n549_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT103), .ZN(new_n621_));
  OAI21_X1  g420(.A(G1gat), .B1(new_n621_), .B2(new_n366_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n610_), .A2(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(KEYINPUT38), .B1(new_n608_), .B2(new_n609_), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n623_), .A2(new_n624_), .ZN(G1324gat));
  INV_X1    g424(.A(new_n289_), .ZN(new_n626_));
  AND3_X1   g425(.A1(new_n606_), .A2(new_n626_), .A3(new_n533_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT104), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n617_), .A2(new_n626_), .A3(new_n619_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n629_), .A2(G8gat), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT39), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n630_), .A2(KEYINPUT39), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n628_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT40), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n628_), .A2(new_n632_), .A3(KEYINPUT40), .A4(new_n631_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(G1325gat));
  INV_X1    g436(.A(G15gat), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT103), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n620_), .B(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n638_), .B1(new_n640_), .B2(new_n424_), .ZN(new_n641_));
  XOR2_X1   g440(.A(KEYINPUT105), .B(KEYINPUT41), .Z(new_n642_));
  OR2_X1    g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n606_), .A2(new_n638_), .A3(new_n424_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n641_), .A2(new_n642_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n643_), .A2(new_n644_), .A3(new_n645_), .ZN(G1326gat));
  INV_X1    g445(.A(G22gat), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n606_), .A2(new_n647_), .A3(new_n397_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT42), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n640_), .A2(new_n397_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n649_), .B1(new_n650_), .B2(G22gat), .ZN(new_n651_));
  AOI211_X1 g450(.A(KEYINPUT42), .B(new_n647_), .C1(new_n640_), .C2(new_n397_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n648_), .B1(new_n651_), .B2(new_n652_), .ZN(G1327gat));
  NAND2_X1  g452(.A1(new_n616_), .A2(new_n549_), .ZN(new_n654_));
  NOR4_X1   g453(.A1(new_n615_), .A2(new_n577_), .A3(new_n618_), .A4(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(G29gat), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n655_), .A2(new_n656_), .A3(new_n367_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n605_), .A2(new_n578_), .A3(new_n549_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n515_), .B(KEYINPUT106), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  OAI21_X1  g459(.A(KEYINPUT43), .B1(new_n615_), .B2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT43), .ZN(new_n662_));
  INV_X1    g461(.A(new_n515_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n425_), .A2(new_n662_), .A3(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n658_), .B1(new_n661_), .B2(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n366_), .B1(new_n665_), .B2(KEYINPUT44), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT107), .ZN(new_n667_));
  NOR3_X1   g466(.A1(new_n665_), .A2(new_n667_), .A3(KEYINPUT44), .ZN(new_n668_));
  INV_X1    g467(.A(new_n658_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n662_), .B1(new_n425_), .B2(new_n659_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n663_), .A2(new_n662_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n615_), .A2(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n669_), .B1(new_n670_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT44), .ZN(new_n674_));
  AOI21_X1  g473(.A(KEYINPUT107), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n666_), .B1(new_n668_), .B2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT108), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n676_), .A2(new_n677_), .A3(G29gat), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n677_), .B1(new_n676_), .B2(G29gat), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n657_), .B1(new_n678_), .B2(new_n679_), .ZN(G1328gat));
  INV_X1    g479(.A(G36gat), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n655_), .A2(new_n681_), .A3(new_n626_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT45), .ZN(new_n683_));
  OAI211_X1 g482(.A(KEYINPUT44), .B(new_n669_), .C1(new_n670_), .C2(new_n672_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(new_n626_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n667_), .B1(new_n665_), .B2(KEYINPUT44), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n673_), .A2(KEYINPUT107), .A3(new_n674_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n685_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n683_), .B1(new_n688_), .B2(new_n681_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT46), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  OAI211_X1 g490(.A(new_n683_), .B(KEYINPUT46), .C1(new_n688_), .C2(new_n681_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(G1329gat));
  AND2_X1   g492(.A1(new_n424_), .A2(G43gat), .ZN(new_n694_));
  OAI211_X1 g493(.A(new_n684_), .B(new_n694_), .C1(new_n668_), .C2(new_n675_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n655_), .A2(new_n424_), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n696_), .A2(G43gat), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT47), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT47), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n695_), .A2(new_n700_), .A3(new_n697_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(G1330gat));
  AOI21_X1  g501(.A(G50gat), .B1(new_n655_), .B2(new_n397_), .ZN(new_n703_));
  AOI22_X1  g502(.A1(new_n686_), .A2(new_n687_), .B1(KEYINPUT44), .B2(new_n665_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n397_), .A2(G50gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n703_), .B1(new_n704_), .B2(new_n705_), .ZN(G1331gat));
  AND2_X1   g505(.A1(new_n553_), .A2(new_n618_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n707_), .A2(KEYINPUT109), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n707_), .A2(KEYINPUT109), .ZN(new_n709_));
  NOR4_X1   g508(.A1(new_n708_), .A2(new_n709_), .A3(new_n615_), .A4(new_n578_), .ZN(new_n710_));
  INV_X1    g509(.A(G57gat), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n710_), .A2(new_n711_), .A3(new_n367_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n550_), .A2(new_n577_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n605_), .A2(new_n713_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n617_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  OAI21_X1  g515(.A(G57gat), .B1(new_n716_), .B2(new_n366_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n712_), .A2(new_n717_), .ZN(G1332gat));
  INV_X1    g517(.A(G64gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n719_), .B1(new_n715_), .B2(new_n626_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(KEYINPUT110), .B(KEYINPUT48), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n720_), .B(new_n721_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n710_), .A2(new_n719_), .A3(new_n626_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(G1333gat));
  INV_X1    g523(.A(G71gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n725_), .B1(new_n715_), .B2(new_n424_), .ZN(new_n726_));
  XOR2_X1   g525(.A(new_n726_), .B(KEYINPUT49), .Z(new_n727_));
  NAND3_X1  g526(.A1(new_n710_), .A2(new_n725_), .A3(new_n424_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1334gat));
  INV_X1    g528(.A(G78gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n730_), .B1(new_n715_), .B2(new_n397_), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT50), .Z(new_n732_));
  NAND3_X1  g531(.A1(new_n710_), .A2(new_n730_), .A3(new_n397_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1335gat));
  NOR4_X1   g533(.A1(new_n615_), .A2(new_n578_), .A3(new_n605_), .A4(new_n654_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n735_), .A2(new_n464_), .A3(new_n367_), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n605_), .A2(new_n578_), .A3(new_n550_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n737_), .B1(new_n670_), .B2(new_n672_), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n738_), .A2(new_n366_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n736_), .B1(new_n740_), .B2(new_n464_), .ZN(G1336gat));
  OAI21_X1  g540(.A(G92gat), .B1(new_n738_), .B2(new_n289_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n735_), .A2(new_n465_), .A3(new_n626_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  XOR2_X1   g543(.A(new_n744_), .B(KEYINPUT111), .Z(G1337gat));
  OAI211_X1 g544(.A(new_n735_), .B(new_n424_), .C1(new_n460_), .C2(new_n461_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT112), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n746_), .B(new_n747_), .ZN(new_n748_));
  OAI21_X1  g547(.A(G99gat), .B1(new_n738_), .B2(new_n310_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT51), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT51), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n748_), .A2(new_n752_), .A3(new_n749_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n751_), .A2(new_n753_), .ZN(G1338gat));
  XNOR2_X1  g553(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n397_), .B(new_n737_), .C1(new_n670_), .C2(new_n672_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(G106gat), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT52), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n735_), .A2(new_n432_), .A3(new_n397_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n755_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n757_), .A2(KEYINPUT52), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT52), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n762_), .B1(new_n756_), .B2(G106gat), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n759_), .B(new_n755_), .C1(new_n761_), .C2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n760_), .A2(new_n765_), .ZN(G1339gat));
  AOI22_X1  g565(.A1(new_n573_), .A2(new_n575_), .B1(new_n591_), .B2(new_n596_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT55), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n584_), .A2(new_n587_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n768_), .B1(new_n582_), .B2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT12), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n589_), .A2(new_n771_), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n588_), .A2(new_n772_), .A3(KEYINPUT55), .A4(new_n580_), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n584_), .B(new_n580_), .C1(new_n581_), .C2(KEYINPUT12), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n586_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n770_), .A2(new_n773_), .A3(new_n775_), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n776_), .A2(KEYINPUT56), .A3(new_n595_), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT56), .B1(new_n776_), .B2(new_n595_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n767_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n560_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n559_), .A2(new_n566_), .A3(new_n562_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n780_), .A2(new_n558_), .A3(new_n781_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n575_), .A2(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n783_), .B1(new_n603_), .B2(new_n597_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n779_), .A2(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(KEYINPUT57), .B1(new_n785_), .B2(new_n514_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n599_), .A2(new_n783_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n776_), .A2(KEYINPUT56), .A3(new_n595_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n788_), .B1(new_n778_), .B2(KEYINPUT114), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT114), .ZN(new_n790_));
  AOI211_X1 g589(.A(new_n790_), .B(KEYINPUT56), .C1(new_n776_), .C2(new_n595_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n787_), .B1(new_n789_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT58), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n515_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  OAI211_X1 g593(.A(KEYINPUT58), .B(new_n787_), .C1(new_n789_), .C2(new_n791_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n786_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n785_), .A2(KEYINPUT57), .A3(new_n514_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n550_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT54), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n618_), .A2(new_n713_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n799_), .B1(new_n800_), .B2(new_n515_), .ZN(new_n801_));
  NOR4_X1   g600(.A1(new_n618_), .A2(new_n663_), .A3(KEYINPUT54), .A4(new_n713_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n798_), .A2(new_n803_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n626_), .A2(new_n397_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n805_), .A2(new_n367_), .A3(new_n424_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n804_), .A2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(G113gat), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n807_), .A2(new_n808_), .A3(new_n578_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT59), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n807_), .A2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n797_), .B1(new_n796_), .B2(KEYINPUT115), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT115), .ZN(new_n813_));
  AOI211_X1 g612(.A(new_n813_), .B(new_n786_), .C1(new_n795_), .C2(new_n794_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n549_), .B1(new_n812_), .B2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT116), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n803_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  OAI211_X1 g616(.A(KEYINPUT116), .B(new_n549_), .C1(new_n812_), .C2(new_n814_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n806_), .A2(KEYINPUT59), .ZN(new_n820_));
  AOI211_X1 g619(.A(new_n577_), .B(new_n811_), .C1(new_n819_), .C2(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n809_), .B1(new_n821_), .B2(new_n808_), .ZN(G1340gat));
  INV_X1    g621(.A(G120gat), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(new_n605_), .B2(KEYINPUT60), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n807_), .B(new_n824_), .C1(KEYINPUT60), .C2(new_n823_), .ZN(new_n825_));
  AOI211_X1 g624(.A(new_n605_), .B(new_n811_), .C1(new_n819_), .C2(new_n820_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n825_), .B1(new_n826_), .B2(new_n823_), .ZN(G1341gat));
  AOI21_X1  g626(.A(G127gat), .B1(new_n807_), .B2(new_n550_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n811_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n550_), .A2(G127gat), .ZN(new_n830_));
  XOR2_X1   g629(.A(new_n830_), .B(KEYINPUT117), .Z(new_n831_));
  AOI21_X1  g630(.A(new_n828_), .B1(new_n829_), .B2(new_n831_), .ZN(G1342gat));
  AOI21_X1  g631(.A(G134gat), .B1(new_n807_), .B2(new_n616_), .ZN(new_n833_));
  XOR2_X1   g632(.A(KEYINPUT118), .B(G134gat), .Z(new_n834_));
  NOR2_X1   g633(.A1(new_n515_), .A2(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n833_), .B1(new_n829_), .B2(new_n835_), .ZN(G1343gat));
  NAND4_X1  g635(.A1(new_n289_), .A2(new_n367_), .A3(new_n397_), .A4(new_n310_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(KEYINPUT119), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n804_), .A2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n578_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g640(.A1(new_n839_), .A2(new_n618_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g642(.A1(new_n839_), .A2(new_n550_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(KEYINPUT61), .B(G155gat), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n844_), .B(new_n845_), .ZN(G1346gat));
  NAND3_X1  g645(.A1(new_n839_), .A2(G162gat), .A3(new_n659_), .ZN(new_n847_));
  NOR3_X1   g646(.A1(new_n804_), .A2(new_n514_), .A3(new_n838_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n847_), .B1(new_n848_), .B2(G162gat), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(KEYINPUT120), .ZN(G1347gat));
  INV_X1    g649(.A(KEYINPUT121), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n851_), .A2(KEYINPUT62), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n626_), .A2(new_n368_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n398_), .ZN(new_n855_));
  AOI211_X1 g654(.A(new_n577_), .B(new_n855_), .C1(new_n817_), .C2(new_n818_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n222_), .B1(new_n851_), .B2(KEYINPUT62), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n852_), .B1(new_n856_), .B2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n852_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n855_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n819_), .A2(new_n861_), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n857_), .B(new_n860_), .C1(new_n862_), .C2(new_n577_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n856_), .A2(new_n219_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n859_), .A2(new_n863_), .A3(new_n864_), .ZN(G1348gat));
  NOR2_X1   g664(.A1(new_n804_), .A2(new_n397_), .ZN(new_n866_));
  AND4_X1   g665(.A1(G176gat), .A2(new_n866_), .A3(new_n618_), .A4(new_n854_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT122), .ZN(new_n868_));
  AOI211_X1 g667(.A(new_n605_), .B(new_n855_), .C1(new_n817_), .C2(new_n818_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n868_), .B1(new_n869_), .B2(G176gat), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n819_), .A2(new_n618_), .A3(new_n861_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n871_), .A2(KEYINPUT122), .A3(new_n221_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n867_), .B1(new_n870_), .B2(new_n872_), .ZN(G1349gat));
  NOR2_X1   g672(.A1(new_n549_), .A2(new_n234_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(KEYINPUT123), .B1(new_n862_), .B2(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n855_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT123), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n877_), .A2(new_n878_), .A3(new_n874_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n866_), .A2(new_n550_), .A3(new_n854_), .ZN(new_n880_));
  INV_X1    g679(.A(G183gat), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  AND3_X1   g681(.A1(new_n876_), .A2(new_n879_), .A3(new_n882_), .ZN(G1350gat));
  OAI21_X1  g682(.A(G190gat), .B1(new_n862_), .B2(new_n515_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n877_), .A2(new_n230_), .A3(new_n616_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(G1351gat));
  NAND3_X1  g685(.A1(new_n626_), .A2(new_n422_), .A3(new_n310_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n804_), .A2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(new_n578_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g689(.A1(new_n888_), .A2(new_n618_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT124), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n892_), .B2(G204gat), .ZN(new_n893_));
  XNOR2_X1  g692(.A(KEYINPUT124), .B(G204gat), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n891_), .B2(new_n894_), .ZN(G1353gat));
  NAND2_X1  g694(.A1(new_n888_), .A2(new_n550_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT63), .ZN(new_n897_));
  INV_X1    g696(.A(G211gat), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n896_), .A2(new_n897_), .A3(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT126), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  NAND4_X1  g700(.A1(new_n896_), .A2(KEYINPUT126), .A3(new_n897_), .A4(new_n898_), .ZN(new_n902_));
  XOR2_X1   g701(.A(KEYINPUT63), .B(G211gat), .Z(new_n903_));
  INV_X1    g702(.A(new_n903_), .ZN(new_n904_));
  OR3_X1    g703(.A1(new_n896_), .A2(KEYINPUT125), .A3(new_n904_), .ZN(new_n905_));
  OAI21_X1  g704(.A(KEYINPUT125), .B1(new_n896_), .B2(new_n904_), .ZN(new_n906_));
  AOI22_X1  g705(.A1(new_n901_), .A2(new_n902_), .B1(new_n905_), .B2(new_n906_), .ZN(G1354gat));
  INV_X1    g706(.A(G218gat), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n888_), .A2(new_n908_), .A3(new_n616_), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n804_), .A2(new_n515_), .A3(new_n887_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n909_), .B1(new_n910_), .B2(new_n908_), .ZN(new_n911_));
  XOR2_X1   g710(.A(new_n911_), .B(KEYINPUT127), .Z(G1355gat));
endmodule


