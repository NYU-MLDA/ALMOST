//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 0 1 0 1 1 1 0 1 0 1 1 1 1 0 0 0 1 0 0 0 1 1 0 0 1 0 1 1 1 1 0 1 1 1 1 1 1 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n834_, new_n835_, new_n836_, new_n837_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n923_, new_n924_, new_n925_, new_n927_, new_n928_,
    new_n929_, new_n931_, new_n932_, new_n933_, new_n935_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n946_, new_n947_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n958_,
    new_n960_, new_n962_, new_n963_, new_n964_, new_n965_, new_n966_,
    new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n978_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n987_, new_n988_,
    new_n989_, new_n990_, new_n991_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT87), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  AND2_X1   g006(.A1(KEYINPUT84), .A2(KEYINPUT23), .ZN(new_n208_));
  NOR2_X1   g007(.A1(KEYINPUT84), .A2(KEYINPUT23), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n207_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n206_), .A2(new_n211_), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n210_), .B(new_n212_), .C1(G183gat), .C2(G190gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT85), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  NOR3_X1   g014(.A1(KEYINPUT85), .A2(KEYINPUT22), .A3(G176gat), .ZN(new_n216_));
  INV_X1    g015(.A(G169gat), .ZN(new_n217_));
  OR3_X1    g016(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n217_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n213_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT86), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n206_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n206_), .A2(KEYINPUT23), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n222_), .A2(new_n224_), .ZN(new_n225_));
  OR3_X1    g024(.A1(KEYINPUT83), .A2(G169gat), .A3(G176gat), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT83), .B1(G169gat), .B2(G176gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n226_), .A2(KEYINPUT24), .A3(new_n227_), .A4(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT24), .ZN(new_n230_));
  INV_X1    g029(.A(new_n227_), .ZN(new_n231_));
  NOR3_X1   g030(.A1(KEYINPUT83), .A2(G169gat), .A3(G176gat), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n230_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT25), .B(G183gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT26), .B(G190gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n225_), .A2(new_n229_), .A3(new_n233_), .A4(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n220_), .A2(new_n221_), .A3(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n221_), .B1(new_n220_), .B2(new_n237_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G71gat), .B(G99gat), .ZN(new_n242_));
  INV_X1    g041(.A(G43gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT30), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n241_), .B(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G227gat), .A2(G233gat), .ZN(new_n247_));
  INV_X1    g046(.A(G15gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n205_), .B1(new_n246_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT31), .ZN(new_n252_));
  OR2_X1    g051(.A1(new_n241_), .A2(new_n245_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n241_), .A2(new_n245_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n253_), .A2(new_n249_), .A3(new_n254_), .ZN(new_n255_));
  AND3_X1   g054(.A1(new_n251_), .A2(new_n252_), .A3(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n252_), .B1(new_n251_), .B2(new_n255_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n204_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n246_), .A2(new_n250_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n259_), .A2(KEYINPUT87), .A3(new_n255_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT31), .ZN(new_n261_));
  INV_X1    g060(.A(new_n204_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n251_), .A2(new_n252_), .A3(new_n255_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n261_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n258_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT103), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n220_), .A2(new_n237_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT86), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G197gat), .B(G204gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G211gat), .B(G218gat), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT21), .ZN(new_n272_));
  NOR3_X1   g071(.A1(new_n270_), .A2(new_n271_), .A3(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT93), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n271_), .ZN(new_n276_));
  XOR2_X1   g075(.A(G197gat), .B(G204gat), .Z(new_n277_));
  NAND3_X1  g076(.A1(new_n276_), .A2(KEYINPUT21), .A3(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT93), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT92), .ZN(new_n280_));
  INV_X1    g079(.A(G197gat), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n280_), .A2(new_n281_), .A3(G204gat), .ZN(new_n282_));
  OAI211_X1 g081(.A(KEYINPUT21), .B(new_n282_), .C1(new_n277_), .C2(new_n280_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n276_), .B1(new_n272_), .B2(new_n270_), .ZN(new_n284_));
  AOI22_X1  g083(.A1(new_n275_), .A2(new_n279_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n269_), .A2(new_n285_), .A3(new_n238_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n228_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT22), .B(G169gat), .ZN(new_n288_));
  INV_X1    g087(.A(G176gat), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n287_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(G183gat), .A2(G190gat), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n292_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT98), .B1(new_n291_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT98), .ZN(new_n295_));
  AND2_X1   g094(.A1(new_n222_), .A2(new_n224_), .ZN(new_n296_));
  OAI211_X1 g095(.A(new_n295_), .B(new_n290_), .C1(new_n296_), .C2(new_n292_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n294_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT97), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n229_), .A2(new_n233_), .A3(new_n236_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n210_), .A2(new_n212_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n299_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  AND3_X1   g101(.A1(new_n229_), .A2(new_n233_), .A3(new_n236_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n301_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n303_), .A2(KEYINPUT97), .A3(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n298_), .B1(new_n302_), .B2(new_n305_), .ZN(new_n306_));
  OAI211_X1 g105(.A(new_n286_), .B(KEYINPUT20), .C1(new_n306_), .C2(new_n285_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G226gat), .A2(G233gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT19), .ZN(new_n309_));
  XOR2_X1   g108(.A(new_n309_), .B(KEYINPUT96), .Z(new_n310_));
  OAI21_X1  g109(.A(new_n267_), .B1(new_n307_), .B2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n303_), .A2(new_n304_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n290_), .B1(new_n296_), .B2(new_n292_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT102), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n312_), .A2(KEYINPUT102), .A3(new_n313_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n316_), .A2(new_n285_), .A3(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n275_), .A2(new_n279_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n284_), .A2(new_n283_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n321_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n318_), .A2(KEYINPUT20), .A3(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(new_n309_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT20), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n325_), .B1(new_n241_), .B2(new_n285_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n298_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n305_), .A2(new_n302_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n285_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n310_), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n326_), .A2(new_n330_), .A3(KEYINPUT103), .A4(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n311_), .A2(new_n324_), .A3(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G8gat), .B(G36gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT18), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G64gat), .B(G92gat), .ZN(new_n336_));
  XOR2_X1   g135(.A(new_n335_), .B(new_n336_), .Z(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT32), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n333_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G1gat), .B(G29gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(G85gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT0), .B(G57gat), .ZN(new_n343_));
  XOR2_X1   g142(.A(new_n342_), .B(new_n343_), .Z(new_n344_));
  NAND2_X1  g143(.A1(G225gat), .A2(G233gat), .ZN(new_n345_));
  INV_X1    g144(.A(G141gat), .ZN(new_n346_));
  INV_X1    g145(.A(G148gat), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT3), .ZN(new_n348_));
  OAI211_X1 g147(.A(new_n346_), .B(new_n347_), .C1(new_n348_), .C2(KEYINPUT90), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(KEYINPUT90), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n348_), .A2(new_n346_), .A3(new_n347_), .A4(KEYINPUT90), .ZN(new_n352_));
  AND3_X1   g151(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n353_));
  AOI21_X1  g152(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n351_), .A2(new_n352_), .A3(new_n355_), .ZN(new_n356_));
  AND2_X1   g155(.A1(G155gat), .A2(G162gat), .ZN(new_n357_));
  NOR2_X1   g156(.A1(G155gat), .A2(G162gat), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n356_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT88), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT1), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n361_), .B1(new_n357_), .B2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G155gat), .A2(G162gat), .ZN(new_n364_));
  OAI22_X1  g163(.A1(new_n358_), .A2(KEYINPUT89), .B1(new_n364_), .B2(KEYINPUT1), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT89), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n357_), .A2(new_n366_), .A3(new_n362_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n364_), .A2(KEYINPUT88), .A3(KEYINPUT1), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n363_), .A2(new_n365_), .A3(new_n367_), .A4(new_n368_), .ZN(new_n369_));
  XOR2_X1   g168(.A(G141gat), .B(G148gat), .Z(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n360_), .A2(new_n371_), .A3(new_n204_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(KEYINPUT99), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n204_), .B1(new_n360_), .B2(new_n371_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n360_), .A2(new_n371_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT99), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n376_), .A2(new_n377_), .A3(new_n262_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(KEYINPUT4), .B1(new_n375_), .B2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n376_), .A2(new_n262_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n381_), .A2(KEYINPUT4), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n345_), .B1(new_n380_), .B2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n381_), .A2(KEYINPUT99), .A3(new_n372_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n385_), .A2(new_n345_), .A3(new_n378_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n344_), .B1(new_n384_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n345_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT4), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n390_), .B1(new_n385_), .B2(new_n378_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n389_), .B1(new_n391_), .B2(new_n382_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n344_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n392_), .A2(new_n386_), .A3(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n388_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n286_), .A2(KEYINPUT20), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n310_), .B1(new_n396_), .B2(new_n329_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n327_), .A2(new_n328_), .A3(new_n285_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n309_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n322_), .A2(new_n398_), .A3(KEYINPUT20), .A4(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n397_), .A2(new_n400_), .A3(new_n338_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n340_), .A2(new_n395_), .A3(new_n401_), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n397_), .A2(new_n337_), .A3(new_n400_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n337_), .B1(new_n397_), .B2(new_n400_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT33), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n392_), .A2(new_n386_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n406_), .B1(new_n407_), .B2(new_n344_), .ZN(new_n408_));
  AOI211_X1 g207(.A(KEYINPUT33), .B(new_n393_), .C1(new_n392_), .C2(new_n386_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n405_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT100), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n380_), .A2(new_n411_), .A3(new_n345_), .A4(new_n383_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n385_), .A2(new_n378_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n344_), .B1(new_n413_), .B2(new_n389_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n391_), .A2(new_n382_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n411_), .B1(new_n416_), .B2(new_n345_), .ZN(new_n417_));
  OAI21_X1  g216(.A(KEYINPUT101), .B1(new_n415_), .B2(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n380_), .A2(new_n345_), .A3(new_n383_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT100), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT101), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n420_), .A2(new_n421_), .A3(new_n412_), .A4(new_n414_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n418_), .A2(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n402_), .B1(new_n410_), .B2(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n285_), .B1(KEYINPUT29), .B2(new_n376_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT94), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G228gat), .A2(G233gat), .ZN(new_n427_));
  XOR2_X1   g226(.A(new_n427_), .B(KEYINPUT91), .Z(new_n428_));
  NAND3_X1  g227(.A1(new_n425_), .A2(new_n426_), .A3(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n376_), .A2(KEYINPUT29), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n430_), .A2(new_n321_), .A3(new_n428_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT94), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n429_), .A2(new_n432_), .ZN(new_n433_));
  OR2_X1    g232(.A1(new_n425_), .A2(new_n427_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G22gat), .B(G50gat), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT28), .B1(new_n376_), .B2(KEYINPUT29), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NOR3_X1   g238(.A1(new_n376_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n437_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  OR3_X1    g240(.A1(new_n376_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n442_), .A2(new_n438_), .A3(new_n436_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n441_), .A2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n435_), .A2(KEYINPUT95), .A3(new_n444_), .ZN(new_n445_));
  NOR3_X1   g244(.A1(new_n439_), .A2(new_n440_), .A3(new_n437_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n436_), .B1(new_n442_), .B2(new_n438_), .ZN(new_n447_));
  OAI21_X1  g246(.A(KEYINPUT95), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT95), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n441_), .A2(new_n449_), .A3(new_n443_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n448_), .A2(new_n450_), .A3(new_n434_), .A4(new_n433_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n445_), .A2(new_n451_), .ZN(new_n452_));
  XOR2_X1   g251(.A(G78gat), .B(G106gat), .Z(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n445_), .A2(new_n451_), .A3(new_n453_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n424_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT27), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n403_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n337_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n333_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n461_), .A2(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n460_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n395_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n266_), .B1(new_n459_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n395_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n258_), .A2(new_n264_), .A3(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n464_), .A2(new_n465_), .ZN(new_n472_));
  NOR3_X1   g271(.A1(new_n471_), .A2(new_n457_), .A3(new_n472_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n469_), .A2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G29gat), .B(G36gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT77), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G43gat), .B(G50gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT15), .ZN(new_n479_));
  XOR2_X1   g278(.A(G15gat), .B(G22gat), .Z(new_n480_));
  NAND2_X1  g279(.A1(G1gat), .A2(G8gat), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n480_), .B1(KEYINPUT14), .B2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT80), .ZN(new_n483_));
  XOR2_X1   g282(.A(G1gat), .B(G8gat), .Z(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT80), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n482_), .B(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n484_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n485_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  OR2_X1    g290(.A1(new_n479_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n477_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n476_), .B(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n491_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G229gat), .A2(G233gat), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n492_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n490_), .B(new_n478_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n496_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n497_), .A2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G113gat), .B(G141gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G169gat), .B(G197gat), .ZN(new_n503_));
  XOR2_X1   g302(.A(new_n502_), .B(new_n503_), .Z(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n501_), .A2(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n497_), .A2(new_n500_), .A3(new_n504_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n474_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT75), .ZN(new_n511_));
  XNOR2_X1  g310(.A(KEYINPUT67), .B(KEYINPUT6), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G99gat), .A2(G106gat), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n512_), .B(new_n514_), .ZN(new_n515_));
  XOR2_X1   g314(.A(G85gat), .B(G92gat), .Z(new_n516_));
  XOR2_X1   g315(.A(KEYINPUT66), .B(G92gat), .Z(new_n517_));
  INV_X1    g316(.A(G85gat), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n518_), .A2(KEYINPUT9), .ZN(new_n519_));
  AOI22_X1  g318(.A1(KEYINPUT9), .A2(new_n516_), .B1(new_n517_), .B2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT65), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT10), .B(G99gat), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(KEYINPUT64), .B(G106gat), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n521_), .B1(new_n523_), .B2(new_n525_), .ZN(new_n526_));
  NOR3_X1   g325(.A1(new_n522_), .A2(new_n524_), .A3(KEYINPUT65), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n515_), .B(new_n520_), .C1(new_n526_), .C2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT8), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n516_), .A2(new_n529_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(G99gat), .A2(G106gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT7), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n530_), .B1(new_n515_), .B2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT68), .B(KEYINPUT6), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(new_n514_), .ZN(new_n535_));
  OR2_X1    g334(.A1(KEYINPUT68), .A2(KEYINPUT6), .ZN(new_n536_));
  NAND2_X1  g335(.A1(KEYINPUT68), .A2(KEYINPUT6), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n536_), .A2(new_n513_), .A3(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n532_), .A2(new_n535_), .A3(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n529_), .B1(new_n539_), .B2(new_n516_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT72), .ZN(new_n541_));
  NOR3_X1   g340(.A1(new_n533_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n539_), .A2(new_n516_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT8), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n512_), .B(new_n513_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n532_), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n529_), .B(new_n516_), .C1(new_n545_), .C2(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(KEYINPUT72), .B1(new_n544_), .B2(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n528_), .B1(new_n542_), .B2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G57gat), .B(G64gat), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT69), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(G64gat), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(G57gat), .ZN(new_n554_));
  INV_X1    g353(.A(G57gat), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(G64gat), .ZN(new_n556_));
  AND3_X1   g355(.A1(new_n554_), .A2(new_n556_), .A3(new_n551_), .ZN(new_n557_));
  OAI21_X1  g356(.A(KEYINPUT11), .B1(new_n552_), .B2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G71gat), .B(G78gat), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n554_), .A2(new_n556_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(KEYINPUT69), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n550_), .A2(new_n551_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT11), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n562_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n558_), .A2(new_n560_), .A3(new_n565_), .ZN(new_n566_));
  OAI211_X1 g365(.A(KEYINPUT11), .B(new_n559_), .C1(new_n552_), .C2(new_n557_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT12), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n528_), .B1(new_n533_), .B2(new_n540_), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n566_), .A2(new_n567_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  AOI22_X1  g372(.A1(new_n549_), .A2(new_n570_), .B1(new_n569_), .B2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G230gat), .A2(G233gat), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n575_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT73), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  OAI211_X1 g377(.A(KEYINPUT73), .B(new_n575_), .C1(new_n571_), .C2(new_n572_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n574_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT70), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n582_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n544_), .A2(new_n547_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n584_), .A2(KEYINPUT70), .A3(new_n528_), .A4(new_n568_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n583_), .A2(new_n573_), .A3(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT71), .ZN(new_n587_));
  INV_X1    g386(.A(new_n575_), .ZN(new_n588_));
  AND3_X1   g387(.A1(new_n586_), .A2(new_n587_), .A3(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n587_), .B1(new_n586_), .B2(new_n588_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n581_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  XOR2_X1   g390(.A(G120gat), .B(G148gat), .Z(new_n592_));
  XNOR2_X1  g391(.A(G176gat), .B(G204gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(KEYINPUT74), .B(KEYINPUT5), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n591_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n596_), .ZN(new_n598_));
  OAI211_X1 g397(.A(new_n581_), .B(new_n598_), .C1(new_n589_), .C2(new_n590_), .ZN(new_n599_));
  AND3_X1   g398(.A1(new_n597_), .A2(KEYINPUT13), .A3(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(KEYINPUT13), .B1(new_n597_), .B2(new_n599_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n511_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT13), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n586_), .A2(new_n588_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(KEYINPUT71), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n586_), .A2(new_n587_), .A3(new_n588_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n598_), .B1(new_n607_), .B2(new_n581_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n599_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n603_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n597_), .A2(KEYINPUT13), .A3(new_n599_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n610_), .A2(KEYINPUT75), .A3(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n602_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(KEYINPUT78), .B1(new_n571_), .B2(new_n478_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT78), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n584_), .A2(new_n616_), .A3(new_n494_), .A4(new_n528_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n528_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n584_), .A2(new_n541_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n544_), .A2(KEYINPUT72), .A3(new_n547_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n618_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  OAI211_X1 g420(.A(new_n615_), .B(new_n617_), .C1(new_n621_), .C2(new_n479_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT35), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G190gat), .B(G218gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G134gat), .B(G162gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  AOI22_X1  g425(.A1(new_n622_), .A2(new_n623_), .B1(KEYINPUT36), .B2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(G232gat), .A2(G233gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT35), .ZN(new_n629_));
  XOR2_X1   g428(.A(KEYINPUT76), .B(KEYINPUT34), .Z(new_n630_));
  XOR2_X1   g429(.A(new_n629_), .B(new_n630_), .Z(new_n631_));
  INV_X1    g430(.A(KEYINPUT79), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n631_), .B1(new_n622_), .B2(new_n632_), .ZN(new_n633_));
  OR2_X1    g432(.A1(new_n621_), .A2(new_n479_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n615_), .A2(new_n617_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n631_), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n634_), .A2(KEYINPUT79), .A3(new_n635_), .A4(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n627_), .A2(new_n633_), .A3(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n626_), .A2(KEYINPUT36), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n639_), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n627_), .A2(new_n633_), .A3(new_n637_), .A4(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(KEYINPUT37), .B1(new_n640_), .B2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n640_), .A2(KEYINPUT37), .A3(new_n642_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(G231gat), .A2(G233gat), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n490_), .B(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(new_n568_), .ZN(new_n649_));
  XOR2_X1   g448(.A(G127gat), .B(G155gat), .Z(new_n650_));
  XNOR2_X1  g449(.A(G183gat), .B(G211gat), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n650_), .B(new_n651_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n652_), .B(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT17), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n654_), .A2(KEYINPUT81), .A3(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  OR2_X1    g456(.A1(new_n649_), .A2(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n656_), .B1(new_n655_), .B2(new_n654_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n649_), .A2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n646_), .A2(new_n661_), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n510_), .A2(new_n614_), .A3(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(G1gat), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n663_), .A2(new_n664_), .A3(new_n395_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT104), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT38), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n665_), .A2(KEYINPUT104), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n665_), .A2(KEYINPUT104), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n669_), .A2(KEYINPUT38), .A3(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n388_), .A2(KEYINPUT33), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n407_), .A2(new_n406_), .A3(new_n344_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n674_), .A2(new_n405_), .A3(new_n418_), .A4(new_n422_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n457_), .B1(new_n675_), .B2(new_n402_), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n445_), .A2(new_n451_), .A3(new_n453_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n453_), .B1(new_n445_), .B2(new_n451_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n470_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n679_), .A2(new_n472_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n265_), .B1(new_n676_), .B2(new_n680_), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n266_), .A2(new_n470_), .A3(new_n458_), .A4(new_n466_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n640_), .A2(new_n642_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n602_), .A2(new_n508_), .A3(new_n612_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT105), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n602_), .A2(new_n612_), .A3(KEYINPUT105), .A4(new_n508_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n661_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n688_), .A2(new_n689_), .A3(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(KEYINPUT106), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT106), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n688_), .A2(new_n693_), .A3(new_n689_), .A4(new_n690_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n685_), .B1(new_n692_), .B2(new_n694_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n695_), .A2(new_n395_), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n668_), .B(new_n671_), .C1(new_n664_), .C2(new_n696_), .ZN(G1324gat));
  INV_X1    g496(.A(KEYINPUT40), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n692_), .A2(new_n694_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n683_), .A2(new_n684_), .A3(new_n472_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT107), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n702_), .A2(new_n703_), .A3(G8gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n700_), .B1(new_n692_), .B2(new_n694_), .ZN(new_n705_));
  INV_X1    g504(.A(G8gat), .ZN(new_n706_));
  OAI21_X1  g505(.A(KEYINPUT107), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n704_), .A2(KEYINPUT39), .A3(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT39), .ZN(new_n709_));
  OAI211_X1 g508(.A(KEYINPUT107), .B(new_n709_), .C1(new_n705_), .C2(new_n706_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n663_), .A2(new_n706_), .A3(new_n472_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n698_), .B1(new_n708_), .B2(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n704_), .A2(KEYINPUT39), .A3(new_n707_), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n714_), .A2(KEYINPUT40), .A3(new_n710_), .A4(new_n711_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(G1325gat));
  NAND3_X1  g515(.A1(new_n663_), .A2(new_n248_), .A3(new_n266_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n685_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n699_), .A2(new_n266_), .A3(new_n718_), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n719_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(KEYINPUT41), .B1(new_n719_), .B2(G15gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n717_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT108), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  OAI211_X1 g523(.A(KEYINPUT108), .B(new_n717_), .C1(new_n720_), .C2(new_n721_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(G1326gat));
  INV_X1    g525(.A(G22gat), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n663_), .A2(new_n727_), .A3(new_n457_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT42), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n695_), .A2(new_n457_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n730_), .B2(G22gat), .ZN(new_n731_));
  AOI211_X1 g530(.A(KEYINPUT42), .B(new_n727_), .C1(new_n695_), .C2(new_n457_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n728_), .B1(new_n731_), .B2(new_n732_), .ZN(G1327gat));
  INV_X1    g532(.A(G29gat), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT43), .ZN(new_n735_));
  INV_X1    g534(.A(new_n645_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n736_), .A2(new_n643_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n737_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT109), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n735_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n646_), .B1(new_n469_), .B2(new_n473_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n741_), .A2(KEYINPUT109), .A3(KEYINPUT43), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n688_), .A2(new_n689_), .A3(new_n661_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(KEYINPUT44), .B1(new_n743_), .B2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT44), .ZN(new_n747_));
  AOI211_X1 g546(.A(new_n747_), .B(new_n744_), .C1(new_n740_), .C2(new_n742_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n746_), .A2(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n734_), .B1(new_n749_), .B2(new_n395_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n684_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(new_n661_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n613_), .A2(new_n752_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n510_), .A2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  NOR3_X1   g554(.A1(new_n755_), .A2(G29gat), .A3(new_n470_), .ZN(new_n756_));
  OAI21_X1  g555(.A(KEYINPUT110), .B1(new_n750_), .B2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT110), .ZN(new_n758_));
  INV_X1    g557(.A(new_n756_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n746_), .A2(new_n748_), .A3(new_n470_), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n758_), .B(new_n759_), .C1(new_n760_), .C2(new_n734_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n757_), .A2(new_n761_), .ZN(G1328gat));
  INV_X1    g561(.A(KEYINPUT46), .ZN(new_n763_));
  INV_X1    g562(.A(G36gat), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n764_), .B1(new_n749_), .B2(new_n472_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n754_), .A2(new_n764_), .A3(new_n472_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT45), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n766_), .B(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n763_), .B1(new_n765_), .B2(new_n768_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n766_), .B(KEYINPUT45), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n746_), .A2(new_n748_), .A3(new_n466_), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n770_), .B(KEYINPUT46), .C1(new_n771_), .C2(new_n764_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n769_), .A2(new_n772_), .ZN(G1329gat));
  INV_X1    g572(.A(new_n746_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n743_), .A2(KEYINPUT44), .A3(new_n745_), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n774_), .A2(G43gat), .A3(new_n266_), .A4(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n243_), .B1(new_n755_), .B2(new_n265_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(KEYINPUT47), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT47), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n776_), .A2(new_n780_), .A3(new_n777_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n781_), .ZN(G1330gat));
  INV_X1    g581(.A(G50gat), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n783_), .B1(new_n749_), .B2(new_n457_), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n755_), .A2(G50gat), .A3(new_n458_), .ZN(new_n785_));
  OAI21_X1  g584(.A(KEYINPUT111), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT111), .ZN(new_n787_));
  INV_X1    g586(.A(new_n785_), .ZN(new_n788_));
  NOR3_X1   g587(.A1(new_n746_), .A2(new_n748_), .A3(new_n458_), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n787_), .B(new_n788_), .C1(new_n789_), .C2(new_n783_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n786_), .A2(new_n790_), .ZN(G1331gat));
  NAND2_X1  g590(.A1(new_n662_), .A2(new_n613_), .ZN(new_n792_));
  OR2_X1    g591(.A1(new_n792_), .A2(KEYINPUT112), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n474_), .A2(new_n508_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(KEYINPUT112), .ZN(new_n795_));
  AND3_X1   g594(.A1(new_n793_), .A2(new_n794_), .A3(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n796_), .A2(new_n555_), .A3(new_n395_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n661_), .A2(new_n508_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n613_), .A2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n718_), .A2(new_n395_), .A3(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(G57gat), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n797_), .A2(new_n801_), .ZN(G1332gat));
  NAND3_X1  g601(.A1(new_n796_), .A2(new_n553_), .A3(new_n472_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n718_), .A2(new_n472_), .A3(new_n799_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(KEYINPUT113), .B(KEYINPUT48), .ZN(new_n805_));
  AND3_X1   g604(.A1(new_n804_), .A2(G64gat), .A3(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n805_), .B1(new_n804_), .B2(G64gat), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n803_), .B1(new_n806_), .B2(new_n807_), .ZN(G1333gat));
  NOR2_X1   g607(.A1(new_n265_), .A2(G71gat), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(KEYINPUT114), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n796_), .A2(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n718_), .A2(new_n266_), .A3(new_n799_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(G71gat), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n813_), .A2(KEYINPUT49), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n813_), .A2(KEYINPUT49), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n811_), .B1(new_n814_), .B2(new_n815_), .ZN(G1334gat));
  INV_X1    g615(.A(G78gat), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n796_), .A2(new_n817_), .A3(new_n457_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n718_), .A2(new_n457_), .A3(new_n799_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(G78gat), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n820_), .A2(KEYINPUT50), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n820_), .A2(KEYINPUT50), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n818_), .B1(new_n821_), .B2(new_n822_), .ZN(G1335gat));
  NOR2_X1   g622(.A1(new_n690_), .A2(new_n508_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n613_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT115), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n825_), .B(new_n826_), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n743_), .A2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n518_), .B1(new_n828_), .B2(new_n395_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n614_), .A2(new_n752_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n794_), .A2(new_n830_), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n831_), .A2(G85gat), .A3(new_n470_), .ZN(new_n832_));
  OR2_X1    g631(.A1(new_n829_), .A2(new_n832_), .ZN(G1336gat));
  NAND3_X1  g632(.A1(new_n828_), .A2(new_n517_), .A3(new_n472_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n831_), .A2(new_n466_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n834_), .B1(G92gat), .B2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT116), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n836_), .B(new_n837_), .ZN(G1337gat));
  NOR3_X1   g637(.A1(new_n831_), .A2(new_n522_), .A3(new_n265_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  AND2_X1   g639(.A1(new_n828_), .A2(new_n266_), .ZN(new_n841_));
  INV_X1    g640(.A(G99gat), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n840_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(KEYINPUT51), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT51), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n845_), .B(new_n840_), .C1(new_n841_), .C2(new_n842_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n846_), .ZN(G1338gat));
  XNOR2_X1  g646(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n738_), .A2(new_n739_), .A3(new_n735_), .ZN(new_n849_));
  AOI21_X1  g648(.A(KEYINPUT43), .B1(new_n741_), .B2(KEYINPUT109), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n457_), .B(new_n827_), .C1(new_n849_), .C2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(G106gat), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(KEYINPUT52), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n851_), .A2(new_n854_), .A3(G106gat), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n853_), .A2(new_n855_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n794_), .A2(new_n525_), .A3(new_n457_), .A4(new_n830_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n848_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  AND3_X1   g657(.A1(new_n851_), .A2(new_n854_), .A3(G106gat), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n854_), .B1(new_n851_), .B2(G106gat), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n857_), .B(new_n848_), .C1(new_n859_), .C2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n858_), .A2(new_n862_), .ZN(G1339gat));
  NAND3_X1  g662(.A1(new_n574_), .A2(new_n583_), .A3(new_n585_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n588_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT55), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n581_), .A2(new_n866_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n574_), .A2(new_n580_), .A3(KEYINPUT55), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n865_), .A2(new_n867_), .A3(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n596_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT56), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n869_), .A2(KEYINPUT56), .A3(new_n596_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n874_), .A2(new_n508_), .A3(new_n599_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n504_), .B1(new_n498_), .B2(new_n496_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n492_), .A2(new_n495_), .A3(new_n499_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n507_), .A2(new_n878_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n879_), .B1(new_n597_), .B2(new_n599_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n751_), .B1(new_n875_), .B2(new_n881_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n879_), .A2(new_n609_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n884_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n885_), .A2(KEYINPUT58), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n874_), .A2(KEYINPUT58), .A3(new_n883_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n646_), .ZN(new_n888_));
  OAI22_X1  g687(.A1(new_n882_), .A2(KEYINPUT57), .B1(new_n886_), .B2(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n508_), .A2(new_n599_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n890_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n684_), .B1(new_n891_), .B2(new_n880_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT57), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n661_), .B1(new_n889_), .B2(new_n894_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n798_), .A2(new_n611_), .A3(new_n610_), .ZN(new_n896_));
  OR3_X1    g695(.A1(new_n896_), .A2(new_n646_), .A3(KEYINPUT54), .ZN(new_n897_));
  OAI21_X1  g696(.A(KEYINPUT54), .B1(new_n896_), .B2(new_n646_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n895_), .A2(new_n899_), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n265_), .A2(new_n470_), .A3(new_n472_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n900_), .A2(new_n458_), .A3(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(G113gat), .B1(new_n903_), .B2(new_n508_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT118), .ZN(new_n905_));
  AOI21_X1  g704(.A(KEYINPUT59), .B1(new_n900_), .B2(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(new_n902_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n457_), .B1(new_n895_), .B2(new_n899_), .ZN(new_n908_));
  AOI21_X1  g707(.A(KEYINPUT118), .B1(new_n895_), .B2(new_n899_), .ZN(new_n909_));
  OAI211_X1 g708(.A(new_n908_), .B(new_n901_), .C1(new_n909_), .C2(KEYINPUT59), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n907_), .A2(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n508_), .A2(G113gat), .ZN(new_n912_));
  XOR2_X1   g711(.A(new_n912_), .B(KEYINPUT119), .Z(new_n913_));
  AOI21_X1  g712(.A(new_n904_), .B1(new_n911_), .B2(new_n913_), .ZN(G1340gat));
  NOR2_X1   g713(.A1(new_n614_), .A2(KEYINPUT60), .ZN(new_n915_));
  INV_X1    g714(.A(G120gat), .ZN(new_n916_));
  MUX2_X1   g715(.A(KEYINPUT60), .B(new_n915_), .S(new_n916_), .Z(new_n917_));
  NAND4_X1  g716(.A1(new_n900_), .A2(new_n458_), .A3(new_n901_), .A4(new_n917_), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT120), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n918_), .B(new_n919_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n614_), .B1(new_n907_), .B2(new_n910_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n920_), .B1(new_n921_), .B2(new_n916_), .ZN(G1341gat));
  INV_X1    g721(.A(G127gat), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n903_), .A2(new_n923_), .A3(new_n690_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n661_), .B1(new_n907_), .B2(new_n910_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(new_n925_), .B2(new_n923_), .ZN(G1342gat));
  AOI21_X1  g725(.A(G134gat), .B1(new_n903_), .B2(new_n751_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n646_), .A2(G134gat), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(KEYINPUT121), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n927_), .B1(new_n911_), .B2(new_n929_), .ZN(G1343gat));
  NOR4_X1   g729(.A1(new_n266_), .A2(new_n458_), .A3(new_n470_), .A4(new_n472_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n900_), .A2(new_n931_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n932_), .A2(new_n509_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(new_n346_), .ZN(G1344gat));
  NOR2_X1   g733(.A1(new_n932_), .A2(new_n614_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(new_n347_), .ZN(G1345gat));
  OAI21_X1  g735(.A(KEYINPUT122), .B1(new_n932_), .B2(new_n661_), .ZN(new_n937_));
  INV_X1    g736(.A(KEYINPUT122), .ZN(new_n938_));
  NAND4_X1  g737(.A1(new_n900_), .A2(new_n938_), .A3(new_n690_), .A4(new_n931_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n937_), .A2(new_n939_), .ZN(new_n940_));
  XNOR2_X1  g739(.A(KEYINPUT61), .B(G155gat), .ZN(new_n941_));
  INV_X1    g740(.A(new_n941_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n940_), .A2(new_n942_), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n937_), .A2(new_n939_), .A3(new_n941_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n943_), .A2(new_n944_), .ZN(G1346gat));
  OAI21_X1  g744(.A(G162gat), .B1(new_n932_), .B2(new_n737_), .ZN(new_n946_));
  OR2_X1    g745(.A1(new_n684_), .A2(G162gat), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n946_), .B1(new_n932_), .B2(new_n947_), .ZN(G1347gat));
  NOR2_X1   g747(.A1(new_n471_), .A2(new_n466_), .ZN(new_n949_));
  NAND4_X1  g748(.A1(new_n908_), .A2(new_n508_), .A3(new_n288_), .A4(new_n949_), .ZN(new_n950_));
  INV_X1    g749(.A(KEYINPUT62), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n949_), .A2(new_n508_), .ZN(new_n952_));
  XOR2_X1   g751(.A(new_n952_), .B(KEYINPUT123), .Z(new_n953_));
  NAND2_X1  g752(.A1(new_n908_), .A2(new_n953_), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n951_), .B1(new_n954_), .B2(G169gat), .ZN(new_n955_));
  AOI211_X1 g754(.A(KEYINPUT62), .B(new_n217_), .C1(new_n908_), .C2(new_n953_), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n950_), .B1(new_n955_), .B2(new_n956_), .ZN(G1348gat));
  NAND3_X1  g756(.A1(new_n908_), .A2(new_n613_), .A3(new_n949_), .ZN(new_n958_));
  XNOR2_X1  g757(.A(new_n958_), .B(G176gat), .ZN(G1349gat));
  NAND3_X1  g758(.A1(new_n908_), .A2(new_n690_), .A3(new_n949_), .ZN(new_n960_));
  MUX2_X1   g759(.A(new_n234_), .B(G183gat), .S(new_n960_), .Z(G1350gat));
  NAND2_X1  g760(.A1(new_n751_), .A2(new_n235_), .ZN(new_n962_));
  XNOR2_X1  g761(.A(new_n962_), .B(KEYINPUT124), .ZN(new_n963_));
  NAND3_X1  g762(.A1(new_n908_), .A2(new_n949_), .A3(new_n963_), .ZN(new_n964_));
  AND3_X1   g763(.A1(new_n908_), .A2(new_n646_), .A3(new_n949_), .ZN(new_n965_));
  INV_X1    g764(.A(G190gat), .ZN(new_n966_));
  OAI21_X1  g765(.A(new_n964_), .B1(new_n965_), .B2(new_n966_), .ZN(G1351gat));
  AOI21_X1  g766(.A(new_n737_), .B1(KEYINPUT58), .B2(new_n885_), .ZN(new_n968_));
  OR2_X1    g767(.A1(new_n885_), .A2(KEYINPUT58), .ZN(new_n969_));
  AOI22_X1  g768(.A1(new_n968_), .A2(new_n969_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n970_));
  INV_X1    g769(.A(new_n894_), .ZN(new_n971_));
  NAND2_X1  g770(.A1(new_n970_), .A2(new_n971_), .ZN(new_n972_));
  AOI22_X1  g771(.A1(new_n972_), .A2(new_n661_), .B1(new_n898_), .B2(new_n897_), .ZN(new_n973_));
  NAND3_X1  g772(.A1(new_n265_), .A2(new_n467_), .A3(new_n472_), .ZN(new_n974_));
  NOR2_X1   g773(.A1(new_n973_), .A2(new_n974_), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n975_), .A2(new_n508_), .ZN(new_n976_));
  XNOR2_X1  g775(.A(new_n976_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g776(.A1(new_n975_), .A2(new_n613_), .ZN(new_n978_));
  XNOR2_X1  g777(.A(new_n978_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g778(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n980_));
  XNOR2_X1  g779(.A(new_n980_), .B(KEYINPUT125), .ZN(new_n981_));
  INV_X1    g780(.A(KEYINPUT126), .ZN(new_n982_));
  AOI22_X1  g781(.A1(new_n981_), .A2(new_n982_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n983_));
  NAND3_X1  g782(.A1(new_n975_), .A2(new_n690_), .A3(new_n983_), .ZN(new_n984_));
  NOR2_X1   g783(.A1(new_n981_), .A2(new_n982_), .ZN(new_n985_));
  XNOR2_X1  g784(.A(new_n984_), .B(new_n985_), .ZN(G1354gat));
  AND3_X1   g785(.A1(new_n975_), .A2(G218gat), .A3(new_n646_), .ZN(new_n987_));
  NOR3_X1   g786(.A1(new_n973_), .A2(new_n684_), .A3(new_n974_), .ZN(new_n988_));
  INV_X1    g787(.A(KEYINPUT127), .ZN(new_n989_));
  OR2_X1    g788(.A1(new_n988_), .A2(new_n989_), .ZN(new_n990_));
  AOI21_X1  g789(.A(G218gat), .B1(new_n988_), .B2(new_n989_), .ZN(new_n991_));
  AOI21_X1  g790(.A(new_n987_), .B1(new_n990_), .B2(new_n991_), .ZN(G1355gat));
endmodule


