//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 0 1 0 0 0 1 1 0 0 0 1 0 1 1 0 0 1 1 0 1 1 0 0 0 1 0 0 0 1 1 1 1 0 0 1 1 1 1 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n776_, new_n777_, new_n778_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n862_,
    new_n863_, new_n864_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n873_, new_n874_, new_n875_, new_n876_,
    new_n877_, new_n878_, new_n879_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n920_, new_n921_, new_n922_, new_n924_,
    new_n925_, new_n926_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n933_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_;
  INV_X1    g000(.A(KEYINPUT38), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT74), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT73), .ZN(new_n204_));
  XOR2_X1   g003(.A(G120gat), .B(G148gat), .Z(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT5), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G176gat), .B(G204gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT72), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G57gat), .B(G64gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT11), .ZN(new_n211_));
  XOR2_X1   g010(.A(G71gat), .B(G78gat), .Z(new_n212_));
  OR2_X1    g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n210_), .A2(KEYINPUT11), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n211_), .A2(new_n212_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n213_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  XOR2_X1   g015(.A(KEYINPUT10), .B(G99gat), .Z(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT66), .B(G106gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT67), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT67), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n217_), .A2(new_n221_), .A3(new_n218_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  AOI21_X1  g022(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(KEYINPUT68), .ZN(new_n225_));
  NOR2_X1   g024(.A1(G85gat), .A2(G92gat), .ZN(new_n226_));
  AND2_X1   g025(.A1(G85gat), .A2(G92gat), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n226_), .B1(new_n227_), .B2(KEYINPUT9), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n225_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G99gat), .A2(G106gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(KEYINPUT6), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n223_), .A2(new_n229_), .A3(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT8), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n227_), .A2(new_n226_), .ZN(new_n234_));
  OR3_X1    g033(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n231_), .A2(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT69), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT69), .ZN(new_n239_));
  OAI211_X1 g038(.A(new_n239_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n238_), .A2(new_n240_), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n233_), .B(new_n234_), .C1(new_n236_), .C2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n238_), .A2(new_n240_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT70), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT6), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(KEYINPUT70), .A2(KEYINPUT6), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n246_), .A2(new_n230_), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n230_), .ZN(new_n249_));
  AND2_X1   g048(.A1(KEYINPUT70), .A2(KEYINPUT6), .ZN(new_n250_));
  NOR2_X1   g049(.A1(KEYINPUT70), .A2(KEYINPUT6), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n249_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n243_), .A2(new_n248_), .A3(new_n235_), .A4(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n233_), .B1(new_n253_), .B2(new_n234_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT71), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n242_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  AOI211_X1 g055(.A(KEYINPUT71), .B(new_n233_), .C1(new_n253_), .C2(new_n234_), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n216_), .B(new_n232_), .C1(new_n256_), .C2(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G230gat), .A2(G233gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n258_), .A2(new_n262_), .ZN(new_n263_));
  AND3_X1   g062(.A1(new_n223_), .A2(new_n229_), .A3(new_n231_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n234_), .A2(new_n233_), .ZN(new_n265_));
  AND2_X1   g064(.A1(new_n231_), .A2(new_n235_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n265_), .B1(new_n266_), .B2(new_n243_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n252_), .A2(new_n248_), .A3(new_n235_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n234_), .B1(new_n268_), .B2(new_n241_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(KEYINPUT8), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n267_), .B1(new_n270_), .B2(KEYINPUT71), .ZN(new_n271_));
  INV_X1    g070(.A(new_n257_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n264_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT12), .B1(new_n273_), .B2(new_n216_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n232_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT12), .ZN(new_n276_));
  INV_X1    g075(.A(new_n216_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n275_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n263_), .B1(new_n274_), .B2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n275_), .A2(new_n277_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n262_), .B1(new_n280_), .B2(new_n258_), .ZN(new_n281_));
  OAI211_X1 g080(.A(new_n204_), .B(new_n209_), .C1(new_n279_), .C2(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n261_), .B1(new_n273_), .B2(new_n216_), .ZN(new_n283_));
  AND3_X1   g082(.A1(new_n275_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n276_), .B1(new_n275_), .B2(new_n277_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n283_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n280_), .A2(new_n258_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(new_n261_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n208_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n286_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n282_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n286_), .A2(new_n288_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n204_), .B1(new_n292_), .B2(new_n209_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n203_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n209_), .B1(new_n279_), .B2(new_n281_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(KEYINPUT73), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n296_), .A2(KEYINPUT74), .A3(new_n290_), .A4(new_n282_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n294_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT75), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT13), .ZN(new_n300_));
  OR2_X1    g099(.A1(new_n299_), .A2(KEYINPUT13), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n298_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n294_), .A2(new_n297_), .A3(new_n299_), .A4(KEYINPUT13), .ZN(new_n303_));
  AND2_X1   g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G231gat), .A2(G233gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n216_), .B(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G1gat), .B(G8gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT80), .ZN(new_n309_));
  INV_X1    g108(.A(G15gat), .ZN(new_n310_));
  INV_X1    g109(.A(G22gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G15gat), .A2(G22gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G1gat), .A2(G8gat), .ZN(new_n314_));
  AOI22_X1  g113(.A1(new_n312_), .A2(new_n313_), .B1(KEYINPUT14), .B2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n309_), .B(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n307_), .B(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G127gat), .B(G155gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G183gat), .B(G211gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  XOR2_X1   g121(.A(new_n322_), .B(KEYINPUT17), .Z(new_n323_));
  AND2_X1   g122(.A1(new_n317_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT82), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n322_), .A2(KEYINPUT17), .ZN(new_n327_));
  OR2_X1    g126(.A1(new_n317_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n324_), .A2(new_n325_), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT83), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n330_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT83), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n332_), .A2(new_n333_), .A3(new_n328_), .A4(new_n326_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n331_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G232gat), .A2(G233gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT34), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT35), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G29gat), .B(G36gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT76), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G43gat), .B(G50gat), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n342_), .A2(new_n344_), .ZN(new_n345_));
  OR2_X1    g144(.A1(new_n341_), .A2(KEYINPUT76), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n341_), .A2(KEYINPUT76), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n346_), .A2(new_n347_), .A3(new_n343_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n345_), .A2(new_n348_), .ZN(new_n349_));
  OAI22_X1  g148(.A1(new_n275_), .A2(new_n349_), .B1(KEYINPUT35), .B2(new_n337_), .ZN(new_n350_));
  AND3_X1   g149(.A1(new_n345_), .A2(KEYINPUT15), .A3(new_n348_), .ZN(new_n351_));
  AOI21_X1  g150(.A(KEYINPUT15), .B1(new_n345_), .B2(new_n348_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n273_), .A2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n340_), .B1(new_n350_), .B2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n349_), .ZN(new_n356_));
  AOI22_X1  g155(.A1(new_n273_), .A2(new_n356_), .B1(new_n339_), .B2(new_n338_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n340_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n353_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(new_n275_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n357_), .A2(new_n358_), .A3(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n355_), .A2(new_n361_), .ZN(new_n362_));
  XOR2_X1   g161(.A(G190gat), .B(G218gat), .Z(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT77), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G134gat), .B(G162gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT36), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n362_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT79), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT36), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n366_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n355_), .A2(new_n361_), .A3(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT78), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT78), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n355_), .A2(new_n361_), .A3(new_n375_), .A4(new_n372_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT79), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n362_), .A2(new_n377_), .A3(new_n367_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n369_), .A2(new_n374_), .A3(new_n376_), .A4(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT37), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n368_), .A2(new_n373_), .ZN(new_n381_));
  OR2_X1    g180(.A1(new_n381_), .A2(KEYINPUT37), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n335_), .B1(new_n380_), .B2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  OR3_X1    g183(.A1(new_n305_), .A2(KEYINPUT84), .A3(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n359_), .A2(new_n316_), .ZN(new_n386_));
  OR2_X1    g185(.A1(new_n316_), .A2(new_n349_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G229gat), .A2(G233gat), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n386_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n316_), .B(new_n349_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n388_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n389_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G113gat), .B(G141gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G169gat), .B(G197gat), .ZN(new_n396_));
  XOR2_X1   g195(.A(new_n395_), .B(new_n396_), .Z(new_n397_));
  AOI21_X1  g196(.A(KEYINPUT85), .B1(new_n394_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT85), .ZN(new_n399_));
  INV_X1    g198(.A(new_n397_), .ZN(new_n400_));
  NOR3_X1   g199(.A1(new_n393_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n401_));
  OAI22_X1  g200(.A1(new_n398_), .A2(new_n401_), .B1(new_n394_), .B2(new_n397_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G8gat), .B(G36gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(KEYINPUT18), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G64gat), .B(G92gat), .ZN(new_n406_));
  XOR2_X1   g205(.A(new_n405_), .B(new_n406_), .Z(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  XOR2_X1   g207(.A(KEYINPUT95), .B(G204gat), .Z(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(G197gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT96), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT21), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT94), .B(G197gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(G204gat), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT96), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n409_), .A2(new_n415_), .A3(G197gat), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n411_), .A2(new_n412_), .A3(new_n414_), .A4(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G211gat), .B(G218gat), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  OAI22_X1  g218(.A1(new_n409_), .A2(G197gat), .B1(new_n413_), .B2(G204gat), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n419_), .B1(new_n420_), .B2(KEYINPUT21), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n417_), .A2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n411_), .A2(new_n414_), .A3(new_n416_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n418_), .A2(new_n412_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n422_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT91), .ZN(new_n428_));
  XOR2_X1   g227(.A(KEYINPUT90), .B(G176gat), .Z(new_n429_));
  INV_X1    g228(.A(G169gat), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT22), .B1(new_n430_), .B2(KEYINPUT89), .ZN(new_n431_));
  OR2_X1    g230(.A1(new_n430_), .A2(KEYINPUT22), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n429_), .B(new_n431_), .C1(KEYINPUT89), .C2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(G176gat), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n430_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT23), .ZN(new_n437_));
  INV_X1    g236(.A(G183gat), .ZN(new_n438_));
  INV_X1    g237(.A(G190gat), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n437_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n440_), .B(new_n441_), .C1(G183gat), .C2(G190gat), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n433_), .A2(new_n436_), .A3(new_n442_), .ZN(new_n443_));
  AND2_X1   g242(.A1(new_n440_), .A2(new_n441_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(G169gat), .A2(G176gat), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT24), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n444_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT88), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n444_), .A2(KEYINPUT88), .A3(new_n447_), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NOR3_X1   g251(.A1(new_n435_), .A2(new_n446_), .A3(new_n445_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT25), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n455_), .A2(G183gat), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT86), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT26), .ZN(new_n459_));
  AOI22_X1  g258(.A1(new_n455_), .A2(G183gat), .B1(new_n459_), .B2(G190gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n458_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT87), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n462_), .B1(new_n459_), .B2(G190gat), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n439_), .A2(KEYINPUT87), .A3(KEYINPUT26), .ZN(new_n464_));
  OAI211_X1 g263(.A(new_n463_), .B(new_n464_), .C1(new_n456_), .C2(new_n457_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n454_), .B1(new_n461_), .B2(new_n465_), .ZN(new_n466_));
  OAI211_X1 g265(.A(new_n428_), .B(new_n443_), .C1(new_n452_), .C2(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n466_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n443_), .ZN(new_n469_));
  OAI21_X1  g268(.A(KEYINPUT91), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n427_), .B1(new_n467_), .B2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G226gat), .A2(G233gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n472_), .B(KEYINPUT19), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT22), .B(G169gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n429_), .A2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n476_), .A2(new_n442_), .A3(new_n436_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT100), .ZN(new_n478_));
  XNOR2_X1  g277(.A(KEYINPUT25), .B(G183gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(KEYINPUT26), .B(G190gat), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n453_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT98), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n482_), .B1(new_n444_), .B2(new_n447_), .ZN(new_n483_));
  AND4_X1   g282(.A1(new_n482_), .A2(new_n440_), .A3(new_n447_), .A4(new_n441_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n481_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT99), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  OAI211_X1 g286(.A(new_n481_), .B(KEYINPUT99), .C1(new_n483_), .C2(new_n484_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n478_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n474_), .B1(new_n489_), .B2(new_n426_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT20), .ZN(new_n491_));
  NOR3_X1   g290(.A1(new_n471_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n491_), .B1(new_n489_), .B2(new_n426_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n427_), .A2(new_n467_), .A3(new_n470_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n474_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n408_), .B1(new_n492_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n495_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n467_), .A2(new_n470_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(new_n426_), .ZN(new_n499_));
  OR2_X1    g298(.A1(new_n489_), .A2(new_n426_), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n499_), .A2(new_n500_), .A3(KEYINPUT20), .A4(new_n474_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n497_), .A2(new_n501_), .A3(new_n407_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n496_), .A2(new_n502_), .A3(KEYINPUT101), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT27), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT101), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n505_), .B(new_n408_), .C1(new_n492_), .C2(new_n495_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n503_), .A2(new_n504_), .A3(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT29), .ZN(new_n508_));
  NOR2_X1   g307(.A1(KEYINPUT93), .A2(KEYINPUT3), .ZN(new_n509_));
  INV_X1    g308(.A(G141gat), .ZN(new_n510_));
  INV_X1    g309(.A(G148gat), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n509_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G141gat), .A2(G148gat), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT2), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  OAI22_X1  g314(.A1(KEYINPUT93), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n516_));
  NAND3_X1  g315(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n512_), .A2(new_n515_), .A3(new_n516_), .A4(new_n517_), .ZN(new_n518_));
  OR2_X1    g317(.A1(G155gat), .A2(G162gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G155gat), .A2(G162gat), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n518_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n510_), .A2(new_n511_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(KEYINPUT1), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(new_n519_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n520_), .A2(KEYINPUT1), .ZN(new_n525_));
  OAI211_X1 g324(.A(new_n522_), .B(new_n513_), .C1(new_n524_), .C2(new_n525_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n521_), .A2(new_n526_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n426_), .B1(new_n508_), .B2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G228gat), .A2(G233gat), .ZN(new_n529_));
  XOR2_X1   g328(.A(new_n528_), .B(new_n529_), .Z(new_n530_));
  NAND2_X1  g329(.A1(new_n521_), .A2(new_n526_), .ZN(new_n531_));
  OR3_X1    g330(.A1(new_n531_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n532_));
  OAI21_X1  g331(.A(KEYINPUT28), .B1(new_n531_), .B2(KEYINPUT29), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G22gat), .B(G50gat), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  AND3_X1   g334(.A1(new_n532_), .A2(new_n533_), .A3(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n535_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G78gat), .B(G106gat), .ZN(new_n538_));
  OR3_X1    g337(.A1(new_n536_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT97), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n540_), .B(new_n538_), .C1(new_n536_), .C2(new_n537_), .ZN(new_n541_));
  AND3_X1   g340(.A1(new_n530_), .A2(new_n539_), .A3(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n530_), .B1(new_n539_), .B2(new_n541_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n471_), .A2(new_n491_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n427_), .A2(new_n485_), .A3(new_n477_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n474_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  AND3_X1   g346(.A1(new_n493_), .A2(new_n474_), .A3(new_n494_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n408_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n549_), .A2(KEYINPUT27), .A3(new_n502_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n507_), .A2(new_n544_), .A3(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT105), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n507_), .A2(KEYINPUT105), .A3(new_n544_), .A4(new_n550_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G227gat), .A2(G233gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(new_n310_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT30), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT31), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G71gat), .B(G99gat), .ZN(new_n560_));
  INV_X1    g359(.A(G43gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n498_), .B(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(G127gat), .B(G134gat), .Z(new_n565_));
  XOR2_X1   g364(.A(G113gat), .B(G120gat), .Z(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT92), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G127gat), .B(G134gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G113gat), .B(G120gat), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n567_), .A2(new_n568_), .A3(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n569_), .A2(new_n570_), .A3(KEYINPUT92), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n564_), .A2(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n563_), .A2(new_n573_), .A3(new_n572_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n559_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n575_), .A2(new_n559_), .A3(new_n576_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  XOR2_X1   g379(.A(G1gat), .B(G29gat), .Z(new_n581_));
  XNOR2_X1  g380(.A(G57gat), .B(G85gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(KEYINPUT103), .B(KEYINPUT0), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n574_), .A2(new_n531_), .ZN(new_n586_));
  OAI211_X1 g385(.A(G225gat), .B(G233gat), .C1(new_n586_), .C2(KEYINPUT4), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n567_), .A2(new_n571_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n527_), .A2(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n590_), .A2(KEYINPUT4), .A3(new_n586_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n588_), .A2(KEYINPUT102), .A3(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G225gat), .A2(G233gat), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n590_), .A2(new_n586_), .A3(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT102), .ZN(new_n596_));
  INV_X1    g395(.A(new_n591_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n596_), .B1(new_n597_), .B2(new_n587_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n585_), .B1(new_n595_), .B2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n585_), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n598_), .A2(new_n592_), .A3(new_n601_), .A4(new_n594_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n580_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n555_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT104), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n407_), .A2(KEYINPUT32), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n497_), .A2(new_n501_), .A3(new_n608_), .A4(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n609_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n611_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n497_), .A2(new_n501_), .A3(new_n609_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(KEYINPUT104), .ZN(new_n614_));
  AND4_X1   g413(.A1(new_n610_), .A2(new_n612_), .A3(new_n614_), .A4(new_n603_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n592_), .A2(new_n594_), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n616_), .A2(KEYINPUT33), .A3(new_n601_), .A4(new_n598_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT33), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n602_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n590_), .A2(new_n586_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n593_), .B1(new_n586_), .B2(KEYINPUT4), .ZN(new_n621_));
  OAI221_X1 g420(.A(new_n585_), .B1(new_n620_), .B2(new_n593_), .C1(new_n597_), .C2(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n617_), .A2(new_n619_), .A3(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n623_), .B1(new_n503_), .B2(new_n506_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n544_), .B1(new_n615_), .B2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n544_), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n626_), .A2(new_n507_), .A3(new_n604_), .A4(new_n550_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n625_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n580_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n403_), .B1(new_n607_), .B2(new_n630_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n385_), .A2(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(KEYINPUT84), .B1(new_n305_), .B2(new_n384_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n604_), .A2(G1gat), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n632_), .A2(new_n633_), .A3(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(KEYINPUT106), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n635_), .A2(KEYINPUT106), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n202_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n635_), .A2(KEYINPUT106), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n640_), .A2(KEYINPUT38), .A3(new_n636_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT107), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n381_), .B(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n643_), .B1(new_n607_), .B2(new_n630_), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n304_), .A2(new_n402_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n329_), .A2(new_n330_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n644_), .A2(new_n645_), .A3(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(G1gat), .B1(new_n647_), .B2(new_n604_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n639_), .A2(new_n641_), .A3(new_n648_), .ZN(G1324gat));
  NAND2_X1  g448(.A1(new_n507_), .A2(new_n550_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(G8gat), .B1(new_n647_), .B2(new_n651_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT39), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n651_), .A2(G8gat), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n385_), .A2(new_n631_), .A3(new_n633_), .A4(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT108), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n653_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT40), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n653_), .A2(new_n656_), .A3(KEYINPUT40), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(G1325gat));
  OAI21_X1  g460(.A(G15gat), .B1(new_n647_), .B2(new_n629_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT41), .Z(new_n663_));
  AND2_X1   g462(.A1(new_n632_), .A2(new_n633_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n664_), .A2(new_n310_), .A3(new_n580_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n663_), .A2(new_n665_), .ZN(G1326gat));
  NAND3_X1  g465(.A1(new_n664_), .A2(new_n311_), .A3(new_n626_), .ZN(new_n667_));
  OAI21_X1  g466(.A(G22gat), .B1(new_n647_), .B2(new_n544_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT42), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(G1327gat));
  INV_X1    g469(.A(new_n643_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n335_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n605_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n580_), .B1(new_n625_), .B2(new_n627_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n673_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n304_), .A2(new_n402_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(G29gat), .B1(new_n678_), .B2(new_n603_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n645_), .A2(new_n335_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n380_), .A2(new_n382_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n682_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(KEYINPUT43), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT43), .ZN(new_n685_));
  OAI211_X1 g484(.A(new_n685_), .B(new_n682_), .C1(new_n674_), .C2(new_n675_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n680_), .B1(new_n684_), .B2(new_n686_), .ZN(new_n687_));
  XOR2_X1   g486(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n688_));
  NOR2_X1   g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n684_), .A2(new_n686_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n677_), .A2(new_n672_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n690_), .A2(KEYINPUT44), .A3(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n689_), .A2(new_n693_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n603_), .A2(G29gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n679_), .B1(new_n694_), .B2(new_n695_), .ZN(G1328gat));
  OAI211_X1 g495(.A(new_n692_), .B(new_n650_), .C1(new_n687_), .C2(new_n688_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(G36gat), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT112), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n699_), .A2(KEYINPUT46), .ZN(new_n700_));
  XOR2_X1   g499(.A(KEYINPUT110), .B(KEYINPUT45), .Z(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n651_), .A2(G36gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(KEYINPUT111), .B1(new_n678_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT111), .ZN(new_n705_));
  INV_X1    g504(.A(new_n703_), .ZN(new_n706_));
  NOR4_X1   g505(.A1(new_n676_), .A2(new_n677_), .A3(new_n705_), .A4(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n702_), .B1(new_n704_), .B2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n607_), .A2(new_n630_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n645_), .A2(new_n709_), .A3(new_n673_), .A4(new_n703_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(new_n705_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n678_), .A2(KEYINPUT111), .A3(new_n703_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n711_), .A2(new_n712_), .A3(new_n701_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n700_), .B1(new_n708_), .B2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n699_), .A2(KEYINPUT46), .ZN(new_n715_));
  AND3_X1   g514(.A1(new_n698_), .A2(new_n714_), .A3(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n715_), .B1(new_n698_), .B2(new_n714_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n716_), .A2(new_n717_), .ZN(G1329gat));
  NOR2_X1   g517(.A1(new_n629_), .A2(new_n561_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n694_), .A2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT47), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n678_), .A2(new_n580_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(new_n561_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n720_), .A2(new_n721_), .A3(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n719_), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n689_), .A2(new_n693_), .A3(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n723_), .ZN(new_n727_));
  OAI21_X1  g526(.A(KEYINPUT47), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n724_), .A2(new_n728_), .ZN(G1330gat));
  AOI21_X1  g528(.A(G50gat), .B1(new_n678_), .B2(new_n626_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n626_), .A2(G50gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n694_), .B2(new_n731_), .ZN(G1331gat));
  NAND2_X1  g531(.A1(new_n709_), .A2(new_n403_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n305_), .A2(new_n383_), .ZN(new_n734_));
  OR3_X1    g533(.A1(new_n733_), .A2(KEYINPUT113), .A3(new_n734_), .ZN(new_n735_));
  OAI21_X1  g534(.A(KEYINPUT113), .B1(new_n733_), .B2(new_n734_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(G57gat), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n737_), .A2(new_n738_), .A3(new_n603_), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n304_), .A2(new_n335_), .A3(new_n402_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n644_), .A2(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(G57gat), .B1(new_n741_), .B2(new_n604_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n739_), .A2(new_n742_), .ZN(G1332gat));
  INV_X1    g542(.A(G64gat), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n735_), .A2(new_n744_), .A3(new_n650_), .A4(new_n736_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT48), .ZN(new_n746_));
  INV_X1    g545(.A(new_n741_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(new_n650_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n746_), .B1(new_n748_), .B2(G64gat), .ZN(new_n749_));
  AOI211_X1 g548(.A(KEYINPUT48), .B(new_n744_), .C1(new_n747_), .C2(new_n650_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n745_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT114), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n751_), .B(new_n752_), .ZN(G1333gat));
  INV_X1    g552(.A(G71gat), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n580_), .A2(new_n754_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT116), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n737_), .A2(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n754_), .B1(new_n747_), .B2(new_n580_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(KEYINPUT115), .B(KEYINPUT49), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n758_), .A2(new_n759_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n757_), .B1(new_n760_), .B2(new_n761_), .ZN(G1334gat));
  INV_X1    g561(.A(G78gat), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n737_), .A2(new_n763_), .A3(new_n626_), .ZN(new_n764_));
  OAI21_X1  g563(.A(G78gat), .B1(new_n741_), .B2(new_n544_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT50), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(G1335gat));
  AND4_X1   g566(.A1(new_n305_), .A2(new_n709_), .A3(new_n403_), .A4(new_n673_), .ZN(new_n768_));
  AOI21_X1  g567(.A(G85gat), .B1(new_n768_), .B2(new_n603_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n305_), .A2(new_n335_), .A3(new_n403_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n770_), .B1(new_n684_), .B2(new_n686_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT117), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n603_), .A2(G85gat), .ZN(new_n773_));
  XOR2_X1   g572(.A(new_n773_), .B(KEYINPUT118), .Z(new_n774_));
  AOI21_X1  g573(.A(new_n769_), .B1(new_n772_), .B2(new_n774_), .ZN(G1336gat));
  INV_X1    g574(.A(G92gat), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n768_), .A2(new_n776_), .A3(new_n650_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n772_), .A2(new_n650_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n777_), .B1(new_n778_), .B2(new_n776_), .ZN(G1337gat));
  NAND3_X1  g578(.A1(new_n768_), .A2(new_n217_), .A3(new_n580_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT119), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n780_), .B(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT51), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n771_), .A2(new_n580_), .ZN(new_n784_));
  INV_X1    g583(.A(G99gat), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n782_), .B(new_n783_), .C1(new_n784_), .C2(new_n785_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n780_), .B(KEYINPUT119), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n784_), .A2(new_n785_), .ZN(new_n788_));
  OAI21_X1  g587(.A(KEYINPUT51), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n786_), .A2(new_n789_), .ZN(G1338gat));
  NAND3_X1  g589(.A1(new_n768_), .A2(new_n218_), .A3(new_n626_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT52), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n771_), .A2(new_n626_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n792_), .B1(new_n793_), .B2(G106gat), .ZN(new_n794_));
  INV_X1    g593(.A(G106gat), .ZN(new_n795_));
  AOI211_X1 g594(.A(KEYINPUT52), .B(new_n795_), .C1(new_n771_), .C2(new_n626_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n791_), .B1(new_n794_), .B2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT53), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT53), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n799_), .B(new_n791_), .C1(new_n794_), .C2(new_n796_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n798_), .A2(new_n800_), .ZN(G1339gat));
  NAND3_X1  g600(.A1(new_n555_), .A2(new_n580_), .A3(new_n603_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n398_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n401_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n386_), .A2(new_n387_), .A3(new_n391_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n397_), .B1(new_n390_), .B2(new_n388_), .ZN(new_n806_));
  AOI22_X1  g605(.A1(new_n803_), .A2(new_n804_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n258_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n261_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n286_), .A2(new_n810_), .ZN(new_n811_));
  OAI211_X1 g610(.A(KEYINPUT55), .B(new_n283_), .C1(new_n284_), .C2(new_n285_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n809_), .A2(new_n811_), .A3(new_n812_), .ZN(new_n813_));
  AND3_X1   g612(.A1(new_n813_), .A2(KEYINPUT56), .A3(new_n209_), .ZN(new_n814_));
  AOI21_X1  g613(.A(KEYINPUT56), .B1(new_n813_), .B2(new_n209_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n807_), .B(new_n290_), .C1(new_n814_), .C2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT58), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n290_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n813_), .A2(new_n209_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT56), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n813_), .A2(KEYINPUT56), .A3(new_n209_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n819_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n824_), .A2(KEYINPUT58), .A3(new_n807_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n818_), .A2(new_n682_), .A3(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT57), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n298_), .A2(new_n807_), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n290_), .B(new_n402_), .C1(new_n814_), .C2(new_n815_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n827_), .B1(new_n830_), .B2(new_n671_), .ZN(new_n831_));
  AOI211_X1 g630(.A(KEYINPUT57), .B(new_n643_), .C1(new_n828_), .C2(new_n829_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n826_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n646_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n304_), .A2(new_n836_), .A3(new_n383_), .A4(new_n403_), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n383_), .A2(new_n303_), .A3(new_n302_), .A4(new_n403_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT54), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n802_), .B1(new_n835_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(G113gat), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n841_), .A2(new_n842_), .A3(new_n402_), .ZN(new_n843_));
  AOI22_X1  g642(.A1(new_n833_), .A2(new_n335_), .B1(new_n839_), .B2(new_n837_), .ZN(new_n844_));
  NOR3_X1   g643(.A1(new_n844_), .A2(KEYINPUT59), .A3(new_n802_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT120), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT59), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n846_), .B1(new_n841_), .B2(new_n847_), .ZN(new_n848_));
  AOI22_X1  g647(.A1(new_n833_), .A2(new_n834_), .B1(new_n839_), .B2(new_n837_), .ZN(new_n849_));
  OAI211_X1 g648(.A(KEYINPUT120), .B(KEYINPUT59), .C1(new_n849_), .C2(new_n802_), .ZN(new_n850_));
  AOI211_X1 g649(.A(new_n403_), .B(new_n845_), .C1(new_n848_), .C2(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n843_), .B1(new_n851_), .B2(new_n842_), .ZN(G1340gat));
  INV_X1    g651(.A(G120gat), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n853_), .B1(new_n304_), .B2(KEYINPUT60), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n841_), .B(new_n854_), .C1(KEYINPUT60), .C2(new_n853_), .ZN(new_n855_));
  AOI211_X1 g654(.A(new_n304_), .B(new_n845_), .C1(new_n848_), .C2(new_n850_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n855_), .B1(new_n856_), .B2(new_n853_), .ZN(G1341gat));
  INV_X1    g656(.A(G127gat), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n841_), .A2(new_n858_), .A3(new_n672_), .ZN(new_n859_));
  AOI211_X1 g658(.A(new_n834_), .B(new_n845_), .C1(new_n848_), .C2(new_n850_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n860_), .B2(new_n858_), .ZN(G1342gat));
  INV_X1    g660(.A(G134gat), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n841_), .A2(new_n862_), .A3(new_n643_), .ZN(new_n863_));
  AOI211_X1 g662(.A(new_n681_), .B(new_n845_), .C1(new_n848_), .C2(new_n850_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n864_), .B2(new_n862_), .ZN(G1343gat));
  NAND2_X1  g664(.A1(new_n835_), .A2(new_n840_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n629_), .A2(new_n626_), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n867_), .A2(new_n604_), .A3(new_n650_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n868_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n869_), .A2(new_n403_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(KEYINPUT121), .B(G141gat), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n870_), .B(new_n871_), .ZN(G1344gat));
  OAI21_X1  g671(.A(KEYINPUT123), .B1(new_n869_), .B2(new_n304_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n868_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n849_), .A2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT123), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n875_), .A2(new_n876_), .A3(new_n305_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n873_), .A2(new_n877_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(KEYINPUT122), .B(G148gat), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n878_), .B(new_n879_), .ZN(G1345gat));
  NAND2_X1  g679(.A1(new_n875_), .A2(new_n672_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(KEYINPUT61), .B(G155gat), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n881_), .B(new_n882_), .ZN(G1346gat));
  INV_X1    g682(.A(G162gat), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n869_), .A2(new_n884_), .A3(new_n681_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n869_), .B2(new_n671_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT124), .ZN(new_n887_));
  OR2_X1    g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n887_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n885_), .B1(new_n888_), .B2(new_n889_), .ZN(G1347gat));
  NAND2_X1  g689(.A1(new_n606_), .A2(new_n650_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(new_n626_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  OAI21_X1  g692(.A(KEYINPUT125), .B1(new_n844_), .B2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT125), .ZN(new_n895_));
  AOI22_X1  g694(.A1(new_n824_), .A2(new_n402_), .B1(new_n298_), .B2(new_n807_), .ZN(new_n896_));
  OAI21_X1  g695(.A(KEYINPUT57), .B1(new_n896_), .B2(new_n643_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n830_), .A2(new_n827_), .A3(new_n671_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n672_), .B1(new_n899_), .B2(new_n826_), .ZN(new_n900_));
  AND2_X1   g699(.A1(new_n837_), .A2(new_n839_), .ZN(new_n901_));
  OAI211_X1 g700(.A(new_n895_), .B(new_n892_), .C1(new_n900_), .C2(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n894_), .A2(new_n902_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n903_), .A2(new_n475_), .A3(new_n402_), .ZN(new_n904_));
  OAI211_X1 g703(.A(new_n402_), .B(new_n892_), .C1(new_n900_), .C2(new_n901_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(G169gat), .ZN(new_n906_));
  AND2_X1   g705(.A1(new_n906_), .A2(KEYINPUT62), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n906_), .A2(KEYINPUT62), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n904_), .B1(new_n907_), .B2(new_n908_), .ZN(G1348gat));
  NOR2_X1   g708(.A1(new_n849_), .A2(new_n626_), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n304_), .A2(new_n891_), .A3(new_n434_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n304_), .B1(new_n894_), .B2(new_n902_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n429_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n912_), .B1(new_n913_), .B2(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT126), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(new_n917_));
  OAI211_X1 g716(.A(new_n912_), .B(KEYINPUT126), .C1(new_n913_), .C2(new_n914_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(G1349gat));
  NOR2_X1   g718(.A1(new_n891_), .A2(new_n335_), .ZN(new_n920_));
  AOI21_X1  g719(.A(G183gat), .B1(new_n910_), .B2(new_n920_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n834_), .A2(new_n479_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n921_), .B1(new_n903_), .B2(new_n922_), .ZN(G1350gat));
  INV_X1    g722(.A(new_n903_), .ZN(new_n924_));
  OAI21_X1  g723(.A(G190gat), .B1(new_n924_), .B2(new_n681_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n903_), .A2(new_n480_), .A3(new_n643_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n925_), .A2(new_n926_), .ZN(G1351gat));
  NOR3_X1   g726(.A1(new_n867_), .A2(new_n651_), .A3(new_n603_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n866_), .A2(new_n928_), .ZN(new_n929_));
  INV_X1    g728(.A(new_n929_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n930_), .A2(new_n402_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g731(.A1(new_n929_), .A2(new_n304_), .ZN(new_n933_));
  MUX2_X1   g732(.A(G204gat), .B(new_n409_), .S(new_n933_), .Z(G1353gat));
  NOR2_X1   g733(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n935_));
  AND2_X1   g734(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n936_));
  NOR4_X1   g735(.A1(new_n929_), .A2(new_n834_), .A3(new_n935_), .A4(new_n936_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n930_), .A2(new_n646_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n937_), .B1(new_n938_), .B2(new_n935_), .ZN(G1354gat));
  XOR2_X1   g738(.A(KEYINPUT127), .B(G218gat), .Z(new_n940_));
  NOR3_X1   g739(.A1(new_n929_), .A2(new_n681_), .A3(new_n940_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n930_), .A2(new_n643_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n941_), .B1(new_n942_), .B2(new_n940_), .ZN(G1355gat));
endmodule


