//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 1 0 1 1 0 0 0 0 0 1 0 1 1 1 1 1 0 1 0 0 0 0 0 0 0 0 0 1 1 0 0 0 1 1 1 1 0 0 1 1 0 1 1 0 1 0 0 1 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n782_, new_n783_, new_n784_,
    new_n785_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n882_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n904_, new_n905_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n912_, new_n913_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_,
    new_n955_, new_n956_, new_n958_, new_n959_, new_n960_, new_n962_,
    new_n963_, new_n964_, new_n965_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n975_, new_n976_,
    new_n977_;
  XNOR2_X1  g000(.A(G15gat), .B(G43gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT83), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT30), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G183gat), .A2(G190gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND3_X1  g006(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n208_));
  OAI211_X1 g007(.A(new_n207_), .B(new_n208_), .C1(G183gat), .C2(G190gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n210_));
  OR3_X1    g009(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n209_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n205_), .A2(KEYINPUT23), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n206_), .A2(G183gat), .A3(G190gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  OR3_X1    g015(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(G183gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT25), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT25), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(G183gat), .ZN(new_n222_));
  INV_X1    g021(.A(G190gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT26), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT26), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(G190gat), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n220_), .A2(new_n222_), .A3(new_n224_), .A4(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G169gat), .A2(G176gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n227_), .A2(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n218_), .B1(new_n232_), .B2(KEYINPUT82), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT25), .B(G183gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT26), .B(G190gat), .ZN(new_n235_));
  AOI22_X1  g034(.A1(new_n234_), .A2(new_n235_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT82), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n213_), .B1(new_n233_), .B2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n204_), .B(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G227gat), .A2(G233gat), .ZN(new_n242_));
  INV_X1    g041(.A(G71gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n241_), .B(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(G127gat), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n247_), .A2(G134gat), .ZN(new_n248_));
  INV_X1    g047(.A(G134gat), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n249_), .A2(G127gat), .ZN(new_n250_));
  INV_X1    g049(.A(G113gat), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n251_), .A2(G120gat), .ZN(new_n252_));
  INV_X1    g051(.A(G120gat), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n253_), .A2(G113gat), .ZN(new_n254_));
  OAI22_X1  g053(.A1(new_n248_), .A2(new_n250_), .B1(new_n252_), .B2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G127gat), .B(G134gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G113gat), .B(G120gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  AND3_X1   g057(.A1(new_n255_), .A2(new_n258_), .A3(KEYINPUT84), .ZN(new_n259_));
  AOI21_X1  g058(.A(KEYINPUT84), .B1(new_n255_), .B2(new_n258_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT31), .ZN(new_n262_));
  INV_X1    g061(.A(G99gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n246_), .B(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G226gat), .A2(G233gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT19), .ZN(new_n268_));
  XOR2_X1   g067(.A(new_n268_), .B(KEYINPUT92), .Z(new_n269_));
  OR2_X1    g068(.A1(G197gat), .A2(G204gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G197gat), .A2(G204gat), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n270_), .A2(KEYINPUT21), .A3(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT21), .ZN(new_n273_));
  AND2_X1   g072(.A1(G197gat), .A2(G204gat), .ZN(new_n274_));
  NOR2_X1   g073(.A1(G197gat), .A2(G204gat), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n273_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G211gat), .B(G218gat), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n272_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  NOR3_X1   g077(.A1(new_n274_), .A2(new_n275_), .A3(new_n273_), .ZN(new_n279_));
  XOR2_X1   g078(.A(G211gat), .B(G218gat), .Z(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n278_), .A2(new_n281_), .ZN(new_n282_));
  AND2_X1   g081(.A1(new_n216_), .A2(new_n217_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n283_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n232_), .A2(KEYINPUT82), .ZN(new_n285_));
  OAI211_X1 g084(.A(new_n282_), .B(new_n212_), .C1(new_n284_), .C2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n286_), .A2(KEYINPUT93), .A3(KEYINPUT20), .ZN(new_n287_));
  INV_X1    g086(.A(new_n282_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n212_), .B1(new_n232_), .B2(new_n218_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n287_), .A2(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(KEYINPUT93), .B1(new_n286_), .B2(KEYINPUT20), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n269_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT20), .B1(new_n288_), .B2(new_n289_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n294_), .B1(new_n240_), .B2(new_n288_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n268_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G8gat), .B(G36gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT18), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G64gat), .B(G92gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n293_), .A2(new_n297_), .A3(new_n302_), .ZN(new_n303_));
  OR2_X1    g102(.A1(new_n303_), .A2(KEYINPUT97), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(KEYINPUT97), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT27), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n286_), .A2(KEYINPUT20), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT93), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n269_), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n309_), .A2(new_n310_), .A3(new_n290_), .A4(new_n287_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n311_), .B1(new_n296_), .B2(new_n295_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n306_), .B1(new_n312_), .B2(new_n301_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n304_), .A2(new_n305_), .A3(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n293_), .A2(new_n297_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(new_n301_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(new_n303_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(new_n306_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n314_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(G141gat), .ZN(new_n320_));
  INV_X1    g119(.A(G148gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT2), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G141gat), .A2(G148gat), .ZN(new_n324_));
  AOI22_X1  g123(.A1(new_n322_), .A2(KEYINPUT3), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT87), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND4_X1  g127(.A1(KEYINPUT87), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT86), .ZN(new_n331_));
  NOR2_X1   g130(.A1(G141gat), .A2(G148gat), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT3), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n331_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  NOR4_X1   g133(.A1(KEYINPUT86), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n325_), .B(new_n330_), .C1(new_n334_), .C2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT88), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(G155gat), .A2(G162gat), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT85), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n341_), .B1(G155gat), .B2(G162gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G155gat), .A2(G162gat), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n343_), .A2(KEYINPUT85), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n340_), .B1(new_n342_), .B2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT89), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n343_), .A2(KEYINPUT85), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n341_), .A2(G155gat), .A3(G162gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT89), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n349_), .A2(new_n350_), .A3(new_n340_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n346_), .A2(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(KEYINPUT86), .B1(new_n322_), .B2(KEYINPUT3), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n332_), .A2(new_n331_), .A3(new_n333_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n355_), .A2(KEYINPUT88), .A3(new_n330_), .A4(new_n325_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n338_), .A2(new_n352_), .A3(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT29), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n349_), .A2(KEYINPUT1), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(new_n340_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n349_), .A2(KEYINPUT1), .ZN(new_n361_));
  OAI211_X1 g160(.A(new_n322_), .B(new_n324_), .C1(new_n360_), .C2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n357_), .A2(new_n358_), .A3(new_n362_), .ZN(new_n363_));
  XOR2_X1   g162(.A(KEYINPUT90), .B(KEYINPUT28), .Z(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G228gat), .A2(G233gat), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT91), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n366_), .B1(new_n282_), .B2(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G22gat), .B(G50gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n365_), .A2(new_n370_), .ZN(new_n371_));
  XOR2_X1   g170(.A(new_n368_), .B(new_n369_), .Z(new_n372_));
  OR2_X1    g171(.A1(new_n363_), .A2(new_n364_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n363_), .A2(new_n364_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n372_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n371_), .A2(new_n375_), .ZN(new_n376_));
  AOI211_X1 g175(.A(KEYINPUT89), .B(new_n339_), .C1(new_n347_), .C2(new_n348_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n350_), .B1(new_n349_), .B2(new_n340_), .ZN(new_n378_));
  OAI22_X1  g177(.A1(new_n336_), .A2(new_n337_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n324_), .A2(new_n323_), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n382_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n383_));
  AOI21_X1  g182(.A(KEYINPUT88), .B1(new_n383_), .B2(new_n330_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n362_), .B1(new_n379_), .B2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT29), .ZN(new_n386_));
  INV_X1    g185(.A(G78gat), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n386_), .A2(new_n387_), .A3(new_n288_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(G106gat), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n387_), .B1(new_n386_), .B2(new_n288_), .ZN(new_n391_));
  NOR3_X1   g190(.A1(new_n389_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n386_), .A2(new_n288_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(G78gat), .ZN(new_n394_));
  AOI21_X1  g193(.A(G106gat), .B1(new_n394_), .B2(new_n388_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n376_), .B1(new_n392_), .B2(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n390_), .B1(new_n389_), .B2(new_n391_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n394_), .A2(G106gat), .A3(new_n388_), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n397_), .A2(new_n398_), .A3(new_n375_), .A4(new_n371_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n396_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n261_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n385_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n255_), .A2(new_n258_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n357_), .A2(new_n362_), .A3(new_n403_), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G225gat), .A2(G233gat), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n402_), .A2(KEYINPUT4), .A3(new_n404_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(KEYINPUT94), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n261_), .B1(new_n357_), .B2(new_n362_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT4), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n409_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  AOI22_X1  g211(.A1(new_n405_), .A2(new_n406_), .B1(new_n407_), .B2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G1gat), .B(G29gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(G85gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(KEYINPUT0), .B(G57gat), .ZN(new_n416_));
  XOR2_X1   g215(.A(new_n415_), .B(new_n416_), .Z(new_n417_));
  AND2_X1   g216(.A1(new_n407_), .A2(new_n412_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n402_), .A2(new_n404_), .A3(new_n406_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(new_n417_), .ZN(new_n420_));
  OAI22_X1  g219(.A1(new_n413_), .A2(new_n417_), .B1(new_n418_), .B2(new_n420_), .ZN(new_n421_));
  NOR4_X1   g220(.A1(new_n266_), .A2(new_n319_), .A3(new_n400_), .A4(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT33), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n423_), .B1(new_n418_), .B2(new_n420_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n417_), .B1(new_n405_), .B2(new_n408_), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n407_), .B(new_n406_), .C1(KEYINPUT4), .C2(new_n402_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  AND3_X1   g226(.A1(new_n419_), .A2(KEYINPUT33), .A3(new_n417_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n407_), .A2(new_n412_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n424_), .A2(new_n427_), .A3(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT95), .B1(new_n431_), .B2(new_n317_), .ZN(new_n432_));
  AND3_X1   g231(.A1(new_n293_), .A2(new_n297_), .A3(new_n302_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n302_), .B1(new_n293_), .B2(new_n297_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  AOI22_X1  g234(.A1(new_n426_), .A2(new_n425_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT95), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n435_), .A2(new_n436_), .A3(new_n437_), .A4(new_n424_), .ZN(new_n438_));
  AND2_X1   g237(.A1(new_n302_), .A2(KEYINPUT32), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n312_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(KEYINPUT96), .ZN(new_n441_));
  OR2_X1    g240(.A1(new_n315_), .A2(new_n439_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT96), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n312_), .A2(new_n443_), .A3(new_n439_), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n441_), .A2(new_n421_), .A3(new_n442_), .A4(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n432_), .A2(new_n438_), .A3(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n400_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n421_), .B1(new_n396_), .B2(new_n399_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n449_), .A2(new_n314_), .A3(KEYINPUT98), .A4(new_n318_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT98), .ZN(new_n451_));
  INV_X1    g250(.A(new_n421_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n400_), .A2(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n451_), .B1(new_n319_), .B2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n448_), .A2(new_n450_), .A3(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n422_), .B1(new_n455_), .B2(new_n266_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G15gat), .B(G22gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(KEYINPUT74), .ZN(new_n458_));
  INV_X1    g257(.A(G1gat), .ZN(new_n459_));
  INV_X1    g258(.A(G8gat), .ZN(new_n460_));
  OAI21_X1  g259(.A(KEYINPUT14), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT75), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n458_), .A2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G1gat), .B(G8gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n465_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n458_), .A2(new_n467_), .A3(new_n463_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G29gat), .B(G36gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G43gat), .B(G50gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n466_), .A2(new_n468_), .A3(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT79), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n466_), .A2(KEYINPUT79), .A3(new_n468_), .A4(new_n471_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G229gat), .A2(G233gat), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n468_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n467_), .B1(new_n458_), .B2(new_n463_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n476_), .B(new_n478_), .C1(new_n481_), .C2(new_n471_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G113gat), .B(G141gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G169gat), .B(G197gat), .ZN(new_n484_));
  XOR2_X1   g283(.A(new_n483_), .B(new_n484_), .Z(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT80), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n466_), .A2(new_n468_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n471_), .B(KEYINPUT15), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n476_), .A2(new_n491_), .ZN(new_n492_));
  OAI211_X1 g291(.A(new_n482_), .B(new_n488_), .C1(new_n492_), .C2(new_n478_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n478_), .B1(new_n476_), .B2(new_n491_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n471_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n495_));
  AOI211_X1 g294(.A(new_n477_), .B(new_n495_), .C1(new_n474_), .C2(new_n475_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n487_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n493_), .A2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT81), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n456_), .A2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G57gat), .B(G64gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT11), .ZN(new_n502_));
  XNOR2_X1  g301(.A(KEYINPUT66), .B(G71gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(G78gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n502_), .A2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n503_), .B(new_n387_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n501_), .A2(KEYINPUT11), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n505_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT17), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G127gat), .B(G155gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT16), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G183gat), .B(G211gat), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT16), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n511_), .B(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n513_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n510_), .B1(new_n514_), .B2(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n481_), .B1(KEYINPUT76), .B2(new_n519_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n516_), .A2(new_n517_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n512_), .A2(new_n513_), .ZN(new_n522_));
  OAI21_X1  g321(.A(KEYINPUT17), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT76), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n489_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G231gat), .A2(G233gat), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n520_), .A2(new_n525_), .A3(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n527_), .B1(new_n520_), .B2(new_n525_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n509_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n530_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n509_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n532_), .A2(new_n533_), .A3(new_n528_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n521_), .A2(new_n522_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(new_n510_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n531_), .A2(new_n534_), .A3(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT77), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT77), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n531_), .A2(new_n534_), .A3(new_n539_), .A4(new_n536_), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n538_), .A2(KEYINPUT78), .A3(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(KEYINPUT78), .B1(new_n538_), .B2(new_n540_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G99gat), .A2(G106gat), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n544_), .A2(KEYINPUT6), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n544_), .A2(KEYINPUT6), .ZN(new_n546_));
  OR2_X1    g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  XOR2_X1   g346(.A(KEYINPUT10), .B(G99gat), .Z(new_n548_));
  XOR2_X1   g347(.A(KEYINPUT64), .B(G106gat), .Z(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  XOR2_X1   g349(.A(G85gat), .B(G92gat), .Z(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(KEYINPUT9), .ZN(new_n552_));
  XNOR2_X1  g351(.A(KEYINPUT65), .B(G85gat), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT9), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n553_), .A2(new_n554_), .A3(G92gat), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n547_), .A2(new_n550_), .A3(new_n552_), .A4(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n557_));
  OR3_X1    g356(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n557_), .B(new_n558_), .C1(new_n545_), .C2(new_n546_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT8), .ZN(new_n560_));
  AND3_X1   g359(.A1(new_n559_), .A2(new_n560_), .A3(new_n551_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n560_), .B1(new_n559_), .B2(new_n551_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n556_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n490_), .A2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G232gat), .A2(G233gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT35), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n471_), .B(new_n556_), .C1(new_n561_), .C2(new_n562_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n564_), .A2(new_n569_), .A3(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n567_), .A2(new_n568_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n572_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n564_), .A2(new_n574_), .A3(new_n569_), .A4(new_n570_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n573_), .A2(KEYINPUT73), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT36), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G190gat), .B(G218gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT71), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT72), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G134gat), .B(G162gat), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n580_), .B(new_n581_), .Z(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n576_), .A2(new_n577_), .A3(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n573_), .A2(new_n582_), .A3(new_n575_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n577_), .B1(new_n576_), .B2(new_n583_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n588_), .A2(KEYINPUT37), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT37), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n590_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n589_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n543_), .A2(new_n592_), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n563_), .A2(new_n509_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT67), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n563_), .A2(new_n509_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n594_), .A2(new_n595_), .A3(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(G230gat), .A2(G233gat), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  OAI211_X1 g398(.A(new_n597_), .B(new_n599_), .C1(new_n595_), .C2(new_n596_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT68), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n596_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT12), .ZN(new_n603_));
  AOI21_X1  g402(.A(KEYINPUT68), .B1(new_n563_), .B2(new_n509_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT12), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n603_), .A2(new_n598_), .A3(new_n606_), .A4(new_n594_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n600_), .A2(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G120gat), .B(G148gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT5), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G176gat), .B(G204gat), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n610_), .B(new_n611_), .Z(new_n612_));
  NAND2_X1  g411(.A1(new_n608_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n612_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n600_), .A2(new_n607_), .A3(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n613_), .A2(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n616_), .B1(KEYINPUT69), .B2(KEYINPUT13), .ZN(new_n617_));
  AND2_X1   g416(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n618_));
  NOR2_X1   g417(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n619_));
  OAI211_X1 g418(.A(new_n613_), .B(new_n615_), .C1(new_n618_), .C2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n617_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n593_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n500_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n421_), .A2(new_n459_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT99), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n627_), .A2(KEYINPUT38), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n621_), .A2(new_n498_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n529_), .A2(new_n530_), .ZN(new_n630_));
  AOI22_X1  g429(.A1(new_n630_), .A2(new_n533_), .B1(new_n510_), .B2(new_n535_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n539_), .B1(new_n631_), .B2(new_n531_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n540_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n629_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n455_), .A2(new_n266_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n422_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT100), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n640_), .A2(new_n641_), .A3(new_n588_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n588_), .ZN(new_n643_));
  OAI21_X1  g442(.A(KEYINPUT100), .B1(new_n456_), .B2(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n637_), .B1(new_n642_), .B2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  OAI21_X1  g445(.A(G1gat), .B1(new_n646_), .B2(new_n452_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n627_), .A2(KEYINPUT38), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n628_), .A2(new_n647_), .A3(new_n648_), .ZN(G1324gat));
  AOI21_X1  g448(.A(new_n460_), .B1(new_n645_), .B2(new_n319_), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n650_), .A2(KEYINPUT39), .ZN(new_n651_));
  INV_X1    g450(.A(new_n624_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n319_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n653_), .A2(G8gat), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n652_), .A2(KEYINPUT101), .A3(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT101), .ZN(new_n656_));
  INV_X1    g455(.A(new_n654_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n656_), .B1(new_n624_), .B2(new_n657_), .ZN(new_n658_));
  AOI22_X1  g457(.A1(new_n650_), .A2(KEYINPUT39), .B1(new_n655_), .B2(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n651_), .A2(new_n659_), .A3(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(new_n651_), .B2(new_n659_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1325gat));
  INV_X1    g462(.A(G15gat), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n664_), .B1(new_n645_), .B2(new_n265_), .ZN(new_n665_));
  XOR2_X1   g464(.A(KEYINPUT103), .B(KEYINPUT41), .Z(new_n666_));
  OR2_X1    g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n652_), .A2(new_n664_), .A3(new_n265_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n665_), .A2(new_n666_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n667_), .A2(new_n668_), .A3(new_n669_), .ZN(G1326gat));
  INV_X1    g469(.A(G22gat), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n652_), .A2(new_n671_), .A3(new_n400_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT42), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n645_), .A2(new_n400_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n673_), .B1(new_n674_), .B2(G22gat), .ZN(new_n675_));
  AOI211_X1 g474(.A(KEYINPUT42), .B(new_n671_), .C1(new_n645_), .C2(new_n400_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n672_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(KEYINPUT104), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT104), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n679_), .B(new_n672_), .C1(new_n675_), .C2(new_n676_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(G1327gat));
  INV_X1    g480(.A(new_n543_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n682_), .A2(new_n621_), .A3(new_n643_), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n456_), .A2(new_n683_), .A3(new_n499_), .ZN(new_n684_));
  AOI21_X1  g483(.A(G29gat), .B1(new_n684_), .B2(new_n421_), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n543_), .A2(new_n629_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT43), .ZN(new_n688_));
  INV_X1    g487(.A(new_n592_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n640_), .B2(new_n689_), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n456_), .A2(KEYINPUT43), .A3(new_n592_), .ZN(new_n691_));
  OAI211_X1 g490(.A(KEYINPUT44), .B(new_n687_), .C1(new_n690_), .C2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(KEYINPUT105), .ZN(new_n693_));
  OAI21_X1  g492(.A(KEYINPUT43), .B1(new_n456_), .B2(new_n592_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n449_), .A2(new_n318_), .A3(new_n314_), .ZN(new_n695_));
  AOI22_X1  g494(.A1(new_n446_), .A2(new_n447_), .B1(new_n695_), .B2(new_n451_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n265_), .B1(new_n696_), .B2(new_n450_), .ZN(new_n697_));
  OAI211_X1 g496(.A(new_n688_), .B(new_n689_), .C1(new_n697_), .C2(new_n422_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n686_), .B1(new_n694_), .B2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT105), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n699_), .A2(new_n700_), .A3(KEYINPUT44), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n693_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n699_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n702_), .A2(new_n705_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n421_), .A2(G29gat), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n685_), .B1(new_n706_), .B2(new_n707_), .ZN(G1328gat));
  INV_X1    g507(.A(KEYINPUT46), .ZN(new_n709_));
  INV_X1    g508(.A(G36gat), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n319_), .B1(new_n699_), .B2(KEYINPUT44), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n710_), .B1(new_n702_), .B2(new_n712_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n653_), .A2(G36gat), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n684_), .A2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT106), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT106), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n684_), .A2(new_n717_), .A3(new_n714_), .ZN(new_n718_));
  AOI21_X1  g517(.A(KEYINPUT45), .B1(new_n716_), .B2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n716_), .A2(KEYINPUT45), .A3(new_n718_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n709_), .B1(new_n713_), .B2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n721_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n724_), .A2(new_n719_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n711_), .B1(new_n693_), .B2(new_n701_), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n725_), .B(KEYINPUT46), .C1(new_n710_), .C2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n723_), .A2(new_n727_), .ZN(G1329gat));
  AND2_X1   g527(.A1(new_n265_), .A2(G43gat), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n692_), .A2(KEYINPUT105), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n700_), .B1(new_n699_), .B2(KEYINPUT44), .ZN(new_n731_));
  OAI211_X1 g530(.A(new_n705_), .B(new_n729_), .C1(new_n730_), .C2(new_n731_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n684_), .A2(new_n265_), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n733_), .A2(G43gat), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT47), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT47), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n732_), .A2(new_n737_), .A3(new_n734_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(G1330gat));
  AOI21_X1  g538(.A(G50gat), .B1(new_n684_), .B2(new_n400_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n400_), .A2(G50gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n706_), .B2(new_n741_), .ZN(G1331gat));
  NAND2_X1  g541(.A1(new_n642_), .A2(new_n644_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT78), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n744_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n538_), .A2(KEYINPUT78), .A3(new_n540_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n745_), .A2(new_n499_), .A3(new_n746_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n747_), .A2(new_n621_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n743_), .A2(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(G57gat), .B1(new_n749_), .B2(new_n452_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n456_), .A2(new_n498_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n593_), .A2(new_n621_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  OR3_X1    g552(.A1(new_n753_), .A2(G57gat), .A3(new_n452_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n750_), .A2(new_n754_), .ZN(G1332gat));
  OAI21_X1  g554(.A(G64gat), .B1(new_n749_), .B2(new_n653_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n756_), .A2(KEYINPUT48), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n756_), .A2(KEYINPUT48), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n653_), .A2(G64gat), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT107), .ZN(new_n760_));
  OAI22_X1  g559(.A1(new_n757_), .A2(new_n758_), .B1(new_n753_), .B2(new_n760_), .ZN(G1333gat));
  INV_X1    g560(.A(new_n753_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n762_), .A2(new_n243_), .A3(new_n265_), .ZN(new_n763_));
  OAI21_X1  g562(.A(G71gat), .B1(new_n749_), .B2(new_n266_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n764_), .A2(KEYINPUT49), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n764_), .A2(KEYINPUT49), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n763_), .B1(new_n765_), .B2(new_n766_), .ZN(G1334gat));
  NAND3_X1  g566(.A1(new_n762_), .A2(new_n387_), .A3(new_n400_), .ZN(new_n768_));
  OAI21_X1  g567(.A(G78gat), .B1(new_n749_), .B2(new_n447_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n769_), .A2(KEYINPUT50), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n769_), .A2(KEYINPUT50), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n768_), .B1(new_n770_), .B2(new_n771_), .ZN(G1335gat));
  NOR3_X1   g571(.A1(new_n543_), .A2(new_n621_), .A3(new_n588_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n751_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(G85gat), .B1(new_n775_), .B2(new_n421_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n694_), .A2(new_n698_), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n543_), .A2(new_n498_), .A3(new_n621_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n421_), .A2(new_n553_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n776_), .B1(new_n779_), .B2(new_n780_), .ZN(G1336gat));
  INV_X1    g580(.A(G92gat), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n782_), .B1(new_n774_), .B2(new_n653_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT108), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n653_), .A2(new_n782_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n784_), .B1(new_n779_), .B2(new_n785_), .ZN(G1337gat));
  NAND3_X1  g585(.A1(new_n775_), .A2(new_n265_), .A3(new_n548_), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n777_), .A2(new_n265_), .A3(new_n778_), .ZN(new_n788_));
  OAI211_X1 g587(.A(KEYINPUT110), .B(new_n787_), .C1(new_n788_), .C2(new_n263_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT109), .ZN(new_n790_));
  NAND2_X1  g589(.A1(KEYINPUT109), .A2(KEYINPUT51), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n787_), .B(new_n791_), .C1(new_n788_), .C2(new_n263_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT51), .ZN(new_n793_));
  AOI22_X1  g592(.A1(new_n790_), .A2(new_n792_), .B1(new_n793_), .B2(new_n789_), .ZN(G1338gat));
  NAND2_X1  g593(.A1(new_n400_), .A2(new_n549_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n774_), .A2(new_n795_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT111), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT112), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n777_), .A2(new_n400_), .A3(new_n778_), .ZN(new_n801_));
  OAI21_X1  g600(.A(G106gat), .B1(new_n798_), .B2(KEYINPUT112), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n800_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n797_), .A2(new_n803_), .ZN(new_n804_));
  NOR3_X1   g603(.A1(new_n801_), .A2(new_n800_), .A3(new_n802_), .ZN(new_n805_));
  OAI21_X1  g604(.A(KEYINPUT53), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n805_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n807_), .A2(new_n808_), .A3(new_n803_), .A4(new_n797_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n806_), .A2(new_n809_), .ZN(G1339gat));
  INV_X1    g609(.A(KEYINPUT117), .ZN(new_n811_));
  XNOR2_X1  g610(.A(KEYINPUT116), .B(KEYINPUT58), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n594_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n604_), .A2(new_n605_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n599_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT114), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n607_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n814_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n820_), .A2(KEYINPUT55), .A3(new_n598_), .A4(new_n606_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT114), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n822_), .B(new_n599_), .C1(new_n814_), .C2(new_n815_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n817_), .A2(new_n819_), .A3(new_n821_), .A4(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n612_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT56), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n824_), .A2(KEYINPUT56), .A3(new_n612_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n477_), .B1(new_n476_), .B2(new_n491_), .ZN(new_n830_));
  AOI211_X1 g629(.A(new_n478_), .B(new_n495_), .C1(new_n474_), .C2(new_n475_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n486_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n485_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n832_), .A2(new_n833_), .A3(new_n615_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT115), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n832_), .A2(new_n833_), .A3(new_n615_), .A4(KEYINPUT115), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n813_), .B1(new_n829_), .B2(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n811_), .B1(new_n839_), .B2(new_n592_), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n827_), .A2(new_n828_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(KEYINPUT58), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n689_), .B(KEYINPUT117), .C1(new_n841_), .C2(new_n813_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n840_), .A2(new_n842_), .A3(new_n843_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n498_), .A2(new_n615_), .ZN(new_n845_));
  AND3_X1   g644(.A1(new_n824_), .A2(KEYINPUT56), .A3(new_n612_), .ZN(new_n846_));
  AOI21_X1  g645(.A(KEYINPUT56), .B1(new_n824_), .B2(new_n612_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n845_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n616_), .A2(new_n832_), .A3(new_n833_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(KEYINPUT57), .B1(new_n850_), .B2(new_n588_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT57), .ZN(new_n852_));
  AOI211_X1 g651(.A(new_n852_), .B(new_n643_), .C1(new_n848_), .C2(new_n849_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n851_), .A2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n543_), .B1(new_n844_), .B2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT113), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n856_), .B1(new_n543_), .B2(new_n499_), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n745_), .A2(new_n499_), .A3(new_n856_), .A4(new_n746_), .ZN(new_n858_));
  AOI22_X1  g657(.A1(new_n589_), .A2(new_n591_), .B1(new_n617_), .B2(new_n620_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(KEYINPUT54), .B1(new_n857_), .B2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n747_), .A2(KEYINPUT113), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT54), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n862_), .A2(new_n863_), .A3(new_n858_), .A4(new_n859_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n861_), .A2(new_n864_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n855_), .A2(new_n865_), .ZN(new_n866_));
  NOR4_X1   g665(.A1(new_n266_), .A2(new_n319_), .A3(new_n400_), .A4(new_n452_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT59), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n866_), .A2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n844_), .A2(new_n854_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n635_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n861_), .A2(new_n864_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n872_), .A2(KEYINPUT118), .A3(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT118), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n634_), .B1(new_n844_), .B2(new_n854_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(new_n876_), .B2(new_n865_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n874_), .A2(new_n877_), .A3(new_n867_), .ZN(new_n878_));
  AOI211_X1 g677(.A(new_n499_), .B(new_n870_), .C1(new_n878_), .C2(KEYINPUT59), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n498_), .A2(new_n251_), .ZN(new_n880_));
  OAI22_X1  g679(.A1(new_n879_), .A2(new_n251_), .B1(new_n878_), .B2(new_n880_), .ZN(G1340gat));
  AOI211_X1 g680(.A(new_n621_), .B(new_n870_), .C1(new_n878_), .C2(KEYINPUT59), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n253_), .B1(new_n621_), .B2(KEYINPUT60), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n883_), .B1(KEYINPUT60), .B2(new_n253_), .ZN(new_n884_));
  OAI22_X1  g683(.A1(new_n882_), .A2(new_n253_), .B1(new_n878_), .B2(new_n884_), .ZN(G1341gat));
  AOI211_X1 g684(.A(new_n635_), .B(new_n870_), .C1(new_n878_), .C2(KEYINPUT59), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n543_), .A2(new_n247_), .ZN(new_n887_));
  OAI22_X1  g686(.A1(new_n886_), .A2(new_n247_), .B1(new_n878_), .B2(new_n887_), .ZN(G1342gat));
  OAI21_X1  g687(.A(new_n249_), .B1(new_n878_), .B2(new_n588_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT119), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  OAI211_X1 g690(.A(KEYINPUT119), .B(new_n249_), .C1(new_n878_), .C2(new_n588_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n870_), .B1(new_n878_), .B2(KEYINPUT59), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n592_), .A2(new_n249_), .ZN(new_n894_));
  AOI22_X1  g693(.A1(new_n891_), .A2(new_n892_), .B1(new_n893_), .B2(new_n894_), .ZN(G1343gat));
  NOR2_X1   g694(.A1(new_n447_), .A2(new_n265_), .ZN(new_n896_));
  AND3_X1   g695(.A1(new_n874_), .A2(new_n877_), .A3(new_n896_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n319_), .A2(new_n452_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n498_), .ZN(new_n900_));
  OAI21_X1  g699(.A(G141gat), .B1(new_n899_), .B2(new_n900_), .ZN(new_n901_));
  NAND4_X1  g700(.A1(new_n897_), .A2(new_n320_), .A3(new_n498_), .A4(new_n898_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1344gat));
  OAI21_X1  g702(.A(G148gat), .B1(new_n899_), .B2(new_n621_), .ZN(new_n904_));
  NAND4_X1  g703(.A1(new_n897_), .A2(new_n321_), .A3(new_n622_), .A4(new_n898_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(G1345gat));
  XNOR2_X1  g705(.A(KEYINPUT61), .B(G155gat), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n907_), .B1(new_n899_), .B2(new_n682_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n907_), .ZN(new_n909_));
  NAND4_X1  g708(.A1(new_n897_), .A2(new_n543_), .A3(new_n898_), .A4(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n908_), .A2(new_n910_), .ZN(G1346gat));
  OAI21_X1  g710(.A(G162gat), .B1(new_n899_), .B2(new_n592_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n588_), .A2(G162gat), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n897_), .A2(new_n898_), .A3(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n912_), .A2(new_n914_), .ZN(G1347gat));
  OR2_X1    g714(.A1(new_n855_), .A2(new_n865_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n653_), .A2(new_n421_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(new_n265_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n918_), .A2(new_n400_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n916_), .A2(new_n498_), .A3(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(G169gat), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(KEYINPUT120), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT120), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n920_), .A2(new_n923_), .A3(G169gat), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n922_), .A2(KEYINPUT62), .A3(new_n924_), .ZN(new_n925_));
  XOR2_X1   g724(.A(KEYINPUT22), .B(G169gat), .Z(new_n926_));
  NOR2_X1   g725(.A1(new_n920_), .A2(new_n926_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n923_), .B1(new_n920_), .B2(G169gat), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT62), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n927_), .B1(new_n928_), .B2(new_n929_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n925_), .A2(new_n930_), .ZN(G1348gat));
  AND3_X1   g730(.A1(new_n874_), .A2(new_n877_), .A3(new_n447_), .ZN(new_n932_));
  INV_X1    g731(.A(G176gat), .ZN(new_n933_));
  NOR3_X1   g732(.A1(new_n918_), .A2(new_n933_), .A3(new_n621_), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n916_), .A2(new_n622_), .A3(new_n919_), .ZN(new_n935_));
  AOI22_X1  g734(.A1(new_n932_), .A2(new_n934_), .B1(new_n935_), .B2(new_n933_), .ZN(G1349gat));
  NOR2_X1   g735(.A1(new_n918_), .A2(new_n682_), .ZN(new_n937_));
  NAND4_X1  g736(.A1(new_n874_), .A2(new_n877_), .A3(new_n447_), .A4(new_n937_), .ZN(new_n938_));
  AND2_X1   g737(.A1(new_n938_), .A2(new_n219_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n635_), .A2(new_n234_), .ZN(new_n940_));
  OAI211_X1 g739(.A(new_n919_), .B(new_n940_), .C1(new_n855_), .C2(new_n865_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(KEYINPUT121), .ZN(new_n942_));
  OAI21_X1  g741(.A(KEYINPUT122), .B1(new_n939_), .B2(new_n942_), .ZN(new_n943_));
  INV_X1    g742(.A(KEYINPUT121), .ZN(new_n944_));
  XNOR2_X1  g743(.A(new_n941_), .B(new_n944_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n938_), .A2(new_n219_), .ZN(new_n946_));
  INV_X1    g745(.A(KEYINPUT122), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n945_), .A2(new_n946_), .A3(new_n947_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n943_), .A2(new_n948_), .ZN(G1350gat));
  NAND3_X1  g748(.A1(new_n916_), .A2(new_n689_), .A3(new_n919_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n950_), .A2(G190gat), .ZN(new_n951_));
  NAND4_X1  g750(.A1(new_n916_), .A2(new_n235_), .A3(new_n643_), .A4(new_n919_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n951_), .A2(new_n952_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n953_), .A2(KEYINPUT123), .ZN(new_n954_));
  INV_X1    g753(.A(KEYINPUT123), .ZN(new_n955_));
  NAND3_X1  g754(.A1(new_n951_), .A2(new_n955_), .A3(new_n952_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n954_), .A2(new_n956_), .ZN(G1351gat));
  NAND4_X1  g756(.A1(new_n874_), .A2(new_n877_), .A3(new_n896_), .A4(new_n917_), .ZN(new_n958_));
  NOR2_X1   g757(.A1(new_n958_), .A2(new_n900_), .ZN(new_n959_));
  INV_X1    g758(.A(G197gat), .ZN(new_n960_));
  XNOR2_X1  g759(.A(new_n959_), .B(new_n960_), .ZN(G1352gat));
  NOR2_X1   g760(.A1(new_n958_), .A2(new_n621_), .ZN(new_n962_));
  AND2_X1   g761(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n963_));
  NOR2_X1   g762(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n964_));
  OAI21_X1  g763(.A(new_n962_), .B1(new_n963_), .B2(new_n964_), .ZN(new_n965_));
  OAI21_X1  g764(.A(new_n965_), .B1(new_n962_), .B2(new_n964_), .ZN(G1353gat));
  NAND2_X1  g765(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n634_), .A2(new_n967_), .ZN(new_n968_));
  NOR2_X1   g767(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n969_));
  AND2_X1   g768(.A1(new_n969_), .A2(KEYINPUT125), .ZN(new_n970_));
  NOR3_X1   g769(.A1(new_n958_), .A2(new_n968_), .A3(new_n970_), .ZN(new_n971_));
  OR2_X1    g770(.A1(new_n958_), .A2(new_n968_), .ZN(new_n972_));
  XNOR2_X1  g771(.A(new_n969_), .B(KEYINPUT125), .ZN(new_n973_));
  AOI21_X1  g772(.A(new_n971_), .B1(new_n972_), .B2(new_n973_), .ZN(G1354gat));
  XOR2_X1   g773(.A(KEYINPUT126), .B(G218gat), .Z(new_n975_));
  NOR3_X1   g774(.A1(new_n958_), .A2(new_n592_), .A3(new_n975_), .ZN(new_n976_));
  NAND3_X1  g775(.A1(new_n897_), .A2(new_n643_), .A3(new_n917_), .ZN(new_n977_));
  AOI21_X1  g776(.A(new_n976_), .B1(new_n977_), .B2(new_n975_), .ZN(G1355gat));
endmodule


