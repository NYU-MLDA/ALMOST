//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 1 0 1 1 0 0 1 1 0 0 0 1 1 0 0 0 1 1 0 1 0 1 0 1 0 1 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 0 1 1 0 1 0 0 1 1 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n761_, new_n762_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n783_, new_n784_, new_n785_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n798_, new_n799_, new_n800_, new_n802_, new_n803_,
    new_n804_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n913_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n923_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n942_, new_n943_, new_n944_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n957_, new_n958_,
    new_n959_, new_n960_, new_n961_, new_n963_, new_n964_, new_n966_,
    new_n967_, new_n968_, new_n969_, new_n970_, new_n971_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n980_,
    new_n981_, new_n982_, new_n983_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n990_, new_n991_;
  XNOR2_X1  g000(.A(G120gat), .B(G148gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT5), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G176gat), .B(G204gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(KEYINPUT69), .ZN(new_n206_));
  INV_X1    g005(.A(G57gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n207_), .A2(G64gat), .ZN(new_n208_));
  INV_X1    g007(.A(G64gat), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n209_), .A2(G57gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n206_), .B1(new_n208_), .B2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT11), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n209_), .A2(G57gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n207_), .A2(G64gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n213_), .A2(new_n214_), .A3(KEYINPUT69), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n211_), .A2(new_n212_), .A3(new_n215_), .ZN(new_n216_));
  XOR2_X1   g015(.A(G71gat), .B(G78gat), .Z(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT70), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n211_), .A2(new_n215_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n219_), .B1(new_n220_), .B2(KEYINPUT11), .ZN(new_n221_));
  AOI211_X1 g020(.A(KEYINPUT70), .B(new_n212_), .C1(new_n211_), .C2(new_n215_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n218_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  AND3_X1   g022(.A1(new_n213_), .A2(new_n214_), .A3(KEYINPUT69), .ZN(new_n224_));
  AOI21_X1  g023(.A(KEYINPUT69), .B1(new_n213_), .B2(new_n214_), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT11), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT70), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n220_), .A2(new_n219_), .A3(KEYINPUT11), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n227_), .A2(new_n228_), .A3(new_n216_), .A4(new_n217_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G85gat), .A2(G92gat), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(G85gat), .A2(G92gat), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(KEYINPUT68), .A2(KEYINPUT6), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(KEYINPUT68), .A2(KEYINPUT6), .ZN(new_n236_));
  OAI211_X1 g035(.A(G99gat), .B(G106gat), .C1(new_n235_), .C2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n236_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G99gat), .A2(G106gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n238_), .A2(new_n239_), .A3(new_n234_), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n237_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  NOR4_X1   g041(.A1(KEYINPUT67), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n244_));
  NOR2_X1   g043(.A1(G99gat), .A2(G106gat), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT7), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n244_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n243_), .A2(new_n247_), .ZN(new_n248_));
  OAI211_X1 g047(.A(KEYINPUT8), .B(new_n233_), .C1(new_n242_), .C2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT6), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n239_), .A2(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n251_), .A2(new_n241_), .A3(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n233_), .B1(new_n248_), .B2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT8), .ZN(new_n255_));
  NAND3_X1  g054(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT66), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n256_), .B1(new_n232_), .B2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT65), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT9), .ZN(new_n260_));
  AND3_X1   g059(.A1(new_n230_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n259_), .B1(new_n230_), .B2(new_n260_), .ZN(new_n262_));
  OAI221_X1 g061(.A(new_n258_), .B1(new_n257_), .B2(new_n256_), .C1(new_n261_), .C2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n251_), .A2(new_n252_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT10), .B(G99gat), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(G106gat), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n264_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  AOI22_X1  g067(.A1(new_n254_), .A2(new_n255_), .B1(new_n263_), .B2(new_n268_), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n223_), .A2(new_n229_), .A3(new_n249_), .A4(new_n269_), .ZN(new_n270_));
  OR2_X1    g069(.A1(new_n270_), .A2(KEYINPUT71), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n254_), .A2(new_n255_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n263_), .A2(new_n268_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n272_), .A2(new_n249_), .A3(new_n273_), .ZN(new_n274_));
  NOR3_X1   g073(.A1(new_n221_), .A2(new_n222_), .A3(new_n218_), .ZN(new_n275_));
  AOI22_X1  g074(.A1(new_n227_), .A2(new_n228_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n274_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT72), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n223_), .A2(new_n229_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n280_), .A2(KEYINPUT72), .A3(new_n274_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n270_), .A2(KEYINPUT71), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n271_), .A2(new_n279_), .A3(new_n281_), .A4(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G230gat), .A2(G233gat), .ZN(new_n284_));
  XOR2_X1   g083(.A(new_n284_), .B(KEYINPUT64), .Z(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n283_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n277_), .A2(KEYINPUT12), .A3(new_n270_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT12), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n280_), .A2(new_n290_), .A3(new_n274_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n286_), .B1(new_n289_), .B2(new_n291_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n205_), .B1(new_n288_), .B2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n289_), .A2(new_n291_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(new_n285_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n205_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n287_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n293_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT13), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n293_), .A2(KEYINPUT13), .A3(new_n297_), .ZN(new_n301_));
  AND2_X1   g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  XOR2_X1   g102(.A(G29gat), .B(G36gat), .Z(new_n304_));
  XOR2_X1   g103(.A(G43gat), .B(G50gat), .Z(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(KEYINPUT15), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT15), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n306_), .A2(new_n309_), .ZN(new_n310_));
  AND2_X1   g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(new_n274_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G232gat), .A2(G233gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT34), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT35), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n315_), .A2(new_n316_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n269_), .A2(new_n306_), .A3(new_n249_), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n312_), .A2(new_n318_), .A3(new_n319_), .A4(new_n320_), .ZN(new_n321_));
  XOR2_X1   g120(.A(new_n321_), .B(KEYINPUT74), .Z(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n319_), .ZN(new_n323_));
  OR2_X1    g122(.A1(new_n323_), .A2(KEYINPUT73), .ZN(new_n324_));
  AOI22_X1  g123(.A1(new_n323_), .A2(KEYINPUT73), .B1(new_n311_), .B2(new_n274_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n318_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT36), .ZN(new_n328_));
  XOR2_X1   g127(.A(G134gat), .B(G162gat), .Z(new_n329_));
  XNOR2_X1  g128(.A(G190gat), .B(G218gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n322_), .A2(new_n327_), .A3(new_n328_), .A4(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n328_), .ZN(new_n333_));
  OR2_X1    g132(.A1(new_n331_), .A2(new_n328_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n321_), .B(KEYINPUT74), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n333_), .B(new_n334_), .C1(new_n335_), .C2(new_n326_), .ZN(new_n336_));
  AND3_X1   g135(.A1(new_n332_), .A2(KEYINPUT37), .A3(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(KEYINPUT37), .B1(new_n332_), .B2(new_n336_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT75), .B(G1gat), .ZN(new_n340_));
  INV_X1    g139(.A(G8gat), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT14), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G15gat), .B(G22gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G1gat), .B(G8gat), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n342_), .A2(new_n343_), .A3(new_n345_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G231gat), .A2(G233gat), .ZN(new_n350_));
  XOR2_X1   g149(.A(new_n349_), .B(new_n350_), .Z(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(new_n280_), .ZN(new_n352_));
  XOR2_X1   g151(.A(G127gat), .B(G155gat), .Z(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT16), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G183gat), .B(G211gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT17), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  AND2_X1   g157(.A1(new_n356_), .A2(new_n357_), .ZN(new_n359_));
  OR3_X1    g158(.A1(new_n352_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n352_), .A2(new_n358_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n339_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G226gat), .A2(G233gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT19), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT25), .B(G183gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT26), .B(G190gat), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT24), .ZN(new_n369_));
  NOR2_X1   g168(.A1(G169gat), .A2(G176gat), .ZN(new_n370_));
  AOI22_X1  g169(.A1(new_n367_), .A2(new_n368_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT79), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n373_));
  AND2_X1   g172(.A1(G169gat), .A2(G176gat), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n372_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(G169gat), .ZN(new_n376_));
  INV_X1    g175(.A(G176gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G169gat), .A2(G176gat), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n378_), .A2(KEYINPUT79), .A3(KEYINPUT24), .A4(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n375_), .A2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n371_), .A2(new_n381_), .A3(new_n385_), .ZN(new_n386_));
  OR2_X1    g185(.A1(G197gat), .A2(G204gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G197gat), .A2(G204gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT21), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n387_), .A2(KEYINPUT21), .A3(new_n388_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G211gat), .B(G218gat), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n391_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  OR2_X1    g193(.A1(new_n392_), .A2(new_n393_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G183gat), .A2(G190gat), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT23), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(G183gat), .ZN(new_n399_));
  INV_X1    g198(.A(G190gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n398_), .A2(new_n401_), .A3(new_n382_), .ZN(new_n402_));
  OAI21_X1  g201(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT22), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n404_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n402_), .A2(new_n403_), .A3(new_n405_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n386_), .A2(new_n394_), .A3(new_n395_), .A4(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT20), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n405_), .A2(new_n403_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n402_), .A2(KEYINPUT89), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT89), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n398_), .A2(new_n401_), .A3(new_n411_), .A4(new_n382_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n409_), .B1(new_n410_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n378_), .A2(KEYINPUT24), .A3(new_n379_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n371_), .A2(new_n385_), .A3(new_n415_), .ZN(new_n416_));
  AOI22_X1  g215(.A1(new_n414_), .A2(new_n416_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n366_), .B1(new_n408_), .B2(new_n417_), .ZN(new_n418_));
  XOR2_X1   g217(.A(G8gat), .B(G36gat), .Z(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(KEYINPUT18), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G64gat), .B(G92gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT20), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n386_), .A2(new_n406_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n394_), .A2(new_n395_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n423_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n366_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n394_), .A2(new_n395_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n428_), .A2(new_n414_), .A3(new_n416_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n426_), .A2(new_n427_), .A3(new_n429_), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n418_), .A2(new_n422_), .A3(new_n430_), .ZN(new_n431_));
  XOR2_X1   g230(.A(new_n431_), .B(KEYINPUT101), .Z(new_n432_));
  NAND2_X1  g231(.A1(new_n399_), .A2(KEYINPUT25), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT25), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(G183gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n400_), .A2(KEYINPUT26), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT26), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(G190gat), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n433_), .A2(new_n435_), .A3(new_n436_), .A4(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n370_), .A2(new_n369_), .ZN(new_n440_));
  AND4_X1   g239(.A1(new_n385_), .A2(new_n439_), .A3(new_n440_), .A4(new_n415_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n425_), .B1(new_n413_), .B2(new_n441_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n442_), .A2(new_n407_), .A3(KEYINPUT20), .A4(new_n427_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(KEYINPUT97), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n409_), .B1(new_n385_), .B2(new_n401_), .ZN(new_n445_));
  AND3_X1   g244(.A1(new_n439_), .A2(new_n385_), .A3(new_n440_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n445_), .B1(new_n446_), .B2(new_n381_), .ZN(new_n447_));
  OAI21_X1  g246(.A(KEYINPUT20), .B1(new_n447_), .B2(new_n428_), .ZN(new_n448_));
  NOR3_X1   g247(.A1(new_n425_), .A2(new_n413_), .A3(new_n441_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n366_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  AND2_X1   g249(.A1(new_n444_), .A2(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n423_), .B1(new_n447_), .B2(new_n428_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT97), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n452_), .A2(new_n453_), .A3(new_n427_), .A4(new_n442_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n422_), .B1(new_n451_), .B2(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(KEYINPUT27), .B1(new_n432_), .B2(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n422_), .B1(new_n418_), .B2(new_n430_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n431_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  OR2_X1    g258(.A1(new_n459_), .A2(KEYINPUT27), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n456_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT85), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  OAI211_X1 g264(.A(KEYINPUT85), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(G141gat), .ZN(new_n468_));
  INV_X1    g267(.A(G148gat), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n468_), .A2(new_n469_), .A3(KEYINPUT84), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT84), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n471_), .B1(G141gat), .B2(G148gat), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT3), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n470_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G141gat), .A2(G148gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT86), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT2), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT2), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n475_), .A2(KEYINPUT86), .A3(new_n478_), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n467_), .A2(new_n474_), .A3(new_n477_), .A4(new_n479_), .ZN(new_n480_));
  XOR2_X1   g279(.A(G155gat), .B(G162gat), .Z(new_n481_));
  NOR2_X1   g280(.A1(G141gat), .A2(G148gat), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n475_), .B1(new_n482_), .B2(KEYINPUT82), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n483_), .B1(KEYINPUT82), .B2(new_n482_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G155gat), .A2(G162gat), .ZN(new_n485_));
  OR3_X1    g284(.A1(new_n485_), .A2(KEYINPUT83), .A3(KEYINPUT1), .ZN(new_n486_));
  NOR2_X1   g285(.A1(G155gat), .A2(G162gat), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n485_), .B1(new_n487_), .B2(KEYINPUT1), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT83), .B1(new_n485_), .B2(KEYINPUT1), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n486_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  AOI22_X1  g289(.A1(new_n480_), .A2(new_n481_), .B1(new_n484_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT29), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n425_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(G228gat), .ZN(new_n494_));
  INV_X1    g293(.A(G233gat), .ZN(new_n495_));
  OAI21_X1  g294(.A(KEYINPUT88), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n493_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(G78gat), .ZN(new_n498_));
  INV_X1    g297(.A(G78gat), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n493_), .A2(new_n499_), .A3(new_n496_), .ZN(new_n500_));
  AOI21_X1  g299(.A(G106gat), .B1(new_n498_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n498_), .A2(G106gat), .A3(new_n500_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n491_), .A2(new_n492_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G22gat), .B(G50gat), .ZN(new_n505_));
  XOR2_X1   g304(.A(new_n504_), .B(new_n505_), .Z(new_n506_));
  AND3_X1   g305(.A1(new_n502_), .A2(new_n503_), .A3(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n506_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n509_));
  NOR3_X1   g308(.A1(new_n494_), .A2(new_n495_), .A3(KEYINPUT88), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  OR3_X1    g311(.A1(new_n507_), .A2(new_n508_), .A3(new_n512_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n512_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n462_), .A2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G127gat), .B(G134gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G113gat), .B(G120gat), .ZN(new_n518_));
  AND2_X1   g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n517_), .A2(new_n518_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT31), .ZN(new_n523_));
  OAI21_X1  g322(.A(KEYINPUT81), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n524_), .B1(new_n523_), .B2(new_n522_), .ZN(new_n525_));
  XOR2_X1   g324(.A(G71gat), .B(G99gat), .Z(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G227gat), .A2(G233gat), .ZN(new_n528_));
  INV_X1    g327(.A(G15gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT30), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n424_), .B(new_n531_), .ZN(new_n532_));
  XOR2_X1   g331(.A(KEYINPUT80), .B(G43gat), .Z(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n527_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n527_), .A2(new_n534_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G1gat), .B(G29gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(G85gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(KEYINPUT0), .B(G57gat), .ZN(new_n540_));
  XOR2_X1   g339(.A(new_n539_), .B(new_n540_), .Z(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G225gat), .A2(G233gat), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT90), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n544_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n517_), .ZN(new_n546_));
  XOR2_X1   g345(.A(G113gat), .B(G120gat), .Z(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n517_), .A2(new_n518_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n548_), .A2(KEYINPUT90), .A3(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n545_), .B1(new_n491_), .B2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n480_), .A2(new_n481_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n484_), .A2(new_n490_), .ZN(new_n553_));
  AND4_X1   g352(.A1(new_n552_), .A2(new_n545_), .A3(new_n553_), .A4(new_n550_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n543_), .B1(new_n551_), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(KEYINPUT92), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n552_), .A2(new_n553_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n557_), .A2(new_n544_), .A3(new_n522_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n491_), .A2(new_n545_), .A3(new_n550_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT92), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n560_), .A2(new_n561_), .A3(new_n543_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n556_), .A2(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(KEYINPUT4), .B1(new_n551_), .B2(new_n554_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n543_), .ZN(new_n565_));
  XOR2_X1   g364(.A(KEYINPUT91), .B(KEYINPUT4), .Z(new_n566_));
  NAND3_X1  g365(.A1(new_n557_), .A2(new_n521_), .A3(new_n566_), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n564_), .A2(new_n565_), .A3(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n542_), .B1(new_n563_), .B2(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n564_), .A2(new_n565_), .A3(new_n567_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n570_), .A2(new_n556_), .A3(new_n541_), .A4(new_n562_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n537_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n516_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n515_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT33), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n458_), .B1(new_n571_), .B2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n564_), .A2(new_n543_), .A3(new_n567_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n541_), .B1(new_n560_), .B2(new_n565_), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n579_), .A2(KEYINPUT96), .A3(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(KEYINPUT96), .B1(new_n579_), .B2(new_n580_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n578_), .A2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(KEYINPUT94), .B(KEYINPUT33), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n571_), .A2(KEYINPUT93), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n561_), .B1(new_n560_), .B2(new_n543_), .ZN(new_n588_));
  AOI211_X1 g387(.A(KEYINPUT92), .B(new_n565_), .C1(new_n558_), .C2(new_n559_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT93), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n590_), .A2(new_n591_), .A3(new_n541_), .A4(new_n570_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n586_), .B1(new_n587_), .B2(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n584_), .B1(new_n593_), .B2(KEYINPUT95), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n593_), .A2(KEYINPUT95), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n418_), .A2(new_n430_), .ZN(new_n597_));
  AND2_X1   g396(.A1(new_n422_), .A2(KEYINPUT32), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n599_), .B1(new_n569_), .B2(new_n571_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n444_), .A2(new_n450_), .A3(new_n454_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(new_n598_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT98), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT98), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n601_), .A2(new_n604_), .A3(new_n598_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n603_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n600_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(KEYINPUT99), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT99), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n600_), .A2(new_n609_), .A3(new_n606_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n610_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n576_), .B1(new_n596_), .B2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT100), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT95), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n587_), .A2(new_n592_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n615_), .B1(new_n616_), .B2(new_n586_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n593_), .A2(KEYINPUT95), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n617_), .A2(new_n618_), .A3(new_n584_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n599_), .ZN(new_n620_));
  AND4_X1   g419(.A1(new_n609_), .A2(new_n572_), .A3(new_n606_), .A4(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n609_), .B1(new_n600_), .B2(new_n606_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n515_), .B1(new_n619_), .B2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(KEYINPUT100), .ZN(new_n625_));
  INV_X1    g424(.A(new_n572_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n515_), .A2(new_n461_), .A3(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n614_), .A2(new_n625_), .A3(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n575_), .B1(new_n628_), .B2(new_n537_), .ZN(new_n629_));
  XOR2_X1   g428(.A(G113gat), .B(G141gat), .Z(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT78), .ZN(new_n631_));
  XNOR2_X1  g430(.A(G169gat), .B(G197gat), .ZN(new_n632_));
  XOR2_X1   g431(.A(new_n631_), .B(new_n632_), .Z(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT77), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n349_), .A2(new_n306_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(G229gat), .A2(G233gat), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT76), .ZN(new_n639_));
  INV_X1    g438(.A(new_n349_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n311_), .A2(new_n639_), .A3(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n640_), .A2(new_n308_), .A3(new_n310_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(KEYINPUT76), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n638_), .B1(new_n641_), .B2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n640_), .A2(new_n307_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(new_n636_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n648_), .A2(new_n637_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n635_), .B1(new_n645_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n635_), .ZN(new_n652_));
  NOR3_X1   g451(.A1(new_n644_), .A2(new_n649_), .A3(new_n652_), .ZN(new_n653_));
  OR2_X1    g452(.A1(new_n651_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  OAI21_X1  g454(.A(KEYINPUT102), .B1(new_n629_), .B2(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n627_), .B1(new_n624_), .B2(KEYINPUT100), .ZN(new_n657_));
  AOI211_X1 g456(.A(new_n613_), .B(new_n515_), .C1(new_n619_), .C2(new_n623_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n537_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(new_n574_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT102), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n660_), .A2(new_n661_), .A3(new_n654_), .ZN(new_n662_));
  AOI211_X1 g461(.A(new_n303_), .B(new_n364_), .C1(new_n656_), .C2(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n663_), .A2(new_n572_), .A3(new_n340_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n665_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n332_), .A2(new_n336_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n629_), .A2(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n302_), .A2(KEYINPUT104), .A3(new_n654_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n300_), .A2(new_n654_), .A3(new_n301_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT104), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n671_), .A2(new_n363_), .A3(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n670_), .A2(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(G1gat), .B1(new_n676_), .B2(new_n626_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n666_), .A2(new_n667_), .A3(new_n677_), .ZN(G1324gat));
  NAND3_X1  g477(.A1(new_n663_), .A2(new_n341_), .A3(new_n462_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT39), .ZN(new_n680_));
  OAI21_X1  g479(.A(G8gat), .B1(new_n680_), .B2(KEYINPUT105), .ZN(new_n681_));
  INV_X1    g480(.A(new_n676_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n681_), .B1(new_n682_), .B2(new_n462_), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n683_), .A2(KEYINPUT105), .A3(new_n680_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n683_), .B1(KEYINPUT105), .B2(new_n680_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n679_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT40), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  OAI211_X1 g487(.A(KEYINPUT40), .B(new_n679_), .C1(new_n684_), .C2(new_n685_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1325gat));
  OAI21_X1  g489(.A(G15gat), .B1(new_n676_), .B2(new_n537_), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT41), .Z(new_n692_));
  INV_X1    g491(.A(new_n537_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n663_), .A2(new_n529_), .A3(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n692_), .A2(new_n694_), .ZN(G1326gat));
  OAI21_X1  g494(.A(G22gat), .B1(new_n676_), .B2(new_n576_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT42), .ZN(new_n697_));
  INV_X1    g496(.A(G22gat), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n663_), .A2(new_n698_), .A3(new_n515_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n697_), .A2(new_n699_), .ZN(G1327gat));
  NOR2_X1   g499(.A1(new_n668_), .A2(new_n363_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n302_), .A2(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n702_), .B1(new_n656_), .B2(new_n662_), .ZN(new_n703_));
  AOI21_X1  g502(.A(G29gat), .B1(new_n703_), .B2(new_n572_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT108), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n671_), .A2(new_n362_), .A3(new_n674_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT106), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n706_), .B(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(KEYINPUT43), .B1(new_n629_), .B2(new_n339_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT43), .ZN(new_n710_));
  INV_X1    g509(.A(new_n339_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n660_), .A2(new_n710_), .A3(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n708_), .B1(new_n709_), .B2(new_n712_), .ZN(new_n713_));
  XOR2_X1   g512(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n714_));
  OAI21_X1  g513(.A(new_n705_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n708_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n710_), .B1(new_n660_), .B2(new_n711_), .ZN(new_n717_));
  AOI211_X1 g516(.A(KEYINPUT43), .B(new_n339_), .C1(new_n659_), .C2(new_n574_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n716_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n714_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n719_), .A2(KEYINPUT108), .A3(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n715_), .A2(new_n721_), .ZN(new_n722_));
  OAI211_X1 g521(.A(KEYINPUT44), .B(new_n716_), .C1(new_n717_), .C2(new_n718_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n572_), .A2(G29gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n704_), .B1(new_n725_), .B2(new_n726_), .ZN(G1328gat));
  INV_X1    g526(.A(KEYINPUT109), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT46), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(G36gat), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n723_), .A2(new_n462_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n731_), .B1(new_n722_), .B2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n702_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n461_), .A2(G36gat), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n629_), .A2(KEYINPUT102), .A3(new_n655_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n661_), .B1(new_n660_), .B2(new_n654_), .ZN(new_n738_));
  OAI211_X1 g537(.A(new_n735_), .B(new_n736_), .C1(new_n737_), .C2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(KEYINPUT45), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT45), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n703_), .A2(new_n741_), .A3(new_n736_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n728_), .A2(new_n729_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n730_), .B1(new_n734_), .B2(new_n745_), .ZN(new_n746_));
  AOI22_X1  g545(.A1(new_n740_), .A2(new_n742_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n730_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n732_), .B1(new_n715_), .B2(new_n721_), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n747_), .B(new_n748_), .C1(new_n749_), .C2(new_n731_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n746_), .A2(new_n750_), .ZN(G1329gat));
  INV_X1    g550(.A(KEYINPUT47), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n703_), .A2(new_n693_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n693_), .A2(G43gat), .ZN(new_n754_));
  OAI221_X1 g553(.A(new_n752_), .B1(G43gat), .B2(new_n753_), .C1(new_n724_), .C2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n723_), .ZN(new_n756_));
  AOI211_X1 g555(.A(new_n754_), .B(new_n756_), .C1(new_n715_), .C2(new_n721_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n753_), .A2(G43gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(KEYINPUT47), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n755_), .A2(new_n759_), .ZN(G1330gat));
  AOI21_X1  g559(.A(G50gat), .B1(new_n703_), .B2(new_n515_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n515_), .A2(G50gat), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n725_), .B2(new_n762_), .ZN(G1331gat));
  NAND2_X1  g562(.A1(new_n363_), .A2(new_n655_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n302_), .A2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n670_), .A2(new_n765_), .ZN(new_n766_));
  OAI21_X1  g565(.A(G57gat), .B1(new_n766_), .B2(new_n626_), .ZN(new_n767_));
  NOR4_X1   g566(.A1(new_n629_), .A2(new_n654_), .A3(new_n302_), .A4(new_n364_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n768_), .A2(new_n207_), .A3(new_n572_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(G1332gat));
  NAND3_X1  g569(.A1(new_n768_), .A2(new_n209_), .A3(new_n462_), .ZN(new_n771_));
  OAI21_X1  g570(.A(G64gat), .B1(new_n766_), .B2(new_n461_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n772_), .A2(KEYINPUT48), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n772_), .A2(KEYINPUT48), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n771_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  XOR2_X1   g574(.A(new_n775_), .B(KEYINPUT110), .Z(G1333gat));
  OAI21_X1  g575(.A(G71gat), .B1(new_n766_), .B2(new_n537_), .ZN(new_n777_));
  XOR2_X1   g576(.A(KEYINPUT111), .B(KEYINPUT49), .Z(new_n778_));
  XNOR2_X1  g577(.A(new_n777_), .B(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(G71gat), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n768_), .A2(new_n780_), .A3(new_n693_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n781_), .ZN(G1334gat));
  OAI21_X1  g581(.A(G78gat), .B1(new_n766_), .B2(new_n576_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT50), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n768_), .A2(new_n499_), .A3(new_n515_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(G1335gat));
  NOR2_X1   g585(.A1(new_n629_), .A2(new_n654_), .ZN(new_n787_));
  NOR3_X1   g586(.A1(new_n302_), .A2(new_n363_), .A3(new_n668_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(G85gat), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n790_), .A2(new_n791_), .A3(new_n572_), .ZN(new_n792_));
  NOR3_X1   g591(.A1(new_n302_), .A2(new_n654_), .A3(new_n363_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n794_), .B1(new_n709_), .B2(new_n712_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n795_), .A2(new_n572_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n792_), .B1(new_n796_), .B2(new_n791_), .ZN(G1336gat));
  INV_X1    g596(.A(G92gat), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n790_), .A2(new_n798_), .A3(new_n462_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n795_), .A2(new_n462_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n799_), .B1(new_n800_), .B2(new_n798_), .ZN(G1337gat));
  NOR3_X1   g600(.A1(new_n789_), .A2(new_n537_), .A3(new_n265_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n795_), .A2(new_n693_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n802_), .B1(new_n803_), .B2(G99gat), .ZN(new_n804_));
  XOR2_X1   g603(.A(new_n804_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g604(.A1(new_n790_), .A2(new_n267_), .A3(new_n515_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n795_), .A2(new_n515_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n807_), .B1(new_n808_), .B2(G106gat), .ZN(new_n809_));
  AOI211_X1 g608(.A(KEYINPUT52), .B(new_n267_), .C1(new_n795_), .C2(new_n515_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n806_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n811_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g611(.A(KEYINPUT112), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n764_), .B(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n814_), .A2(new_n302_), .A3(new_n339_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(KEYINPUT54), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT54), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n814_), .A2(new_n817_), .A3(new_n339_), .A4(new_n302_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n654_), .A2(new_n297_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT56), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n295_), .A2(KEYINPUT55), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n292_), .A2(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n289_), .A2(new_n286_), .A3(new_n291_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT113), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT113), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n289_), .A2(new_n827_), .A3(new_n286_), .A4(new_n291_), .ZN(new_n828_));
  AOI22_X1  g627(.A1(new_n822_), .A2(new_n824_), .B1(new_n826_), .B2(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n821_), .B1(new_n829_), .B2(new_n296_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n826_), .A2(new_n828_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n292_), .A2(new_n823_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n292_), .A2(new_n823_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n831_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n296_), .A2(new_n821_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n820_), .B1(new_n830_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n637_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n636_), .A2(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n839_), .B1(new_n641_), .B2(new_n643_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n648_), .A2(new_n838_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n634_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n633_), .B1(new_n644_), .B2(new_n649_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n298_), .A2(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n668_), .B1(new_n837_), .B2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT57), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  OAI211_X1 g647(.A(KEYINPUT57), .B(new_n668_), .C1(new_n837_), .C2(new_n845_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT115), .ZN(new_n851_));
  INV_X1    g650(.A(new_n835_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n851_), .B1(new_n829_), .B2(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n834_), .A2(KEYINPUT115), .A3(new_n835_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n830_), .A2(new_n853_), .A3(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n844_), .A2(new_n297_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(KEYINPUT114), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT114), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n844_), .A2(new_n297_), .A3(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n855_), .A2(KEYINPUT58), .A3(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT116), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n855_), .A2(KEYINPUT116), .A3(KEYINPUT58), .A4(new_n860_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(KEYINPUT58), .B1(new_n855_), .B2(new_n860_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n866_), .A2(new_n339_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n850_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n819_), .B1(new_n868_), .B2(new_n363_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n626_), .A2(new_n537_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n516_), .A2(new_n870_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n871_), .A2(KEYINPUT59), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n869_), .A2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n654_), .A2(G113gat), .ZN(new_n874_));
  XOR2_X1   g673(.A(new_n874_), .B(KEYINPUT119), .Z(new_n875_));
  INV_X1    g674(.A(KEYINPUT118), .ZN(new_n876_));
  INV_X1    g675(.A(new_n819_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n865_), .A2(new_n867_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(KEYINPUT117), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT117), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n865_), .A2(new_n867_), .A3(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n850_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n879_), .A2(new_n881_), .A3(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n877_), .B1(new_n883_), .B2(new_n362_), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n876_), .B(KEYINPUT59), .C1(new_n884_), .C2(new_n871_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n871_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n850_), .B1(new_n878_), .B2(KEYINPUT117), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n363_), .B1(new_n888_), .B2(new_n881_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n887_), .B1(new_n889_), .B2(new_n877_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n876_), .B1(new_n890_), .B2(KEYINPUT59), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n873_), .B(new_n875_), .C1(new_n886_), .C2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(G113gat), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n893_), .B1(new_n890_), .B2(new_n655_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(KEYINPUT120), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT120), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n892_), .A2(new_n897_), .A3(new_n894_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n896_), .A2(new_n898_), .ZN(G1340gat));
  OAI21_X1  g698(.A(new_n873_), .B1(new_n886_), .B2(new_n891_), .ZN(new_n900_));
  OAI21_X1  g699(.A(G120gat), .B1(new_n900_), .B2(new_n302_), .ZN(new_n901_));
  INV_X1    g700(.A(G120gat), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n902_), .B1(new_n302_), .B2(KEYINPUT60), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n903_), .B1(KEYINPUT60), .B2(new_n902_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n901_), .B1(new_n890_), .B2(new_n904_), .ZN(G1341gat));
  INV_X1    g704(.A(new_n890_), .ZN(new_n906_));
  AOI21_X1  g705(.A(G127gat), .B1(new_n906_), .B2(new_n363_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n900_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n362_), .A2(KEYINPUT121), .ZN(new_n909_));
  MUX2_X1   g708(.A(KEYINPUT121), .B(new_n909_), .S(G127gat), .Z(new_n910_));
  AOI21_X1  g709(.A(new_n907_), .B1(new_n908_), .B2(new_n910_), .ZN(G1342gat));
  OAI21_X1  g710(.A(G134gat), .B1(new_n900_), .B2(new_n339_), .ZN(new_n912_));
  OR2_X1    g711(.A1(new_n668_), .A2(G134gat), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n890_), .B2(new_n913_), .ZN(G1343gat));
  NAND4_X1  g713(.A1(new_n515_), .A2(new_n461_), .A3(new_n572_), .A4(new_n537_), .ZN(new_n915_));
  OAI21_X1  g714(.A(KEYINPUT122), .B1(new_n884_), .B2(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT122), .ZN(new_n917_));
  INV_X1    g716(.A(new_n915_), .ZN(new_n918_));
  OAI211_X1 g717(.A(new_n917_), .B(new_n918_), .C1(new_n889_), .C2(new_n877_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n916_), .A2(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(new_n654_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g721(.A1(new_n920_), .A2(new_n303_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(G148gat), .ZN(G1345gat));
  AND3_X1   g723(.A1(new_n865_), .A2(new_n867_), .A3(new_n880_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n880_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n926_));
  NOR3_X1   g725(.A1(new_n925_), .A2(new_n926_), .A3(new_n850_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n819_), .B1(new_n927_), .B2(new_n363_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n917_), .B1(new_n928_), .B2(new_n918_), .ZN(new_n929_));
  NOR3_X1   g728(.A1(new_n884_), .A2(KEYINPUT122), .A3(new_n915_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n363_), .B1(new_n929_), .B2(new_n930_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n931_), .A2(KEYINPUT123), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT123), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n920_), .A2(new_n933_), .A3(new_n363_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(KEYINPUT61), .B(G155gat), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n932_), .A2(new_n934_), .A3(new_n935_), .ZN(new_n936_));
  INV_X1    g735(.A(new_n935_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n933_), .B1(new_n920_), .B2(new_n363_), .ZN(new_n938_));
  AOI211_X1 g737(.A(KEYINPUT123), .B(new_n362_), .C1(new_n916_), .C2(new_n919_), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n937_), .B1(new_n938_), .B2(new_n939_), .ZN(new_n940_));
  AND2_X1   g739(.A1(new_n936_), .A2(new_n940_), .ZN(G1346gat));
  INV_X1    g740(.A(new_n920_), .ZN(new_n942_));
  OR3_X1    g741(.A1(new_n942_), .A2(G162gat), .A3(new_n668_), .ZN(new_n943_));
  OAI21_X1  g742(.A(G162gat), .B1(new_n942_), .B2(new_n339_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n943_), .A2(new_n944_), .ZN(G1347gat));
  NAND2_X1  g744(.A1(new_n462_), .A2(new_n573_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n946_), .A2(new_n515_), .ZN(new_n947_));
  AND2_X1   g746(.A1(new_n869_), .A2(new_n947_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n948_), .A2(new_n654_), .ZN(new_n949_));
  INV_X1    g748(.A(KEYINPUT124), .ZN(new_n950_));
  NOR2_X1   g749(.A1(new_n950_), .A2(KEYINPUT62), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n376_), .B1(new_n950_), .B2(KEYINPUT62), .ZN(new_n952_));
  AND3_X1   g751(.A1(new_n949_), .A2(new_n951_), .A3(new_n952_), .ZN(new_n953_));
  AOI21_X1  g752(.A(new_n951_), .B1(new_n949_), .B2(new_n952_), .ZN(new_n954_));
  XOR2_X1   g753(.A(KEYINPUT22), .B(G169gat), .Z(new_n955_));
  OAI22_X1  g754(.A1(new_n953_), .A2(new_n954_), .B1(new_n949_), .B2(new_n955_), .ZN(G1348gat));
  AOI21_X1  g755(.A(G176gat), .B1(new_n948_), .B2(new_n303_), .ZN(new_n957_));
  NOR2_X1   g756(.A1(new_n884_), .A2(new_n515_), .ZN(new_n958_));
  INV_X1    g757(.A(new_n946_), .ZN(new_n959_));
  NAND3_X1  g758(.A1(new_n303_), .A2(new_n959_), .A3(G176gat), .ZN(new_n960_));
  INV_X1    g759(.A(new_n960_), .ZN(new_n961_));
  AOI21_X1  g760(.A(new_n957_), .B1(new_n958_), .B2(new_n961_), .ZN(G1349gat));
  NAND3_X1  g761(.A1(new_n958_), .A2(new_n363_), .A3(new_n959_), .ZN(new_n963_));
  NOR2_X1   g762(.A1(new_n362_), .A2(new_n367_), .ZN(new_n964_));
  AOI22_X1  g763(.A1(new_n963_), .A2(new_n399_), .B1(new_n948_), .B2(new_n964_), .ZN(G1350gat));
  NAND3_X1  g764(.A1(new_n948_), .A2(new_n368_), .A3(new_n669_), .ZN(new_n966_));
  INV_X1    g765(.A(new_n948_), .ZN(new_n967_));
  OAI21_X1  g766(.A(G190gat), .B1(new_n967_), .B2(new_n339_), .ZN(new_n968_));
  INV_X1    g767(.A(KEYINPUT125), .ZN(new_n969_));
  AND2_X1   g768(.A1(new_n968_), .A2(new_n969_), .ZN(new_n970_));
  NOR2_X1   g769(.A1(new_n968_), .A2(new_n969_), .ZN(new_n971_));
  OAI21_X1  g770(.A(new_n966_), .B1(new_n970_), .B2(new_n971_), .ZN(G1351gat));
  NAND4_X1  g771(.A1(new_n462_), .A2(new_n515_), .A3(new_n626_), .A4(new_n537_), .ZN(new_n973_));
  NOR2_X1   g772(.A1(new_n884_), .A2(new_n973_), .ZN(new_n974_));
  INV_X1    g773(.A(KEYINPUT126), .ZN(new_n975_));
  XNOR2_X1  g774(.A(new_n974_), .B(new_n975_), .ZN(new_n976_));
  AND3_X1   g775(.A1(new_n976_), .A2(G197gat), .A3(new_n654_), .ZN(new_n977_));
  AOI21_X1  g776(.A(G197gat), .B1(new_n976_), .B2(new_n654_), .ZN(new_n978_));
  NOR2_X1   g777(.A1(new_n977_), .A2(new_n978_), .ZN(G1352gat));
  XNOR2_X1  g778(.A(new_n974_), .B(KEYINPUT126), .ZN(new_n980_));
  OAI211_X1 g779(.A(KEYINPUT127), .B(G204gat), .C1(new_n980_), .C2(new_n302_), .ZN(new_n981_));
  NAND2_X1  g780(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n982_));
  NAND3_X1  g781(.A1(new_n976_), .A2(new_n303_), .A3(new_n982_), .ZN(new_n983_));
  NAND2_X1  g782(.A1(new_n981_), .A2(new_n983_), .ZN(G1353gat));
  XNOR2_X1  g783(.A(KEYINPUT63), .B(G211gat), .ZN(new_n985_));
  NOR3_X1   g784(.A1(new_n980_), .A2(new_n362_), .A3(new_n985_), .ZN(new_n986_));
  NAND2_X1  g785(.A1(new_n976_), .A2(new_n363_), .ZN(new_n987_));
  NOR2_X1   g786(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n988_));
  AOI21_X1  g787(.A(new_n986_), .B1(new_n987_), .B2(new_n988_), .ZN(G1354gat));
  OR3_X1    g788(.A1(new_n980_), .A2(G218gat), .A3(new_n668_), .ZN(new_n990_));
  OAI21_X1  g789(.A(G218gat), .B1(new_n980_), .B2(new_n339_), .ZN(new_n991_));
  NAND2_X1  g790(.A1(new_n990_), .A2(new_n991_), .ZN(G1355gat));
endmodule


