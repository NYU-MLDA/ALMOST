//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 0 0 0 0 1 1 1 0 0 0 1 0 0 1 1 1 1 0 0 1 0 0 1 1 0 1 0 0 0 1 0 0 0 0 1 0 1 1 0 0 1 0 0 0 1 0 1 0 1 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n685_, new_n686_, new_n687_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n838_, new_n839_, new_n840_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n851_,
    new_n852_, new_n854_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n871_, new_n873_, new_n875_, new_n876_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n883_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_;
  NOR2_X1   g000(.A1(KEYINPUT70), .A2(KEYINPUT13), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G230gat), .A2(G233gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(G85gat), .B(G92gat), .Z(new_n205_));
  XOR2_X1   g004(.A(KEYINPUT65), .B(KEYINPUT8), .Z(new_n206_));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT6), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT6), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n209_), .A2(G99gat), .A3(G106gat), .ZN(new_n210_));
  AND2_X1   g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT7), .ZN(new_n212_));
  INV_X1    g011(.A(G99gat), .ZN(new_n213_));
  INV_X1    g012(.A(G106gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n212_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n205_), .B(new_n206_), .C1(new_n211_), .C2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT66), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n205_), .B1(new_n211_), .B2(new_n217_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT8), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n208_), .A2(new_n210_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n222_), .A2(new_n216_), .A3(new_n215_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n223_), .A2(new_n224_), .A3(new_n205_), .A4(new_n206_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n219_), .A2(new_n221_), .A3(new_n225_), .ZN(new_n226_));
  XOR2_X1   g025(.A(KEYINPUT10), .B(G99gat), .Z(new_n227_));
  AOI21_X1  g026(.A(new_n211_), .B1(new_n214_), .B2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n205_), .A2(KEYINPUT9), .ZN(new_n229_));
  XOR2_X1   g028(.A(KEYINPUT64), .B(G92gat), .Z(new_n230_));
  INV_X1    g029(.A(KEYINPUT9), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n230_), .A2(new_n231_), .A3(G85gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n228_), .A2(new_n229_), .A3(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(G71gat), .B(G78gat), .Z(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G57gat), .B(G64gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT11), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n235_), .A2(new_n237_), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n236_), .A2(KEYINPUT11), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n234_), .A2(KEYINPUT11), .A3(new_n236_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n238_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  AND3_X1   g041(.A1(new_n226_), .A2(new_n233_), .A3(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n242_), .B1(new_n226_), .B2(new_n233_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT12), .ZN(new_n245_));
  NOR3_X1   g044(.A1(new_n243_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n245_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n204_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n226_), .A2(new_n233_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(new_n241_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n226_), .A2(new_n233_), .A3(new_n242_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n204_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G120gat), .B(G148gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT5), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(G176gat), .ZN(new_n257_));
  INV_X1    g056(.A(G204gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n249_), .A2(new_n254_), .A3(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT68), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n251_), .A2(KEYINPUT12), .A3(new_n252_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(new_n247_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n253_), .B1(new_n265_), .B2(new_n204_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n266_), .A2(KEYINPUT68), .A3(new_n260_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n263_), .A2(new_n267_), .ZN(new_n268_));
  OAI21_X1  g067(.A(KEYINPUT67), .B1(new_n266_), .B2(new_n260_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT67), .ZN(new_n270_));
  INV_X1    g069(.A(new_n204_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n271_), .B1(new_n264_), .B2(new_n247_), .ZN(new_n272_));
  OAI211_X1 g071(.A(new_n270_), .B(new_n259_), .C1(new_n272_), .C2(new_n253_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n269_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT69), .ZN(new_n275_));
  AND3_X1   g074(.A1(new_n268_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n275_), .B1(new_n268_), .B2(new_n274_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n203_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n249_), .A2(new_n254_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n270_), .B1(new_n279_), .B2(new_n259_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n273_), .ZN(new_n281_));
  AOI21_X1  g080(.A(KEYINPUT68), .B1(new_n266_), .B2(new_n260_), .ZN(new_n282_));
  NOR4_X1   g081(.A1(new_n272_), .A2(new_n262_), .A3(new_n253_), .A4(new_n259_), .ZN(new_n283_));
  OAI22_X1  g082(.A1(new_n280_), .A2(new_n281_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT69), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n268_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n286_));
  XOR2_X1   g085(.A(KEYINPUT70), .B(KEYINPUT13), .Z(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n285_), .A2(new_n286_), .A3(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n278_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G229gat), .A2(G233gat), .ZN(new_n291_));
  INV_X1    g090(.A(G8gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT73), .B(G1gat), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT14), .B1(new_n293_), .B2(new_n292_), .ZN(new_n294_));
  INV_X1    g093(.A(G1gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G15gat), .B(G22gat), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n294_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n295_), .B1(new_n294_), .B2(new_n296_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n292_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n299_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n301_), .A2(G8gat), .A3(new_n297_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G29gat), .B(G36gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(G43gat), .ZN(new_n306_));
  INV_X1    g105(.A(G50gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  OR2_X1    g107(.A1(new_n305_), .A2(G43gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n305_), .A2(G43gat), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n309_), .A2(G50gat), .A3(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n308_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT15), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n308_), .A2(KEYINPUT15), .A3(new_n311_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n304_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n312_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n303_), .A2(KEYINPUT79), .A3(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(KEYINPUT79), .B1(new_n303_), .B2(new_n318_), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n291_), .B(new_n317_), .C1(new_n320_), .C2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n321_), .ZN(new_n323_));
  AOI22_X1  g122(.A1(new_n323_), .A2(new_n319_), .B1(new_n304_), .B2(new_n312_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n322_), .B1(new_n324_), .B2(new_n291_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G113gat), .B(G141gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT80), .ZN(new_n327_));
  INV_X1    g126(.A(G169gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(G197gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n325_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n331_), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n322_), .B(new_n333_), .C1(new_n324_), .C2(new_n291_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n290_), .A2(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT102), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G15gat), .B(G43gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT31), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G183gat), .A2(G190gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT23), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n342_), .B1(G183gat), .B2(G190gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G169gat), .A2(G176gat), .ZN(new_n344_));
  AND2_X1   g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT22), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT84), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n346_), .B1(new_n347_), .B2(new_n328_), .ZN(new_n348_));
  NAND4_X1  g147(.A1(KEYINPUT83), .A2(KEYINPUT84), .A3(KEYINPUT22), .A4(G169gat), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n348_), .B(new_n349_), .C1(KEYINPUT83), .C2(G169gat), .ZN(new_n350_));
  INV_X1    g149(.A(G176gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n345_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n328_), .A2(new_n351_), .ZN(new_n354_));
  OR2_X1    g153(.A1(new_n354_), .A2(KEYINPUT24), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n342_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT82), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n354_), .A2(KEYINPUT24), .A3(new_n344_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n342_), .A2(new_n355_), .A3(KEYINPUT82), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT25), .ZN(new_n361_));
  OAI21_X1  g160(.A(KEYINPUT81), .B1(new_n361_), .B2(G183gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT26), .B(G190gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(KEYINPUT25), .B(G183gat), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n362_), .B(new_n363_), .C1(new_n364_), .C2(KEYINPUT81), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n358_), .A2(new_n359_), .A3(new_n360_), .A4(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n353_), .A2(new_n366_), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n367_), .A2(KEYINPUT30), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n367_), .A2(KEYINPUT30), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  XOR2_X1   g169(.A(G71gat), .B(G99gat), .Z(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n371_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n373_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n340_), .B1(new_n372_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT86), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G127gat), .B(G134gat), .ZN(new_n378_));
  OR2_X1    g177(.A1(new_n378_), .A2(KEYINPUT85), .ZN(new_n379_));
  INV_X1    g178(.A(G113gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(KEYINPUT85), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n379_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n380_), .B1(new_n379_), .B2(new_n381_), .ZN(new_n384_));
  INV_X1    g183(.A(G120gat), .ZN(new_n385_));
  NOR3_X1   g184(.A1(new_n383_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n379_), .A2(new_n381_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(G113gat), .ZN(new_n388_));
  AOI21_X1  g187(.A(G120gat), .B1(new_n388_), .B2(new_n382_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n377_), .B1(new_n386_), .B2(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n385_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n388_), .A2(new_n382_), .A3(G120gat), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n391_), .A2(new_n392_), .A3(KEYINPUT86), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n390_), .A2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n394_), .A2(G227gat), .A3(G233gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G227gat), .A2(G233gat), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n390_), .A2(new_n393_), .A3(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n372_), .A2(new_n374_), .A3(new_n340_), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n376_), .A2(new_n395_), .A3(new_n397_), .A4(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n395_), .A2(new_n397_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n398_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n400_), .B1(new_n401_), .B2(new_n375_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n399_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G78gat), .B(G106gat), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(G141gat), .A2(G148gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G155gat), .A2(G162gat), .ZN(new_n408_));
  XOR2_X1   g207(.A(new_n408_), .B(KEYINPUT1), .Z(new_n409_));
  NOR2_X1   g208(.A1(G155gat), .A2(G162gat), .ZN(new_n410_));
  XOR2_X1   g209(.A(new_n410_), .B(KEYINPUT87), .Z(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n407_), .B1(new_n409_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G141gat), .A2(G148gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  AND2_X1   g214(.A1(KEYINPUT88), .A2(KEYINPUT2), .ZN(new_n416_));
  NOR2_X1   g215(.A1(KEYINPUT88), .A2(KEYINPUT2), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n414_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT89), .ZN(new_n419_));
  INV_X1    g218(.A(new_n414_), .ZN(new_n420_));
  AOI22_X1  g219(.A1(new_n418_), .A2(new_n419_), .B1(KEYINPUT2), .B2(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n407_), .B(KEYINPUT3), .ZN(new_n422_));
  OAI211_X1 g221(.A(new_n421_), .B(new_n422_), .C1(new_n419_), .C2(new_n418_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n411_), .B1(G155gat), .B2(G162gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n415_), .A2(new_n425_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n426_), .A2(KEYINPUT29), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n258_), .A2(G197gat), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n330_), .A2(G204gat), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT21), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  XOR2_X1   g229(.A(G211gat), .B(G218gat), .Z(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  OR3_X1    g231(.A1(new_n258_), .A2(KEYINPUT90), .A3(G197gat), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n429_), .A2(KEYINPUT90), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n433_), .B1(new_n434_), .B2(new_n428_), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n430_), .B(new_n432_), .C1(new_n435_), .C2(KEYINPUT21), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n435_), .A2(KEYINPUT21), .A3(new_n431_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  OR3_X1    g238(.A1(new_n427_), .A2(G50gat), .A3(new_n439_), .ZN(new_n440_));
  OAI21_X1  g239(.A(G50gat), .B1(new_n427_), .B2(new_n439_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n406_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n426_), .A2(KEYINPUT29), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT28), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NOR3_X1   g245(.A1(new_n426_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G228gat), .A2(G233gat), .ZN(new_n448_));
  INV_X1    g247(.A(G22gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  OR3_X1    g249(.A1(new_n446_), .A2(new_n447_), .A3(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n450_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n440_), .A2(new_n441_), .A3(new_n406_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n443_), .A2(new_n451_), .A3(new_n452_), .A4(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n451_), .A2(new_n452_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n453_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n455_), .B1(new_n456_), .B2(new_n442_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n454_), .A2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n390_), .A2(new_n393_), .A3(new_n426_), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n415_), .A2(new_n391_), .A3(new_n392_), .A4(new_n425_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G225gat), .A2(G233gat), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n461_), .A2(new_n463_), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n390_), .A2(KEYINPUT96), .A3(new_n393_), .A4(new_n426_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n461_), .A2(KEYINPUT4), .A3(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT4), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n467_), .B1(new_n459_), .B2(KEYINPUT96), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n464_), .B1(new_n469_), .B2(new_n463_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G1gat), .B(G29gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(G85gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n472_), .B(KEYINPUT0), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(G57gat), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n470_), .A2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n462_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n474_), .B1(new_n477_), .B2(new_n464_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n476_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G226gat), .A2(G233gat), .ZN(new_n480_));
  XOR2_X1   g279(.A(new_n480_), .B(KEYINPUT91), .Z(new_n481_));
  XOR2_X1   g280(.A(new_n481_), .B(KEYINPUT19), .Z(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT22), .B(G169gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(new_n351_), .ZN(new_n485_));
  AND3_X1   g284(.A1(new_n343_), .A2(new_n344_), .A3(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n356_), .A2(KEYINPUT94), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT94), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n342_), .A2(new_n355_), .A3(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n344_), .A2(KEYINPUT24), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n490_), .B(KEYINPUT93), .Z(new_n491_));
  AOI22_X1  g290(.A1(new_n487_), .A2(new_n489_), .B1(new_n491_), .B2(new_n354_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n364_), .B(KEYINPUT92), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(new_n363_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n486_), .B1(new_n492_), .B2(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n483_), .B1(new_n495_), .B2(new_n439_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n367_), .A2(new_n438_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n496_), .A2(KEYINPUT20), .A3(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n439_), .A2(new_n353_), .A3(new_n366_), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n499_), .B(KEYINPUT20), .C1(new_n439_), .C2(new_n495_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(new_n483_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n501_), .A2(KEYINPUT95), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT95), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n503_), .B1(new_n500_), .B2(new_n483_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n498_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G8gat), .B(G36gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT18), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(G64gat), .ZN(new_n508_));
  INV_X1    g307(.A(G92gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT32), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  OR2_X1    g311(.A1(new_n505_), .A2(new_n512_), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n495_), .A2(KEYINPUT98), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n495_), .A2(KEYINPUT98), .ZN(new_n515_));
  NOR3_X1   g314(.A1(new_n514_), .A2(new_n515_), .A3(new_n438_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n497_), .A2(KEYINPUT20), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n483_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT99), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  OAI211_X1 g319(.A(KEYINPUT99), .B(new_n483_), .C1(new_n516_), .C2(new_n517_), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n520_), .B(new_n521_), .C1(new_n483_), .C2(new_n500_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(new_n512_), .ZN(new_n523_));
  AND3_X1   g322(.A1(new_n479_), .A2(new_n513_), .A3(new_n523_), .ZN(new_n524_));
  OAI211_X1 g323(.A(new_n498_), .B(new_n510_), .C1(new_n502_), .C2(new_n504_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n510_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n505_), .A2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n459_), .A2(new_n463_), .A3(new_n460_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(new_n474_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT97), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n463_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n525_), .B(new_n527_), .C1(new_n531_), .C2(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(KEYINPUT33), .B1(new_n470_), .B2(new_n475_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT33), .ZN(new_n535_));
  NOR4_X1   g334(.A1(new_n477_), .A2(new_n535_), .A3(new_n464_), .A4(new_n474_), .ZN(new_n536_));
  NOR3_X1   g335(.A1(new_n533_), .A2(new_n534_), .A3(new_n536_), .ZN(new_n537_));
  OAI211_X1 g336(.A(new_n404_), .B(new_n458_), .C1(new_n524_), .C2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n458_), .A2(new_n403_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n454_), .A2(new_n457_), .A3(new_n402_), .A4(new_n399_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(KEYINPUT27), .B1(new_n527_), .B2(new_n525_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n525_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n543_), .B1(new_n522_), .B2(new_n526_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n542_), .B1(new_n544_), .B2(KEYINPUT27), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT100), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n479_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n476_), .A2(KEYINPUT100), .A3(new_n478_), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n541_), .A2(new_n545_), .A3(new_n547_), .A4(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n538_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n316_), .A2(new_n250_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n551_), .B1(new_n312_), .B2(new_n250_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G232gat), .A2(G233gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT34), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n551_), .A2(KEYINPUT71), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n553_), .A2(KEYINPUT35), .A3(new_n555_), .A4(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n556_), .A2(KEYINPUT35), .A3(new_n555_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(new_n552_), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n555_), .A2(KEYINPUT35), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n557_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G190gat), .B(G218gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(G134gat), .ZN(new_n563_));
  INV_X1    g362(.A(G162gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n566_), .A2(KEYINPUT36), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n566_), .A2(KEYINPUT36), .ZN(new_n568_));
  OR3_X1    g367(.A1(new_n561_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n561_), .A2(KEYINPUT72), .A3(new_n567_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(KEYINPUT72), .B1(new_n561_), .B2(new_n567_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n569_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G231gat), .A2(G233gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT74), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n304_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n304_), .A2(new_n576_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(new_n241_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n577_), .A2(new_n242_), .A3(new_n578_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G127gat), .B(G155gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G183gat), .B(G211gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n586_), .B(KEYINPUT17), .Z(new_n587_));
  NAND3_X1  g386(.A1(new_n580_), .A2(new_n581_), .A3(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT77), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n580_), .A2(new_n581_), .A3(KEYINPUT77), .A4(new_n587_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n580_), .A2(new_n581_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n586_), .A2(KEYINPUT17), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n594_), .B(KEYINPUT76), .Z(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n592_), .B1(new_n593_), .B2(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n574_), .A2(new_n597_), .ZN(new_n598_));
  AND3_X1   g397(.A1(new_n337_), .A2(new_n550_), .A3(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n547_), .A2(new_n548_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(G1gat), .B1(new_n600_), .B2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT38), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n573_), .A2(KEYINPUT37), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT37), .ZN(new_n606_));
  OAI211_X1 g405(.A(new_n569_), .B(new_n606_), .C1(new_n571_), .C2(new_n572_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n597_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT78), .ZN(new_n611_));
  INV_X1    g410(.A(new_n336_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n550_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n611_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n602_), .A2(KEYINPUT101), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n602_), .A2(KEYINPUT101), .ZN(new_n618_));
  OAI211_X1 g417(.A(new_n616_), .B(new_n293_), .C1(new_n617_), .C2(new_n618_), .ZN(new_n619_));
  AND3_X1   g418(.A1(new_n619_), .A2(KEYINPUT103), .A3(new_n604_), .ZN(new_n620_));
  AOI21_X1  g419(.A(KEYINPUT103), .B1(new_n619_), .B2(new_n604_), .ZN(new_n621_));
  OAI221_X1 g420(.A(new_n603_), .B1(new_n604_), .B2(new_n619_), .C1(new_n620_), .C2(new_n621_), .ZN(G1324gat));
  INV_X1    g421(.A(new_n545_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n292_), .B1(new_n599_), .B2(new_n623_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n624_), .B(KEYINPUT39), .Z(new_n625_));
  NAND3_X1  g424(.A1(new_n616_), .A2(new_n292_), .A3(new_n623_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  XOR2_X1   g426(.A(new_n627_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g427(.A(G15gat), .B1(new_n600_), .B2(new_n404_), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n629_), .B(KEYINPUT41), .Z(new_n630_));
  NOR3_X1   g429(.A1(new_n615_), .A2(G15gat), .A3(new_n404_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT104), .Z(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(G1326gat));
  INV_X1    g432(.A(new_n458_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n449_), .B1(new_n599_), .B2(new_n634_), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n635_), .B(KEYINPUT42), .Z(new_n636_));
  NAND3_X1  g435(.A1(new_n616_), .A2(new_n449_), .A3(new_n634_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(G1327gat));
  INV_X1    g437(.A(KEYINPUT108), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n608_), .B1(new_n538_), .B2(new_n549_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT43), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n640_), .A2(KEYINPUT106), .A3(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(KEYINPUT106), .B1(new_n640_), .B2(new_n641_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n640_), .A2(new_n641_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n612_), .A2(KEYINPUT102), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT102), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n336_), .A2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n646_), .A2(new_n597_), .A3(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(KEYINPUT105), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT105), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n337_), .A2(new_n651_), .A3(new_n597_), .ZN(new_n652_));
  AOI22_X1  g451(.A1(new_n644_), .A2(new_n645_), .B1(new_n650_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT107), .ZN(new_n654_));
  OAI211_X1 g453(.A(new_n639_), .B(KEYINPUT44), .C1(new_n653_), .C2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n650_), .A2(new_n652_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n640_), .A2(new_n641_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT106), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n640_), .A2(KEYINPUT106), .A3(new_n641_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n659_), .A2(new_n645_), .A3(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n656_), .A2(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(KEYINPUT108), .B1(new_n662_), .B2(KEYINPUT107), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT44), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n664_), .B1(new_n662_), .B2(KEYINPUT108), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n655_), .B1(new_n663_), .B2(new_n665_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n618_), .A2(new_n617_), .ZN(new_n667_));
  OAI21_X1  g466(.A(G29gat), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n574_), .A2(new_n597_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n613_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n602_), .A2(G29gat), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n668_), .B1(new_n671_), .B2(new_n672_), .ZN(G1328gat));
  OAI211_X1 g472(.A(new_n655_), .B(new_n623_), .C1(new_n663_), .C2(new_n665_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(G36gat), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n671_), .A2(G36gat), .A3(new_n545_), .ZN(new_n676_));
  XOR2_X1   g475(.A(KEYINPUT109), .B(KEYINPUT110), .Z(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT45), .ZN(new_n678_));
  XOR2_X1   g477(.A(new_n676_), .B(new_n678_), .Z(new_n679_));
  NAND2_X1  g478(.A1(new_n675_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT46), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n675_), .A2(KEYINPUT46), .A3(new_n679_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(G1329gat));
  NOR3_X1   g483(.A1(new_n671_), .A2(G43gat), .A3(new_n404_), .ZN(new_n685_));
  OAI211_X1 g484(.A(new_n655_), .B(new_n403_), .C1(new_n663_), .C2(new_n665_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n685_), .B1(new_n686_), .B2(G43gat), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g487(.A(G50gat), .B1(new_n666_), .B2(new_n458_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n670_), .A2(new_n307_), .A3(new_n634_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(G1331gat));
  NOR2_X1   g490(.A1(new_n290_), .A2(new_n335_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n550_), .A2(new_n692_), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n693_), .A2(new_n574_), .A3(new_n597_), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n694_), .A2(KEYINPUT111), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(KEYINPUT111), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n695_), .A2(G57gat), .A3(new_n601_), .A4(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(G57gat), .ZN(new_n698_));
  INV_X1    g497(.A(new_n693_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n611_), .A2(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n698_), .B1(new_n700_), .B2(new_n667_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n697_), .A2(new_n701_), .ZN(G1332gat));
  OR3_X1    g501(.A1(new_n700_), .A2(G64gat), .A3(new_n545_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n695_), .A2(new_n623_), .A3(new_n696_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT48), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n704_), .A2(new_n705_), .A3(G64gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n705_), .B1(new_n704_), .B2(G64gat), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n703_), .B1(new_n706_), .B2(new_n707_), .ZN(G1333gat));
  OR3_X1    g507(.A1(new_n700_), .A2(G71gat), .A3(new_n404_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n695_), .A2(new_n403_), .A3(new_n696_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT49), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n710_), .A2(new_n711_), .A3(G71gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n711_), .B1(new_n710_), .B2(G71gat), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n709_), .B1(new_n712_), .B2(new_n713_), .ZN(G1334gat));
  NAND3_X1  g513(.A1(new_n695_), .A2(new_n634_), .A3(new_n696_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT50), .ZN(new_n716_));
  AND3_X1   g515(.A1(new_n715_), .A2(new_n716_), .A3(G78gat), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n716_), .B1(new_n715_), .B2(G78gat), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n458_), .A2(G78gat), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT112), .ZN(new_n720_));
  OAI22_X1  g519(.A1(new_n717_), .A2(new_n718_), .B1(new_n700_), .B2(new_n720_), .ZN(G1335gat));
  AND3_X1   g520(.A1(new_n661_), .A2(new_n597_), .A3(new_n692_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(new_n601_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n693_), .A2(new_n669_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n667_), .A2(G85gat), .ZN(new_n725_));
  AOI22_X1  g524(.A1(new_n723_), .A2(G85gat), .B1(new_n724_), .B2(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT113), .ZN(G1336gat));
  AOI21_X1  g526(.A(G92gat), .B1(new_n724_), .B2(new_n623_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n623_), .A2(new_n230_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n722_), .B2(new_n729_), .ZN(G1337gat));
  NAND3_X1  g529(.A1(new_n661_), .A2(new_n597_), .A3(new_n692_), .ZN(new_n731_));
  OAI21_X1  g530(.A(G99gat), .B1(new_n731_), .B2(new_n404_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n724_), .A2(new_n227_), .A3(new_n403_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT114), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n734_), .B(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT51), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n736_), .B(new_n737_), .ZN(G1338gat));
  AOI21_X1  g537(.A(new_n214_), .B1(new_n722_), .B2(new_n634_), .ZN(new_n739_));
  OR2_X1    g538(.A1(new_n739_), .A2(KEYINPUT52), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n724_), .A2(new_n214_), .A3(new_n634_), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n741_), .B(KEYINPUT115), .Z(new_n742_));
  NAND2_X1  g541(.A1(new_n739_), .A2(KEYINPUT52), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n740_), .A2(new_n742_), .A3(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g544(.A(new_n539_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n545_), .B1(new_n618_), .B2(new_n617_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT54), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT116), .ZN(new_n750_));
  INV_X1    g549(.A(new_n335_), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n751_), .B(new_n592_), .C1(new_n593_), .C2(new_n596_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n750_), .B1(new_n290_), .B2(new_n753_), .ZN(new_n754_));
  AOI211_X1 g553(.A(KEYINPUT116), .B(new_n752_), .C1(new_n278_), .C2(new_n289_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n749_), .B1(new_n756_), .B2(new_n608_), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n276_), .A2(new_n277_), .A3(new_n287_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n202_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n753_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT116), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n290_), .A2(new_n750_), .A3(new_n753_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n761_), .A2(new_n749_), .A3(new_n608_), .A4(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n757_), .A2(new_n764_), .ZN(new_n765_));
  AOI22_X1  g564(.A1(new_n332_), .A2(new_n334_), .B1(new_n263_), .B2(new_n267_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT55), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n249_), .A2(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(KEYINPUT117), .B1(new_n265_), .B2(new_n204_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT117), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n264_), .A2(new_n770_), .A3(new_n271_), .A4(new_n247_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n265_), .A2(KEYINPUT55), .A3(new_n204_), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n768_), .A2(new_n769_), .A3(new_n771_), .A4(new_n772_), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n773_), .A2(KEYINPUT56), .A3(new_n259_), .ZN(new_n774_));
  AOI21_X1  g573(.A(KEYINPUT56), .B1(new_n773_), .B2(new_n259_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n766_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT118), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n291_), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n779_), .B(new_n317_), .C1(new_n320_), .C2(new_n321_), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n331_), .B(new_n780_), .C1(new_n324_), .C2(new_n779_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n334_), .A2(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n782_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n783_));
  OAI211_X1 g582(.A(KEYINPUT118), .B(new_n766_), .C1(new_n774_), .C2(new_n775_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n778_), .A2(new_n783_), .A3(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n573_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT57), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT119), .ZN(new_n789_));
  AOI22_X1  g588(.A1(new_n774_), .A2(new_n789_), .B1(new_n263_), .B2(new_n267_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n773_), .A2(new_n259_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT56), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n773_), .A2(KEYINPUT56), .A3(new_n259_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n793_), .A2(KEYINPUT119), .A3(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n790_), .A2(new_n795_), .A3(new_n782_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT58), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n796_), .A2(KEYINPUT120), .A3(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n607_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n561_), .A2(new_n567_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT72), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n570_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n606_), .B1(new_n803_), .B2(new_n569_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n799_), .A2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n797_), .A2(KEYINPUT120), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n790_), .A2(new_n795_), .A3(new_n806_), .A4(new_n782_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n798_), .A2(new_n805_), .A3(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n785_), .A2(KEYINPUT57), .A3(new_n573_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n788_), .A2(new_n808_), .A3(new_n809_), .ZN(new_n810_));
  AND2_X1   g609(.A1(new_n810_), .A2(new_n597_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n746_), .B(new_n748_), .C1(new_n765_), .C2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(G113gat), .B1(new_n813_), .B2(new_n335_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT121), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT59), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n761_), .A2(new_n608_), .A3(new_n762_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(KEYINPUT54), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n763_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n810_), .A2(new_n597_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n747_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n816_), .B1(new_n821_), .B2(new_n746_), .ZN(new_n822_));
  AOI22_X1  g621(.A1(new_n818_), .A2(new_n763_), .B1(new_n810_), .B2(new_n597_), .ZN(new_n823_));
  NOR4_X1   g622(.A1(new_n823_), .A2(KEYINPUT59), .A3(new_n539_), .A4(new_n747_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n815_), .B1(new_n822_), .B2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n812_), .A2(KEYINPUT59), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n821_), .A2(new_n816_), .A3(new_n746_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(KEYINPUT121), .A3(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n825_), .A2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n335_), .A2(G113gat), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n830_), .B(KEYINPUT122), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n814_), .B1(new_n829_), .B2(new_n831_), .ZN(G1340gat));
  OAI21_X1  g631(.A(new_n385_), .B1(new_n290_), .B2(KEYINPUT60), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n813_), .B(new_n833_), .C1(KEYINPUT60), .C2(new_n385_), .ZN(new_n834_));
  NOR3_X1   g633(.A1(new_n822_), .A2(new_n824_), .A3(new_n290_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n834_), .B1(new_n835_), .B2(new_n385_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n836_), .B(KEYINPUT123), .ZN(G1341gat));
  AOI21_X1  g636(.A(G127gat), .B1(new_n813_), .B2(new_n609_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n609_), .A2(G127gat), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n839_), .B(KEYINPUT124), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n838_), .B1(new_n829_), .B2(new_n840_), .ZN(G1342gat));
  INV_X1    g640(.A(G134gat), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n842_), .B1(new_n829_), .B2(new_n805_), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n812_), .A2(G134gat), .A3(new_n573_), .ZN(new_n844_));
  OAI21_X1  g643(.A(KEYINPUT125), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT125), .ZN(new_n846_));
  INV_X1    g645(.A(new_n844_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n608_), .B1(new_n825_), .B2(new_n828_), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n846_), .B(new_n847_), .C1(new_n848_), .C2(new_n842_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n845_), .A2(new_n849_), .ZN(G1343gat));
  NOR3_X1   g649(.A1(new_n823_), .A2(new_n540_), .A3(new_n747_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n335_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g652(.A1(new_n851_), .A2(new_n289_), .A3(new_n278_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g654(.A1(new_n851_), .A2(new_n609_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(KEYINPUT61), .B(G155gat), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n856_), .B(new_n857_), .ZN(G1346gat));
  AOI21_X1  g657(.A(G162gat), .B1(new_n851_), .B2(new_n574_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n608_), .A2(new_n564_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n859_), .B1(new_n851_), .B2(new_n860_), .ZN(G1347gat));
  NOR3_X1   g660(.A1(new_n823_), .A2(new_n404_), .A3(new_n634_), .ZN(new_n862_));
  NOR3_X1   g661(.A1(new_n618_), .A2(new_n617_), .A3(new_n545_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n328_), .B1(new_n865_), .B2(new_n335_), .ZN(new_n866_));
  OR2_X1    g665(.A1(new_n866_), .A2(KEYINPUT62), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n865_), .A2(new_n335_), .A3(new_n484_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n866_), .A2(KEYINPUT62), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n867_), .A2(new_n868_), .A3(new_n869_), .ZN(G1348gat));
  NOR2_X1   g669(.A1(new_n864_), .A2(new_n290_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(new_n351_), .ZN(G1349gat));
  NOR2_X1   g671(.A1(new_n864_), .A2(new_n597_), .ZN(new_n873_));
  MUX2_X1   g672(.A(G183gat), .B(new_n493_), .S(new_n873_), .Z(G1350gat));
  NAND3_X1  g673(.A1(new_n865_), .A2(new_n574_), .A3(new_n363_), .ZN(new_n875_));
  OAI21_X1  g674(.A(G190gat), .B1(new_n864_), .B2(new_n608_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(G1351gat));
  NOR2_X1   g676(.A1(new_n823_), .A2(new_n601_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n545_), .A2(new_n540_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n880_), .A2(new_n751_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(new_n330_), .ZN(G1352gat));
  NOR2_X1   g681(.A1(new_n880_), .A2(new_n290_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(new_n258_), .ZN(G1353gat));
  INV_X1    g683(.A(new_n880_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n609_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n887_));
  AND2_X1   g686(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n888_));
  NOR3_X1   g687(.A1(new_n886_), .A2(new_n887_), .A3(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n889_), .B1(new_n886_), .B2(new_n887_), .ZN(G1354gat));
  XOR2_X1   g689(.A(KEYINPUT126), .B(G218gat), .Z(new_n891_));
  NOR3_X1   g690(.A1(new_n880_), .A2(new_n608_), .A3(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n885_), .A2(new_n574_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n892_), .B1(new_n893_), .B2(new_n891_), .ZN(G1355gat));
endmodule


