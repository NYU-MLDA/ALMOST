//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 0 0 1 0 1 0 0 1 0 1 0 1 0 0 1 0 1 1 1 1 0 0 1 1 1 1 1 1 1 0 1 1 1 0 1 1 0 1 0 0 0 0 0 1 0 1 1 1 1 1 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n667_, new_n668_, new_n669_, new_n670_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n769_, new_n770_, new_n771_, new_n773_,
    new_n774_, new_n775_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n904_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n938_, new_n939_, new_n941_, new_n942_,
    new_n943_, new_n944_, new_n945_, new_n947_, new_n948_, new_n950_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n957_, new_n958_,
    new_n959_;
  XOR2_X1   g000(.A(G197gat), .B(G204gat), .Z(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT21), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G197gat), .B(G204gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT21), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G211gat), .B(G218gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n203_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  OR3_X1    g007(.A1(new_n204_), .A2(new_n207_), .A3(new_n205_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT91), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT91), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n208_), .A2(new_n212_), .A3(new_n209_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G141gat), .A2(G148gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT3), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n215_), .A2(KEYINPUT88), .A3(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G141gat), .A2(G148gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT2), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT88), .ZN(new_n221_));
  OAI22_X1  g020(.A1(new_n221_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n217_), .A2(new_n220_), .A3(new_n222_), .A4(new_n223_), .ZN(new_n224_));
  XOR2_X1   g023(.A(G155gat), .B(G162gat), .Z(new_n225_));
  INV_X1    g024(.A(G155gat), .ZN(new_n226_));
  INV_X1    g025(.A(G162gat), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT1), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT1), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n229_), .A2(G155gat), .A3(G162gat), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n228_), .B(new_n230_), .C1(G155gat), .C2(G162gat), .ZN(new_n231_));
  INV_X1    g030(.A(new_n215_), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n232_), .A2(new_n218_), .ZN(new_n233_));
  AOI22_X1  g032(.A1(new_n224_), .A2(new_n225_), .B1(new_n231_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT29), .ZN(new_n235_));
  INV_X1    g034(.A(G228gat), .ZN(new_n236_));
  INV_X1    g035(.A(G233gat), .ZN(new_n237_));
  OAI22_X1  g036(.A1(new_n234_), .A2(new_n235_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n214_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT92), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n210_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n236_), .A2(new_n237_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n240_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n241_), .A2(new_n240_), .A3(new_n242_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n239_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G78gat), .B(G106gat), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n245_), .ZN(new_n250_));
  OAI22_X1  g049(.A1(new_n250_), .A2(new_n243_), .B1(new_n214_), .B2(new_n238_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(new_n247_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n249_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G22gat), .B(G50gat), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  XOR2_X1   g054(.A(KEYINPUT90), .B(KEYINPUT28), .Z(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(KEYINPUT89), .B1(new_n234_), .B2(new_n235_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n234_), .A2(KEYINPUT89), .A3(new_n235_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n257_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n260_), .ZN(new_n262_));
  NOR3_X1   g061(.A1(new_n262_), .A2(new_n258_), .A3(new_n256_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n255_), .B1(new_n261_), .B2(new_n263_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n256_), .B1(new_n262_), .B2(new_n258_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n259_), .A2(new_n260_), .A3(new_n257_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n265_), .A2(new_n266_), .A3(new_n254_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n264_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n253_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT93), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n268_), .B1(new_n252_), .B2(new_n249_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT93), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT94), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n275_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n251_), .A2(KEYINPUT94), .A3(new_n247_), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n276_), .A2(new_n277_), .A3(new_n268_), .A4(new_n249_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n272_), .A2(new_n274_), .A3(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT27), .ZN(new_n280_));
  XNOR2_X1  g079(.A(KEYINPUT26), .B(G190gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT25), .B(G183gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT24), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n284_), .B1(G169gat), .B2(G176gat), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n285_), .B1(G169gat), .B2(G176gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n283_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT80), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n283_), .A2(new_n286_), .A3(KEYINPUT80), .ZN(new_n290_));
  INV_X1    g089(.A(G183gat), .ZN(new_n291_));
  INV_X1    g090(.A(G190gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT23), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT23), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n294_), .A2(G183gat), .A3(G190gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  OR3_X1    g095(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(KEYINPUT81), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT81), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n296_), .A2(new_n300_), .A3(new_n297_), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n289_), .A2(new_n290_), .A3(new_n299_), .A4(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT82), .ZN(new_n303_));
  OR2_X1    g102(.A1(new_n295_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n293_), .A2(new_n303_), .A3(new_n295_), .ZN(new_n305_));
  OAI211_X1 g104(.A(new_n304_), .B(new_n305_), .C1(G183gat), .C2(G190gat), .ZN(new_n306_));
  NOR2_X1   g105(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(G169gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n302_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(new_n214_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n282_), .B(KEYINPUT95), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(new_n281_), .ZN(new_n314_));
  AND4_X1   g113(.A1(new_n304_), .A2(new_n286_), .A3(new_n305_), .A4(new_n297_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n296_), .B1(G183gat), .B2(G190gat), .ZN(new_n316_));
  AOI22_X1  g115(.A1(new_n314_), .A2(new_n315_), .B1(new_n308_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n318_), .A2(KEYINPUT96), .A3(new_n210_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT96), .ZN(new_n320_));
  INV_X1    g119(.A(new_n210_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n320_), .B1(new_n317_), .B2(new_n321_), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n312_), .A2(new_n319_), .A3(KEYINPUT20), .A4(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G226gat), .A2(G233gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT19), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n323_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n325_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT20), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n328_), .B1(new_n317_), .B2(new_n321_), .ZN(new_n329_));
  NOR3_X1   g128(.A1(new_n311_), .A2(KEYINPUT97), .A3(new_n214_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT97), .ZN(new_n331_));
  AND2_X1   g130(.A1(new_n211_), .A2(new_n213_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n331_), .B1(new_n332_), .B2(new_n310_), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n327_), .B(new_n329_), .C1(new_n330_), .C2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G8gat), .B(G36gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT18), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G64gat), .B(G92gat), .ZN(new_n337_));
  XOR2_X1   g136(.A(new_n336_), .B(new_n337_), .Z(new_n338_));
  AND3_X1   g137(.A1(new_n326_), .A2(new_n334_), .A3(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n338_), .B1(new_n326_), .B2(new_n334_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n280_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  XOR2_X1   g140(.A(G127gat), .B(G134gat), .Z(new_n342_));
  XOR2_X1   g141(.A(G113gat), .B(G120gat), .Z(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G127gat), .B(G134gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G113gat), .B(G120gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n344_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT84), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n344_), .A2(KEYINPUT84), .A3(new_n347_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n234_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  OR2_X1    g151(.A1(new_n352_), .A2(KEYINPUT4), .ZN(new_n353_));
  AND2_X1   g152(.A1(new_n234_), .A2(new_n348_), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT4), .B1(new_n352_), .B2(new_n354_), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n353_), .A2(new_n355_), .A3(G225gat), .A4(G233gat), .ZN(new_n356_));
  OR2_X1    g155(.A1(new_n352_), .A2(new_n354_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G225gat), .A2(G233gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n356_), .A2(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G1gat), .B(G29gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(G85gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT0), .B(G57gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n360_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n356_), .A2(new_n359_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n364_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n365_), .A2(KEYINPUT100), .A3(new_n368_), .ZN(new_n369_));
  OR3_X1    g168(.A1(new_n366_), .A2(KEYINPUT100), .A3(new_n367_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n328_), .B1(new_n311_), .B2(new_n214_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n372_), .A2(new_n327_), .A3(new_n319_), .A4(new_n322_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n329_), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT97), .B1(new_n311_), .B2(new_n214_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n332_), .A2(new_n310_), .A3(new_n331_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n374_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n373_), .B1(new_n377_), .B2(new_n327_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n338_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n326_), .A2(new_n334_), .A3(new_n338_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n380_), .A2(KEYINPUT27), .A3(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n341_), .A2(new_n371_), .A3(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n302_), .A2(KEYINPUT30), .A3(new_n309_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(KEYINPUT30), .B1(new_n302_), .B2(new_n309_), .ZN(new_n386_));
  OAI21_X1  g185(.A(KEYINPUT83), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n386_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT83), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n388_), .A2(new_n389_), .A3(new_n384_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G71gat), .B(G99gat), .ZN(new_n391_));
  INV_X1    g190(.A(G43gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G227gat), .A2(G233gat), .ZN(new_n394_));
  INV_X1    g193(.A(G15gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n393_), .B(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n387_), .A2(new_n390_), .A3(new_n398_), .ZN(new_n399_));
  AND2_X1   g198(.A1(new_n350_), .A2(new_n351_), .ZN(new_n400_));
  XOR2_X1   g199(.A(new_n400_), .B(KEYINPUT31), .Z(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n388_), .A2(new_n389_), .A3(new_n384_), .A4(new_n397_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n399_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT85), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n404_), .A2(new_n405_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT86), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n399_), .A2(new_n403_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n408_), .B1(new_n409_), .B2(new_n401_), .ZN(new_n410_));
  AOI211_X1 g209(.A(KEYINPUT86), .B(new_n402_), .C1(new_n399_), .C2(new_n403_), .ZN(new_n411_));
  OAI22_X1  g210(.A1(new_n406_), .A2(new_n407_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT87), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT87), .ZN(new_n414_));
  OAI221_X1 g213(.A(new_n414_), .B1(new_n410_), .B2(new_n411_), .C1(new_n406_), .C2(new_n407_), .ZN(new_n415_));
  AOI211_X1 g214(.A(new_n279_), .B(new_n383_), .C1(new_n413_), .C2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n326_), .A2(new_n334_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(new_n379_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n364_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n353_), .A2(new_n355_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n419_), .B1(new_n358_), .B2(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n364_), .B1(new_n356_), .B2(new_n359_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n421_), .B1(KEYINPUT33), .B2(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n418_), .A2(new_n423_), .A3(new_n381_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT98), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT33), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n368_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT98), .B1(new_n422_), .B2(KEYINPUT33), .ZN(new_n428_));
  AND2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT99), .B1(new_n424_), .B2(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n339_), .A2(new_n340_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT99), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n427_), .A2(new_n428_), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n431_), .A2(new_n432_), .A3(new_n433_), .A4(new_n423_), .ZN(new_n434_));
  AND2_X1   g233(.A1(new_n338_), .A2(KEYINPUT32), .ZN(new_n435_));
  OR2_X1    g234(.A1(new_n417_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n378_), .A2(new_n435_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n436_), .A2(new_n370_), .A3(new_n369_), .A4(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n430_), .A2(new_n434_), .A3(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n278_), .B1(new_n273_), .B2(KEYINPUT93), .ZN(new_n440_));
  AND3_X1   g239(.A1(new_n253_), .A2(KEYINPUT93), .A3(new_n269_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n439_), .A2(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT101), .B1(new_n383_), .B2(new_n442_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  NOR3_X1   g245(.A1(new_n383_), .A2(new_n442_), .A3(KEYINPUT101), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n413_), .A2(new_n415_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n416_), .B1(new_n446_), .B2(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G113gat), .B(G141gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G169gat), .B(G197gat), .ZN(new_n452_));
  XOR2_X1   g251(.A(new_n451_), .B(new_n452_), .Z(new_n453_));
  XNOR2_X1  g252(.A(G29gat), .B(G36gat), .ZN(new_n454_));
  XOR2_X1   g253(.A(new_n454_), .B(KEYINPUT70), .Z(new_n455_));
  XNOR2_X1  g254(.A(G43gat), .B(G50gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n454_), .B(KEYINPUT70), .ZN(new_n458_));
  INV_X1    g257(.A(new_n456_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n457_), .A2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G1gat), .B(G8gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(KEYINPUT75), .ZN(new_n463_));
  INV_X1    g262(.A(G1gat), .ZN(new_n464_));
  INV_X1    g263(.A(G8gat), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT14), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT74), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  OAI211_X1 g267(.A(KEYINPUT74), .B(KEYINPUT14), .C1(new_n464_), .C2(new_n465_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G15gat), .B(G22gat), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n468_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n463_), .B(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n461_), .B(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G229gat), .A2(G233gat), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n473_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT15), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n461_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n472_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n457_), .A2(new_n460_), .A3(KEYINPUT15), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n478_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n461_), .A2(new_n472_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n481_), .A2(new_n482_), .A3(new_n474_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n476_), .A2(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n453_), .B1(new_n484_), .B2(KEYINPUT79), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT79), .ZN(new_n486_));
  INV_X1    g285(.A(new_n453_), .ZN(new_n487_));
  AOI211_X1 g286(.A(new_n486_), .B(new_n487_), .C1(new_n476_), .C2(new_n483_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n485_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G120gat), .B(G148gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT5), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G176gat), .B(G204gat), .ZN(new_n493_));
  XOR2_X1   g292(.A(new_n492_), .B(new_n493_), .Z(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G99gat), .A2(G106gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(KEYINPUT6), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT6), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n498_), .A2(G99gat), .A3(G106gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n497_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT65), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n497_), .A2(new_n499_), .A3(KEYINPUT65), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  XOR2_X1   g303(.A(KEYINPUT10), .B(G99gat), .Z(new_n505_));
  INV_X1    g304(.A(G106gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(G85gat), .ZN(new_n508_));
  INV_X1    g307(.A(G92gat), .ZN(new_n509_));
  NOR3_X1   g308(.A1(new_n508_), .A2(new_n509_), .A3(KEYINPUT9), .ZN(new_n510_));
  XOR2_X1   g309(.A(G85gat), .B(G92gat), .Z(new_n511_));
  AOI21_X1  g310(.A(new_n510_), .B1(new_n511_), .B2(KEYINPUT9), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n504_), .A2(new_n507_), .A3(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT8), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n511_), .A2(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(G99gat), .A2(G106gat), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT7), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT66), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n518_), .A2(KEYINPUT66), .A3(new_n519_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n517_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n515_), .B1(new_n504_), .B2(new_n524_), .ZN(new_n525_));
  NOR4_X1   g324(.A1(new_n521_), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n526_));
  AOI21_X1  g325(.A(KEYINPUT66), .B1(new_n518_), .B2(new_n519_), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n500_), .B(new_n516_), .C1(new_n526_), .C2(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n514_), .B1(new_n528_), .B2(new_n511_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n513_), .B1(new_n525_), .B2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(KEYINPUT67), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT67), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n532_), .B(new_n513_), .C1(new_n525_), .C2(new_n529_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G57gat), .B(G64gat), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(KEYINPUT11), .ZN(new_n535_));
  XOR2_X1   g334(.A(G71gat), .B(G78gat), .Z(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n534_), .A2(KEYINPUT11), .ZN(new_n538_));
  OR2_X1    g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  OR2_X1    g338(.A1(new_n535_), .A2(new_n536_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n531_), .A2(new_n533_), .A3(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G230gat), .A2(G233gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT64), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n541_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n528_), .A2(new_n511_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(KEYINPUT8), .ZN(new_n548_));
  INV_X1    g347(.A(new_n515_), .ZN(new_n549_));
  AND3_X1   g348(.A1(new_n497_), .A2(new_n499_), .A3(KEYINPUT65), .ZN(new_n550_));
  AOI21_X1  g349(.A(KEYINPUT65), .B1(new_n497_), .B2(new_n499_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n516_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n549_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n548_), .A2(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n532_), .B1(new_n555_), .B2(new_n513_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n533_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n546_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  XOR2_X1   g357(.A(KEYINPUT69), .B(KEYINPUT12), .Z(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n546_), .A2(new_n530_), .A3(KEYINPUT12), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n545_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n544_), .ZN(new_n564_));
  OAI211_X1 g363(.A(KEYINPUT68), .B(new_n546_), .C1(new_n556_), .C2(new_n557_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT68), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n542_), .A2(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n541_), .B1(new_n531_), .B2(new_n533_), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n564_), .B(new_n565_), .C1(new_n567_), .C2(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n495_), .B1(new_n563_), .B2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n563_), .A2(new_n569_), .A3(new_n495_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n571_), .A2(KEYINPUT13), .A3(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT13), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n563_), .A2(new_n569_), .A3(new_n495_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n574_), .B1(new_n575_), .B2(new_n570_), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n573_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G231gat), .A2(G233gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n541_), .B(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(new_n479_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G127gat), .B(G155gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT16), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G183gat), .B(G211gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(KEYINPUT76), .B(KEYINPUT17), .Z(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT77), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n580_), .A2(new_n587_), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n588_), .A2(KEYINPUT78), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(KEYINPUT78), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n584_), .B(KEYINPUT17), .Z(new_n592_));
  NAND2_X1  g391(.A1(new_n580_), .A2(new_n592_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT73), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT37), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n531_), .A2(new_n461_), .A3(new_n533_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT71), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n531_), .A2(KEYINPUT71), .A3(new_n461_), .A4(new_n533_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(G232gat), .A2(G233gat), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n602_), .B(KEYINPUT34), .Z(new_n603_));
  INV_X1    g402(.A(KEYINPUT35), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n603_), .A2(new_n604_), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n607_), .B(KEYINPUT72), .Z(new_n608_));
  AND2_X1   g407(.A1(new_n478_), .A2(new_n480_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n608_), .B1(new_n609_), .B2(new_n530_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n601_), .A2(new_n606_), .A3(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n606_), .B1(new_n601_), .B2(new_n610_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G190gat), .B(G218gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G134gat), .B(G162gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n616_), .A2(KEYINPUT36), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NOR3_X1   g417(.A1(new_n612_), .A2(new_n613_), .A3(new_n618_), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n616_), .B(KEYINPUT36), .Z(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n601_), .A2(new_n610_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(new_n605_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n621_), .B1(new_n623_), .B2(new_n611_), .ZN(new_n624_));
  OAI211_X1 g423(.A(new_n595_), .B(new_n596_), .C1(new_n619_), .C2(new_n624_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n620_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n623_), .A2(new_n617_), .A3(new_n611_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(KEYINPUT73), .A2(KEYINPUT37), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n595_), .A2(new_n596_), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n626_), .A2(new_n627_), .A3(new_n628_), .A4(new_n629_), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n577_), .A2(new_n594_), .A3(new_n625_), .A4(new_n630_), .ZN(new_n631_));
  NOR3_X1   g430(.A1(new_n450_), .A2(new_n490_), .A3(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT102), .ZN(new_n633_));
  INV_X1    g432(.A(new_n371_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n633_), .A2(new_n464_), .A3(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT38), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n619_), .A2(new_n624_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n450_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n573_), .A2(new_n576_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n640_), .A2(new_n490_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(new_n594_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT103), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n639_), .A2(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT104), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n464_), .B1(new_n645_), .B2(new_n634_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n635_), .A2(new_n636_), .ZN(new_n647_));
  OR3_X1    g446(.A1(new_n637_), .A2(new_n646_), .A3(new_n647_), .ZN(G1324gat));
  INV_X1    g447(.A(KEYINPUT40), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT105), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n341_), .A2(new_n382_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n644_), .A2(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n650_), .B1(new_n652_), .B2(G8gat), .ZN(new_n653_));
  AOI211_X1 g452(.A(KEYINPUT105), .B(new_n465_), .C1(new_n644_), .C2(new_n651_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT39), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n653_), .A2(new_n654_), .A3(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n652_), .A2(G8gat), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n657_), .A2(KEYINPUT105), .A3(new_n655_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n633_), .A2(new_n465_), .A3(new_n651_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n649_), .B1(new_n656_), .B2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n653_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n652_), .A2(new_n650_), .A3(G8gat), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n662_), .A2(KEYINPUT39), .A3(new_n663_), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n664_), .A2(KEYINPUT40), .A3(new_n658_), .A4(new_n659_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n661_), .A2(new_n665_), .ZN(G1325gat));
  NAND3_X1  g465(.A1(new_n633_), .A2(new_n395_), .A3(new_n448_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n645_), .A2(new_n448_), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n668_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(KEYINPUT41), .B1(new_n668_), .B2(G15gat), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n667_), .B1(new_n669_), .B2(new_n670_), .ZN(G1326gat));
  INV_X1    g470(.A(G22gat), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n633_), .A2(new_n672_), .A3(new_n279_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n672_), .B1(new_n645_), .B2(new_n279_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT42), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n674_), .A2(new_n675_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n673_), .B1(new_n676_), .B2(new_n677_), .ZN(G1327gat));
  NOR2_X1   g477(.A1(new_n450_), .A2(new_n490_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n591_), .A2(new_n593_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(new_n638_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n681_), .A2(new_n640_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n679_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(G29gat), .B1(new_n684_), .B2(new_n634_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT43), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n625_), .A2(new_n630_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n686_), .B1(new_n450_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n651_), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n448_), .A2(new_n442_), .A3(new_n371_), .A4(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n444_), .B1(new_n442_), .B2(new_n439_), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n279_), .A2(new_n371_), .A3(new_n341_), .A4(new_n382_), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n413_), .B(new_n415_), .C1(new_n693_), .C2(KEYINPUT101), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n691_), .B1(new_n692_), .B2(new_n694_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n695_), .A2(KEYINPUT43), .A3(new_n687_), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n689_), .A2(new_n680_), .A3(new_n641_), .A4(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n695_), .A2(new_n687_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n594_), .B1(new_n700_), .B2(new_n686_), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n701_), .A2(KEYINPUT44), .A3(new_n641_), .A4(new_n696_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n699_), .A2(new_n702_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n634_), .A2(G29gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n685_), .B1(new_n703_), .B2(new_n704_), .ZN(G1328gat));
  NAND3_X1  g504(.A1(new_n699_), .A2(new_n651_), .A3(new_n702_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(G36gat), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n690_), .A2(G36gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n679_), .A2(new_n682_), .A3(new_n708_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n709_), .B(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n707_), .A2(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(KEYINPUT46), .B1(new_n713_), .B2(KEYINPUT107), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n711_), .B1(new_n706_), .B2(G36gat), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT107), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT46), .ZN(new_n717_));
  NOR3_X1   g516(.A1(new_n715_), .A2(new_n716_), .A3(new_n717_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n714_), .A2(new_n718_), .ZN(G1329gat));
  NAND4_X1  g518(.A1(new_n699_), .A2(new_n702_), .A3(G43gat), .A4(new_n448_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n448_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n392_), .B1(new_n683_), .B2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g523(.A(G50gat), .B1(new_n684_), .B2(new_n279_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n279_), .A2(G50gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n703_), .B2(new_n726_), .ZN(G1331gat));
  NOR2_X1   g526(.A1(new_n450_), .A2(new_n489_), .ZN(new_n728_));
  NOR3_X1   g527(.A1(new_n687_), .A2(new_n577_), .A3(new_n680_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  OR2_X1    g530(.A1(new_n731_), .A2(KEYINPUT108), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(KEYINPUT108), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n732_), .A2(new_n634_), .A3(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(G57gat), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n577_), .A2(new_n489_), .A3(new_n680_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n639_), .A2(new_n736_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n371_), .A2(new_n735_), .ZN(new_n738_));
  AOI22_X1  g537(.A1(new_n734_), .A2(new_n735_), .B1(new_n737_), .B2(new_n738_), .ZN(G1332gat));
  INV_X1    g538(.A(G64gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(new_n737_), .B2(new_n651_), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n741_), .B(KEYINPUT48), .Z(new_n742_));
  NAND3_X1  g541(.A1(new_n731_), .A2(new_n740_), .A3(new_n651_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(G1333gat));
  INV_X1    g543(.A(G71gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n737_), .B2(new_n448_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT49), .Z(new_n747_));
  NAND3_X1  g546(.A1(new_n731_), .A2(new_n745_), .A3(new_n448_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(G1334gat));
  OR3_X1    g548(.A1(new_n730_), .A2(G78gat), .A3(new_n442_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n737_), .A2(new_n279_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(G78gat), .ZN(new_n752_));
  OR2_X1    g551(.A1(new_n752_), .A2(KEYINPUT110), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(KEYINPUT110), .ZN(new_n754_));
  XOR2_X1   g553(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n755_));
  AND3_X1   g554(.A1(new_n753_), .A2(new_n754_), .A3(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n750_), .B1(new_n756_), .B2(new_n757_), .ZN(G1335gat));
  NOR2_X1   g557(.A1(new_n577_), .A2(new_n489_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n701_), .A2(new_n696_), .A3(new_n759_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n371_), .A2(new_n508_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT112), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n760_), .A2(new_n762_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n681_), .A2(new_n577_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n728_), .A2(new_n764_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT111), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(new_n634_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n763_), .B1(new_n767_), .B2(new_n508_), .ZN(G1336gat));
  NAND3_X1  g567(.A1(new_n766_), .A2(new_n509_), .A3(new_n651_), .ZN(new_n769_));
  OAI21_X1  g568(.A(G92gat), .B1(new_n760_), .B2(new_n690_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT113), .ZN(G1337gat));
  NAND3_X1  g571(.A1(new_n766_), .A2(new_n448_), .A3(new_n505_), .ZN(new_n773_));
  OAI21_X1  g572(.A(G99gat), .B1(new_n760_), .B2(new_n721_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g575(.A1(new_n766_), .A2(new_n506_), .A3(new_n279_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n701_), .A2(new_n279_), .A3(new_n696_), .A4(new_n759_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n778_), .A2(new_n779_), .A3(G106gat), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n779_), .B1(new_n778_), .B2(G106gat), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n777_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT53), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n777_), .B(new_n785_), .C1(new_n782_), .C2(new_n781_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(G1339gat));
  NOR2_X1   g586(.A1(new_n721_), .A2(new_n279_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n651_), .A2(new_n371_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n790_), .A2(KEYINPUT59), .ZN(new_n791_));
  NOR3_X1   g590(.A1(new_n687_), .A2(new_n640_), .A3(new_n680_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n792_), .A2(new_n793_), .A3(new_n490_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(KEYINPUT114), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n631_), .A2(new_n489_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT114), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n796_), .A2(new_n797_), .A3(new_n793_), .ZN(new_n798_));
  OAI21_X1  g597(.A(KEYINPUT54), .B1(new_n631_), .B2(new_n489_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n795_), .A2(new_n798_), .A3(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n638_), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n473_), .A2(new_n474_), .ZN(new_n802_));
  AND3_X1   g601(.A1(new_n481_), .A2(new_n482_), .A3(new_n475_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n487_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n484_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n804_), .B1(new_n805_), .B2(new_n487_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n806_), .B1(new_n575_), .B2(new_n570_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(KEYINPUT116), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT116), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n809_), .B(new_n806_), .C1(new_n575_), .C2(new_n570_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n808_), .A2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n489_), .A2(new_n572_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n562_), .B1(new_n568_), .B2(new_n559_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n542_), .A2(new_n544_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n813_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n545_), .A2(new_n561_), .A3(KEYINPUT55), .A4(new_n562_), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n562_), .B(new_n542_), .C1(new_n568_), .C2(new_n559_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n564_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n816_), .A2(new_n817_), .A3(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n494_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT56), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n820_), .A2(KEYINPUT56), .A3(new_n494_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n812_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n811_), .B1(new_n825_), .B2(KEYINPUT115), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n575_), .A2(new_n488_), .A3(new_n485_), .ZN(new_n827_));
  AND3_X1   g626(.A1(new_n820_), .A2(KEYINPUT56), .A3(new_n494_), .ZN(new_n828_));
  AOI21_X1  g627(.A(KEYINPUT56), .B1(new_n820_), .B2(new_n494_), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n827_), .B(KEYINPUT115), .C1(new_n828_), .C2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n801_), .B1(new_n826_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT57), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n827_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT115), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n837_), .A2(new_n830_), .A3(new_n811_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n638_), .A2(new_n833_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n806_), .A2(new_n572_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n840_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n841_));
  AOI22_X1  g640(.A1(new_n841_), .A2(KEYINPUT58), .B1(new_n630_), .B2(new_n625_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT58), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n828_), .A2(new_n829_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n843_), .B1(new_n844_), .B2(new_n840_), .ZN(new_n845_));
  AOI22_X1  g644(.A1(new_n838_), .A2(new_n839_), .B1(new_n842_), .B2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n594_), .B1(new_n834_), .B2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n800_), .B1(new_n847_), .B2(KEYINPUT118), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n838_), .A2(new_n839_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n842_), .A2(new_n845_), .ZN(new_n850_));
  AOI22_X1  g649(.A1(new_n835_), .A2(new_n836_), .B1(new_n808_), .B2(new_n810_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n638_), .B1(new_n851_), .B2(new_n830_), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n849_), .B(new_n850_), .C1(new_n852_), .C2(KEYINPUT57), .ZN(new_n853_));
  AND3_X1   g652(.A1(new_n853_), .A2(KEYINPUT118), .A3(new_n680_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n791_), .B1(new_n848_), .B2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT119), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n797_), .B1(new_n796_), .B2(new_n793_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n799_), .ZN(new_n859_));
  NOR4_X1   g658(.A1(new_n631_), .A2(KEYINPUT114), .A3(KEYINPUT54), .A4(new_n489_), .ZN(new_n860_));
  NOR3_X1   g659(.A1(new_n858_), .A2(new_n859_), .A3(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT117), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n594_), .B1(new_n853_), .B2(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n834_), .A2(KEYINPUT117), .A3(new_n846_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n861_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  OAI21_X1  g664(.A(KEYINPUT59), .B1(new_n865_), .B2(new_n790_), .ZN(new_n866_));
  OAI211_X1 g665(.A(KEYINPUT119), .B(new_n791_), .C1(new_n848_), .C2(new_n854_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n857_), .A2(new_n866_), .A3(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(G113gat), .B1(new_n868_), .B2(new_n490_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n849_), .A2(new_n850_), .ZN(new_n870_));
  AOI21_X1  g669(.A(KEYINPUT57), .B1(new_n838_), .B2(new_n801_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n862_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n872_), .A2(new_n680_), .A3(new_n864_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(new_n800_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n874_), .A2(new_n788_), .A3(new_n789_), .ZN(new_n875_));
  OR2_X1    g674(.A1(new_n490_), .A2(G113gat), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n869_), .B1(new_n875_), .B2(new_n876_), .ZN(G1340gat));
  OAI21_X1  g676(.A(G120gat), .B1(new_n868_), .B2(new_n577_), .ZN(new_n878_));
  INV_X1    g677(.A(G120gat), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n879_), .B1(new_n577_), .B2(KEYINPUT60), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n880_), .B1(KEYINPUT60), .B2(new_n879_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n878_), .B1(new_n875_), .B2(new_n881_), .ZN(G1341gat));
  INV_X1    g681(.A(G127gat), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n680_), .A2(new_n883_), .ZN(new_n884_));
  NAND4_X1  g683(.A1(new_n857_), .A2(new_n866_), .A3(new_n867_), .A4(new_n884_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n883_), .B1(new_n875_), .B2(new_n680_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(KEYINPUT120), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT120), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n885_), .A2(new_n889_), .A3(new_n886_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n888_), .A2(new_n890_), .ZN(G1342gat));
  OAI21_X1  g690(.A(G134gat), .B1(new_n868_), .B2(new_n688_), .ZN(new_n892_));
  OR2_X1    g691(.A1(new_n801_), .A2(G134gat), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n875_), .B2(new_n893_), .ZN(G1343gat));
  INV_X1    g693(.A(KEYINPUT121), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n448_), .A2(new_n442_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n789_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n895_), .B1(new_n865_), .B2(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n897_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n874_), .A2(KEYINPUT121), .A3(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n489_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g702(.A1(new_n901_), .A2(new_n640_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(G148gat), .ZN(G1345gat));
  AOI21_X1  g704(.A(new_n680_), .B1(new_n898_), .B2(new_n900_), .ZN(new_n906_));
  XOR2_X1   g705(.A(KEYINPUT61), .B(G155gat), .Z(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(KEYINPUT122), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(KEYINPUT123), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n906_), .B(new_n909_), .ZN(G1346gat));
  NAND2_X1  g709(.A1(new_n687_), .A2(G162gat), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(KEYINPUT125), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n912_), .B1(new_n898_), .B2(new_n900_), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT124), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n801_), .B1(new_n898_), .B2(new_n900_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n914_), .B1(new_n915_), .B2(G162gat), .ZN(new_n916_));
  AOI21_X1  g715(.A(KEYINPUT121), .B1(new_n874_), .B2(new_n899_), .ZN(new_n917_));
  AOI211_X1 g716(.A(new_n895_), .B(new_n897_), .C1(new_n873_), .C2(new_n800_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n638_), .B1(new_n917_), .B2(new_n918_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n919_), .A2(KEYINPUT124), .A3(new_n227_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n913_), .B1(new_n916_), .B2(new_n920_), .ZN(G1347gat));
  NOR2_X1   g720(.A1(new_n690_), .A2(new_n634_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(new_n448_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(KEYINPUT126), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n924_), .A2(new_n279_), .ZN(new_n925_));
  OAI211_X1 g724(.A(new_n489_), .B(new_n925_), .C1(new_n848_), .C2(new_n854_), .ZN(new_n926_));
  OAI21_X1  g725(.A(G169gat), .B1(new_n926_), .B2(KEYINPUT62), .ZN(new_n927_));
  OAI21_X1  g726(.A(KEYINPUT62), .B1(new_n926_), .B2(KEYINPUT22), .ZN(new_n928_));
  MUX2_X1   g727(.A(G169gat), .B(new_n927_), .S(new_n928_), .Z(G1348gat));
  OR2_X1    g728(.A1(new_n848_), .A2(new_n854_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n930_), .A2(new_n925_), .ZN(new_n931_));
  INV_X1    g730(.A(new_n931_), .ZN(new_n932_));
  AOI21_X1  g731(.A(G176gat), .B1(new_n932_), .B2(new_n640_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n865_), .A2(new_n279_), .ZN(new_n934_));
  INV_X1    g733(.A(new_n924_), .ZN(new_n935_));
  AND3_X1   g734(.A1(new_n935_), .A2(G176gat), .A3(new_n640_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n933_), .B1(new_n934_), .B2(new_n936_), .ZN(G1349gat));
  NOR3_X1   g736(.A1(new_n931_), .A2(new_n313_), .A3(new_n680_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n934_), .A2(new_n594_), .A3(new_n935_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n938_), .B1(new_n291_), .B2(new_n939_), .ZN(G1350gat));
  NAND3_X1  g739(.A1(new_n930_), .A2(new_n687_), .A3(new_n925_), .ZN(new_n941_));
  INV_X1    g740(.A(KEYINPUT127), .ZN(new_n942_));
  AND3_X1   g741(.A1(new_n941_), .A2(new_n942_), .A3(G190gat), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n942_), .B1(new_n941_), .B2(G190gat), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n638_), .A2(new_n281_), .ZN(new_n945_));
  OAI22_X1  g744(.A1(new_n943_), .A2(new_n944_), .B1(new_n931_), .B2(new_n945_), .ZN(G1351gat));
  AND3_X1   g745(.A1(new_n874_), .A2(new_n896_), .A3(new_n922_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n947_), .A2(new_n489_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g748(.A1(new_n947_), .A2(new_n640_), .ZN(new_n950_));
  XNOR2_X1  g749(.A(new_n950_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g750(.A1(new_n947_), .A2(new_n594_), .ZN(new_n952_));
  XNOR2_X1  g751(.A(KEYINPUT63), .B(G211gat), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n952_), .A2(new_n953_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n954_), .B1(new_n952_), .B2(new_n955_), .ZN(G1354gat));
  INV_X1    g755(.A(G218gat), .ZN(new_n957_));
  NAND3_X1  g756(.A1(new_n947_), .A2(new_n957_), .A3(new_n638_), .ZN(new_n958_));
  AND2_X1   g757(.A1(new_n947_), .A2(new_n687_), .ZN(new_n959_));
  OAI21_X1  g758(.A(new_n958_), .B1(new_n959_), .B2(new_n957_), .ZN(G1355gat));
endmodule


