//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 0 1 0 1 0 1 0 0 0 0 1 0 0 1 0 1 0 0 0 1 1 1 1 1 0 1 1 1 1 1 1 1 1 0 1 1 1 1 1 1 1 0 0 1 1 1 1 1 1 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n789_, new_n790_,
    new_n791_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n915_, new_n916_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n923_, new_n925_,
    new_n926_, new_n928_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n945_, new_n946_, new_n947_,
    new_n949_, new_n950_, new_n951_, new_n953_, new_n954_, new_n956_,
    new_n957_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n965_, new_n966_, new_n967_;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G169gat), .B(G197gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G229gat), .A2(G233gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G15gat), .B(G22gat), .ZN(new_n207_));
  INV_X1    g006(.A(G1gat), .ZN(new_n208_));
  INV_X1    g007(.A(G8gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT14), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n207_), .A2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G1gat), .B(G8gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n211_), .B(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G29gat), .B(G36gat), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n215_), .A2(KEYINPUT70), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(KEYINPUT70), .ZN(new_n217_));
  XNOR2_X1  g016(.A(G43gat), .B(G50gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n216_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n215_), .B(KEYINPUT70), .ZN(new_n220_));
  INV_X1    g019(.A(new_n218_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n214_), .A2(new_n219_), .A3(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n219_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(new_n213_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n206_), .B1(new_n223_), .B2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT15), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n224_), .A2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n222_), .A2(KEYINPUT15), .A3(new_n219_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(new_n213_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n224_), .A2(new_n213_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n206_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  AOI211_X1 g033(.A(new_n205_), .B(new_n226_), .C1(new_n231_), .C2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n231_), .A2(new_n234_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n226_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n204_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n235_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G227gat), .A2(G233gat), .ZN(new_n240_));
  INV_X1    g039(.A(G15gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(G71gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT76), .B(G43gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(G99gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n243_), .B(new_n245_), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n246_), .A2(KEYINPUT77), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(KEYINPUT77), .ZN(new_n248_));
  NOR2_X1   g047(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(G169gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G183gat), .A2(G190gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT23), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT23), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n253_), .A2(G183gat), .A3(G190gat), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT75), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n252_), .A2(new_n254_), .A3(new_n255_), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n253_), .A2(KEYINPUT75), .A3(G183gat), .A4(G190gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(G183gat), .A2(G190gat), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n250_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT25), .B(G183gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT26), .B(G190gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  OR2_X1    g062(.A1(G169gat), .A2(G176gat), .ZN(new_n264_));
  OR2_X1    g063(.A1(new_n264_), .A2(KEYINPUT24), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n252_), .A2(new_n254_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G169gat), .A2(G176gat), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n264_), .A2(KEYINPUT24), .A3(new_n267_), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n263_), .A2(new_n265_), .A3(new_n266_), .A4(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n260_), .A2(new_n269_), .ZN(new_n270_));
  XOR2_X1   g069(.A(new_n270_), .B(KEYINPUT30), .Z(new_n271_));
  NAND3_X1  g070(.A1(new_n247_), .A2(new_n248_), .A3(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT80), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n272_), .B(new_n273_), .C1(new_n271_), .C2(new_n247_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT31), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT79), .ZN(new_n276_));
  INV_X1    g075(.A(G113gat), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n277_), .A2(G120gat), .ZN(new_n278_));
  INV_X1    g077(.A(G120gat), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n279_), .A2(G113gat), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT78), .B1(new_n278_), .B2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n279_), .A2(G113gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n277_), .A2(G120gat), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT78), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n282_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G127gat), .B(G134gat), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  AND3_X1   g086(.A1(new_n281_), .A2(new_n285_), .A3(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n287_), .B1(new_n281_), .B2(new_n285_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n276_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n281_), .A2(new_n287_), .A3(new_n285_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT79), .ZN(new_n292_));
  AND2_X1   g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n275_), .B(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(G155gat), .ZN(new_n296_));
  INV_X1    g095(.A(G162gat), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n296_), .A2(new_n297_), .A3(KEYINPUT81), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT81), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n299_), .B1(G155gat), .B2(G162gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G155gat), .A2(G162gat), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n298_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT82), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n298_), .A2(new_n300_), .A3(KEYINPUT82), .A4(new_n301_), .ZN(new_n305_));
  OR3_X1    g104(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G141gat), .A2(G148gat), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT2), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n310_));
  OAI21_X1  g109(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n311_));
  NAND4_X1  g110(.A1(new_n306_), .A2(new_n309_), .A3(new_n310_), .A4(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n304_), .A2(new_n305_), .A3(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(G141gat), .ZN(new_n314_));
  INV_X1    g113(.A(G148gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n301_), .B(KEYINPUT1), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n298_), .A2(new_n300_), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n316_), .B(new_n307_), .C1(new_n317_), .C2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n313_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT29), .ZN(new_n321_));
  INV_X1    g120(.A(G228gat), .ZN(new_n322_));
  INV_X1    g121(.A(G233gat), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(G197gat), .A2(G204gat), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT83), .B(G204gat), .ZN(new_n328_));
  INV_X1    g127(.A(G197gat), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n327_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT21), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  XOR2_X1   g131(.A(G211gat), .B(G218gat), .Z(new_n333_));
  INV_X1    g132(.A(G204gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(KEYINPUT83), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT83), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(G204gat), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n335_), .A2(new_n337_), .A3(new_n329_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n331_), .B1(G197gat), .B2(G204gat), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n333_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n332_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n335_), .A2(new_n337_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n326_), .B1(new_n342_), .B2(G197gat), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT84), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n333_), .A2(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G211gat), .B(G218gat), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n331_), .B1(new_n346_), .B2(KEYINPUT84), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n343_), .A2(new_n345_), .A3(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n341_), .A2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n321_), .A2(new_n325_), .A3(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT85), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n321_), .A2(KEYINPUT85), .A3(new_n325_), .A4(new_n349_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT86), .ZN(new_n354_));
  AND3_X1   g153(.A1(new_n341_), .A2(new_n354_), .A3(new_n348_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n354_), .B1(new_n341_), .B2(new_n348_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n321_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  AOI22_X1  g156(.A1(new_n352_), .A2(new_n353_), .B1(new_n357_), .B2(new_n324_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT87), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G78gat), .B(G106gat), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n362_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT88), .B1(new_n361_), .B2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n352_), .A2(new_n353_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n357_), .A2(new_n324_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT87), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT88), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n368_), .A2(new_n369_), .A3(new_n362_), .A4(new_n360_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n367_), .A2(new_n362_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n320_), .A2(KEYINPUT29), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT28), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G22gat), .B(G50gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n371_), .A2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n364_), .A2(new_n370_), .A3(new_n376_), .ZN(new_n377_));
  AND2_X1   g176(.A1(new_n367_), .A2(new_n362_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n375_), .B1(new_n378_), .B2(new_n371_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n377_), .A2(new_n379_), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n345_), .A2(new_n347_), .ZN(new_n381_));
  AOI22_X1  g180(.A1(new_n381_), .A2(new_n343_), .B1(new_n332_), .B2(new_n340_), .ZN(new_n382_));
  AND3_X1   g181(.A1(new_n263_), .A2(new_n268_), .A3(new_n265_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n258_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n267_), .A2(KEYINPUT89), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT89), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n386_), .A2(G169gat), .A3(G176gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n385_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(G176gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT22), .B(G169gat), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n388_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n259_), .B1(new_n252_), .B2(new_n254_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  AOI22_X1  g192(.A1(new_n383_), .A2(new_n384_), .B1(new_n391_), .B2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n382_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n349_), .A2(new_n270_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G226gat), .A2(G233gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(KEYINPUT19), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n395_), .A2(new_n396_), .A3(KEYINPUT20), .A4(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT20), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n263_), .A2(new_n268_), .A3(new_n265_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n390_), .A2(new_n389_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n403_), .A2(new_n385_), .A3(new_n387_), .ZN(new_n404_));
  OAI22_X1  g203(.A1(new_n402_), .A2(new_n258_), .B1(new_n404_), .B2(new_n392_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n401_), .B1(new_n349_), .B2(new_n405_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n341_), .A2(new_n348_), .A3(new_n260_), .A4(new_n269_), .ZN(new_n407_));
  AOI211_X1 g206(.A(KEYINPUT90), .B(new_n399_), .C1(new_n406_), .C2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT90), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n407_), .B(KEYINPUT20), .C1(new_n382_), .C2(new_n394_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n409_), .B1(new_n410_), .B2(new_n398_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n400_), .B1(new_n408_), .B2(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G8gat), .B(G36gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(KEYINPUT18), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G64gat), .B(G92gat), .ZN(new_n415_));
  XOR2_X1   g214(.A(new_n414_), .B(new_n415_), .Z(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n412_), .A2(new_n417_), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n416_), .B(new_n400_), .C1(new_n408_), .C2(new_n411_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n290_), .A2(new_n320_), .A3(new_n292_), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n313_), .B(new_n319_), .C1(new_n288_), .C2(new_n289_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n420_), .A2(KEYINPUT4), .A3(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G225gat), .A2(G233gat), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT4), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n290_), .A2(new_n320_), .A3(new_n292_), .A4(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n422_), .A2(new_n423_), .A3(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G1gat), .B(G29gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(G85gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(KEYINPUT0), .B(G57gat), .ZN(new_n429_));
  XOR2_X1   g228(.A(new_n428_), .B(new_n429_), .Z(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n423_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n420_), .A2(new_n421_), .A3(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n426_), .A2(new_n431_), .A3(new_n433_), .ZN(new_n434_));
  AND3_X1   g233(.A1(new_n418_), .A2(new_n419_), .A3(new_n434_), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n422_), .A2(KEYINPUT91), .A3(new_n432_), .A4(new_n425_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n420_), .A2(new_n421_), .A3(new_n423_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT33), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT91), .ZN(new_n441_));
  AND3_X1   g240(.A1(new_n420_), .A2(KEYINPUT4), .A3(new_n421_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n425_), .A2(new_n432_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n441_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n439_), .A2(new_n440_), .A3(new_n430_), .A4(new_n444_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n444_), .A2(new_n430_), .A3(new_n437_), .A4(new_n436_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(KEYINPUT33), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n435_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT92), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n416_), .A2(KEYINPUT32), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n349_), .A2(KEYINPUT86), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n341_), .A2(new_n354_), .A3(new_n348_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n453_), .A2(new_n454_), .A3(new_n394_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT93), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(new_n456_), .A3(KEYINPUT20), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(new_n396_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n456_), .B1(new_n455_), .B2(KEYINPUT20), .ZN(new_n459_));
  OAI211_X1 g258(.A(KEYINPUT94), .B(new_n398_), .C1(new_n458_), .C2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n406_), .A2(new_n399_), .A3(new_n407_), .ZN(new_n462_));
  AND2_X1   g261(.A1(new_n462_), .A2(KEYINPUT94), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n455_), .A2(KEYINPUT20), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT93), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n465_), .A2(new_n396_), .A3(new_n457_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n463_), .B1(new_n466_), .B2(new_n398_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n452_), .B1(new_n461_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n444_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n431_), .B1(new_n469_), .B2(new_n438_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n412_), .ZN(new_n471_));
  AOI22_X1  g270(.A1(new_n470_), .A2(new_n446_), .B1(new_n471_), .B2(new_n451_), .ZN(new_n472_));
  AOI22_X1  g271(.A1(new_n449_), .A2(new_n450_), .B1(new_n468_), .B2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n435_), .A2(new_n448_), .A3(KEYINPUT92), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n380_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n470_), .A2(new_n446_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n476_), .B1(new_n377_), .B2(new_n379_), .ZN(new_n477_));
  AOI21_X1  g276(.A(KEYINPUT27), .B1(new_n418_), .B2(new_n419_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n416_), .B(KEYINPUT95), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n479_), .B1(new_n461_), .B2(new_n467_), .ZN(new_n480_));
  AND2_X1   g279(.A1(new_n419_), .A2(KEYINPUT27), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n478_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  AND2_X1   g281(.A1(new_n477_), .A2(new_n482_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n295_), .B1(new_n475_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n476_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n380_), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n294_), .A2(new_n485_), .A3(new_n486_), .A4(new_n482_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n239_), .B1(new_n484_), .B2(new_n487_), .ZN(new_n488_));
  XOR2_X1   g287(.A(G127gat), .B(G155gat), .Z(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT16), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G183gat), .B(G211gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT17), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G231gat), .A2(G233gat), .ZN(new_n494_));
  XOR2_X1   g293(.A(new_n494_), .B(KEYINPUT71), .Z(new_n495_));
  XNOR2_X1  g294(.A(new_n213_), .B(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G71gat), .B(G78gat), .ZN(new_n497_));
  INV_X1    g296(.A(G64gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(G57gat), .ZN(new_n499_));
  INV_X1    g298(.A(G57gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(G64gat), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n497_), .A2(KEYINPUT11), .A3(new_n499_), .A4(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT67), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n499_), .A2(new_n501_), .A3(KEYINPUT11), .ZN(new_n504_));
  INV_X1    g303(.A(G78gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(G71gat), .ZN(new_n506_));
  INV_X1    g305(.A(G71gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(G78gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n504_), .A2(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(KEYINPUT11), .B1(new_n499_), .B2(new_n501_), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n502_), .B(new_n503_), .C1(new_n510_), .C2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT11), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n500_), .A2(G64gat), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n498_), .A2(G57gat), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n514_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n517_), .A2(new_n504_), .A3(new_n509_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n503_), .B1(new_n518_), .B2(new_n502_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n513_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n496_), .A2(new_n520_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n502_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT67), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(new_n512_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n214_), .A2(new_n495_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n495_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n213_), .A2(new_n526_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n524_), .B1(new_n525_), .B2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n493_), .A2(new_n521_), .A3(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n496_), .A2(KEYINPUT72), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT72), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n531_), .B1(new_n525_), .B2(new_n527_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n522_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n530_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT17), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n492_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n533_), .B1(new_n530_), .B2(new_n532_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n529_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT73), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  OAI211_X1 g340(.A(new_n529_), .B(KEYINPUT73), .C1(new_n537_), .C2(new_n538_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G232gat), .A2(G233gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT34), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT64), .ZN(new_n546_));
  NAND2_X1  g345(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n546_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  OR2_X1    g349(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n551_), .A2(KEYINPUT64), .A3(new_n547_), .ZN(new_n552_));
  AOI21_X1  g351(.A(G106gat), .B1(new_n550_), .B2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G99gat), .A2(G106gat), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(KEYINPUT6), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT6), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n556_), .A2(G99gat), .A3(G106gat), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(G85gat), .ZN(new_n559_));
  INV_X1    g358(.A(G92gat), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G85gat), .A2(G92gat), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n561_), .A2(KEYINPUT9), .A3(new_n562_), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n562_), .A2(KEYINPUT9), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n558_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  OR3_X1    g364(.A1(new_n553_), .A2(new_n565_), .A3(KEYINPUT68), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT7), .ZN(new_n567_));
  INV_X1    g366(.A(G99gat), .ZN(new_n568_));
  INV_X1    g367(.A(G106gat), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n567_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT65), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  OAI21_X1  g371(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n567_), .A2(new_n568_), .A3(new_n569_), .A4(KEYINPUT65), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n572_), .A2(new_n558_), .A3(new_n573_), .A4(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n561_), .A2(new_n562_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT66), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n576_), .B1(new_n577_), .B2(KEYINPUT8), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n575_), .A2(new_n578_), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n577_), .A2(KEYINPUT8), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n575_), .A2(new_n578_), .A3(new_n580_), .ZN(new_n583_));
  OAI21_X1  g382(.A(KEYINPUT68), .B1(new_n553_), .B2(new_n565_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n566_), .A2(new_n582_), .A3(new_n583_), .A4(new_n584_), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n230_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n553_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n565_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n582_), .A2(new_n589_), .A3(new_n583_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n590_), .A2(new_n224_), .ZN(new_n591_));
  OAI211_X1 g390(.A(KEYINPUT35), .B(new_n545_), .C1(new_n586_), .C2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G190gat), .B(G218gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G134gat), .B(G162gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n595_), .A2(KEYINPUT36), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT35), .ZN(new_n597_));
  INV_X1    g396(.A(new_n545_), .ZN(new_n598_));
  AOI22_X1  g397(.A1(new_n230_), .A2(new_n585_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n598_), .A2(new_n597_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n591_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n599_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n592_), .A2(new_n596_), .A3(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n595_), .B(KEYINPUT36), .Z(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n607_), .B1(new_n592_), .B2(new_n603_), .ZN(new_n608_));
  OAI21_X1  g407(.A(KEYINPUT37), .B1(new_n605_), .B2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n592_), .A2(new_n603_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(new_n606_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT37), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n611_), .A2(new_n612_), .A3(new_n604_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n543_), .B1(new_n609_), .B2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n590_), .A2(new_n520_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT12), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n533_), .A2(KEYINPUT12), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  AOI22_X1  g417(.A1(new_n615_), .A2(new_n616_), .B1(new_n585_), .B2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(G230gat), .A2(G233gat), .ZN(new_n620_));
  OAI211_X1 g419(.A(KEYINPUT69), .B(new_n620_), .C1(new_n590_), .C2(new_n520_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  AND3_X1   g421(.A1(new_n575_), .A2(new_n580_), .A3(new_n578_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n580_), .B1(new_n575_), .B2(new_n578_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n625_), .A2(new_n524_), .A3(new_n589_), .ZN(new_n626_));
  AOI21_X1  g425(.A(KEYINPUT69), .B1(new_n626_), .B2(new_n620_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n619_), .B1(new_n622_), .B2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n615_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n620_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n628_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(G120gat), .B(G148gat), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT5), .ZN(new_n635_));
  XNOR2_X1  g434(.A(G176gat), .B(G204gat), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n635_), .B(new_n636_), .Z(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n633_), .A2(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n632_), .A2(new_n637_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(KEYINPUT13), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT13), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n643_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n644_));
  AND3_X1   g443(.A1(new_n614_), .A2(new_n642_), .A3(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT74), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n488_), .A2(new_n646_), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n476_), .A2(KEYINPUT96), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n476_), .A2(KEYINPUT96), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NOR3_X1   g450(.A1(new_n647_), .A2(G1gat), .A3(new_n651_), .ZN(new_n652_));
  XOR2_X1   g451(.A(KEYINPUT97), .B(KEYINPUT38), .Z(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n652_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n239_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n605_), .A2(new_n608_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT98), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n658_), .B1(new_n484_), .B2(new_n487_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n539_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n642_), .A2(new_n644_), .ZN(new_n661_));
  AND4_X1   g460(.A1(new_n656_), .A2(new_n659_), .A3(new_n660_), .A4(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(new_n476_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n653_), .B1(new_n663_), .B2(G1gat), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n655_), .B1(new_n664_), .B2(new_n652_), .ZN(G1324gat));
  INV_X1    g464(.A(new_n647_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n482_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n666_), .A2(new_n209_), .A3(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n662_), .A2(new_n667_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(G8gat), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n670_), .A2(KEYINPUT39), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n670_), .A2(KEYINPUT39), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n668_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT40), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  OAI211_X1 g474(.A(KEYINPUT40), .B(new_n668_), .C1(new_n671_), .C2(new_n672_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1325gat));
  NAND3_X1  g476(.A1(new_n666_), .A2(new_n241_), .A3(new_n294_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n662_), .A2(new_n294_), .ZN(new_n679_));
  AND3_X1   g478(.A1(new_n679_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n680_));
  AOI21_X1  g479(.A(KEYINPUT41), .B1(new_n679_), .B2(G15gat), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n678_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT99), .ZN(G1326gat));
  INV_X1    g482(.A(G22gat), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n684_), .B1(new_n662_), .B2(new_n380_), .ZN(new_n685_));
  XOR2_X1   g484(.A(new_n685_), .B(KEYINPUT42), .Z(new_n686_));
  NAND2_X1  g485(.A1(new_n380_), .A2(new_n684_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT100), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n686_), .B1(new_n647_), .B2(new_n688_), .ZN(G1327gat));
  INV_X1    g488(.A(new_n661_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n657_), .A2(new_n543_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n488_), .A2(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(G29gat), .B1(new_n693_), .B2(new_n476_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n543_), .ZN(new_n695_));
  NOR3_X1   g494(.A1(new_n690_), .A2(new_n239_), .A3(new_n695_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n446_), .B(new_n440_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n418_), .A2(new_n419_), .A3(new_n434_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n450_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n468_), .A2(new_n472_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n699_), .A2(new_n700_), .A3(new_n474_), .ZN(new_n701_));
  AOI22_X1  g500(.A1(new_n701_), .A2(new_n486_), .B1(new_n477_), .B2(new_n482_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n487_), .B1(new_n702_), .B2(new_n294_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT43), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n609_), .A2(new_n613_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n703_), .A2(new_n704_), .A3(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n704_), .B1(new_n703_), .B2(new_n706_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n696_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT44), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  OAI211_X1 g510(.A(KEYINPUT44), .B(new_n696_), .C1(new_n707_), .C2(new_n708_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n650_), .A2(G29gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n694_), .B1(new_n713_), .B2(new_n714_), .ZN(G1328gat));
  INV_X1    g514(.A(KEYINPUT46), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n716_), .A2(KEYINPUT102), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n711_), .A2(new_n667_), .A3(new_n712_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(G36gat), .ZN(new_n719_));
  INV_X1    g518(.A(G36gat), .ZN(new_n720_));
  OR2_X1    g519(.A1(new_n667_), .A2(KEYINPUT101), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n667_), .A2(KEYINPUT101), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n693_), .A2(new_n720_), .A3(new_n723_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT45), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n717_), .B1(new_n719_), .B2(new_n725_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n716_), .A2(KEYINPUT102), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n726_), .B(new_n727_), .ZN(G1329gat));
  AOI21_X1  g527(.A(G43gat), .B1(new_n693_), .B2(new_n294_), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT103), .Z(new_n730_));
  NAND3_X1  g529(.A1(new_n713_), .A2(G43gat), .A3(new_n294_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(KEYINPUT47), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT47), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n730_), .A2(new_n731_), .A3(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(G1330gat));
  INV_X1    g535(.A(G50gat), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n693_), .A2(new_n737_), .A3(new_n380_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n711_), .A2(new_n380_), .A3(new_n712_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n739_), .A2(KEYINPUT104), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT104), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n711_), .A2(new_n741_), .A3(new_n380_), .A4(new_n712_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(G50gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n738_), .B1(new_n740_), .B2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT105), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT105), .ZN(new_n746_));
  OAI211_X1 g545(.A(new_n746_), .B(new_n738_), .C1(new_n740_), .C2(new_n743_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n747_), .ZN(G1331gat));
  AOI21_X1  g547(.A(new_n656_), .B1(new_n484_), .B2(new_n487_), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n749_), .A2(new_n614_), .A3(new_n690_), .ZN(new_n750_));
  AOI21_X1  g549(.A(G57gat), .B1(new_n750_), .B2(new_n650_), .ZN(new_n751_));
  AND4_X1   g550(.A1(new_n239_), .A2(new_n659_), .A3(new_n695_), .A4(new_n690_), .ZN(new_n752_));
  XOR2_X1   g551(.A(KEYINPUT106), .B(G57gat), .Z(new_n753_));
  NOR2_X1   g552(.A1(new_n485_), .A2(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n751_), .B1(new_n752_), .B2(new_n754_), .ZN(G1332gat));
  AOI21_X1  g554(.A(new_n498_), .B1(new_n752_), .B2(new_n723_), .ZN(new_n756_));
  XOR2_X1   g555(.A(new_n756_), .B(KEYINPUT48), .Z(new_n757_));
  NAND3_X1  g556(.A1(new_n750_), .A2(new_n498_), .A3(new_n723_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(G1333gat));
  NAND3_X1  g558(.A1(new_n750_), .A2(new_n507_), .A3(new_n294_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n752_), .A2(new_n294_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(G71gat), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n762_), .A2(KEYINPUT49), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n762_), .A2(KEYINPUT49), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n760_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT107), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT107), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n767_), .B(new_n760_), .C1(new_n763_), .C2(new_n764_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(G1334gat));
  NAND3_X1  g568(.A1(new_n750_), .A2(new_n505_), .A3(new_n380_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n752_), .A2(new_n380_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(G78gat), .ZN(new_n772_));
  XNOR2_X1  g571(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n772_), .A2(new_n773_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n770_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(KEYINPUT109), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT109), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n778_), .B(new_n770_), .C1(new_n774_), .C2(new_n775_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(G1335gat));
  AND4_X1   g579(.A1(new_n543_), .A2(new_n749_), .A3(new_n657_), .A4(new_n690_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n781_), .A2(new_n559_), .A3(new_n650_), .ZN(new_n782_));
  OR2_X1    g581(.A1(new_n707_), .A2(new_n708_), .ZN(new_n783_));
  NOR3_X1   g582(.A1(new_n661_), .A2(new_n656_), .A3(new_n695_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT110), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n783_), .A2(new_n785_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n786_), .A2(new_n476_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n782_), .B1(new_n787_), .B2(new_n559_), .ZN(G1336gat));
  AOI21_X1  g587(.A(G92gat), .B1(new_n781_), .B2(new_n667_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT111), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n560_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n786_), .B2(new_n791_), .ZN(G1337gat));
  NAND2_X1  g591(.A1(new_n786_), .A2(new_n294_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n295_), .B1(new_n552_), .B2(new_n550_), .ZN(new_n794_));
  AOI22_X1  g593(.A1(new_n793_), .A2(G99gat), .B1(new_n781_), .B2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT51), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n796_), .A2(KEYINPUT112), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n795_), .B(new_n798_), .ZN(G1338gat));
  NAND3_X1  g598(.A1(new_n781_), .A2(new_n569_), .A3(new_n380_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n783_), .A2(new_n380_), .A3(new_n785_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n802_));
  AND3_X1   g601(.A1(new_n801_), .A2(new_n802_), .A3(G106gat), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n802_), .B1(new_n801_), .B2(G106gat), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n800_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n805_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g605(.A(KEYINPUT113), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT54), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n645_), .A2(new_n807_), .A3(new_n808_), .A4(new_n239_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n614_), .A2(new_n642_), .A3(new_n239_), .A4(new_n644_), .ZN(new_n810_));
  OAI21_X1  g609(.A(KEYINPUT113), .B1(new_n810_), .B2(KEYINPUT54), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(KEYINPUT54), .ZN(new_n812_));
  AND3_X1   g611(.A1(new_n809_), .A2(new_n811_), .A3(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT118), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n814_), .A2(KEYINPUT58), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n628_), .A2(new_n816_), .ZN(new_n817_));
  OAI211_X1 g616(.A(KEYINPUT55), .B(new_n619_), .C1(new_n622_), .C2(new_n627_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n619_), .A2(new_n626_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n630_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n817_), .A2(new_n818_), .A3(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n637_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT56), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n821_), .A2(KEYINPUT56), .A3(new_n637_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n236_), .A2(new_n237_), .A3(new_n204_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n225_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n206_), .B1(new_n828_), .B2(new_n232_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n214_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n223_), .A2(new_n233_), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n829_), .B(new_n205_), .C1(new_n830_), .C2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n827_), .A2(new_n832_), .A3(KEYINPUT116), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n827_), .A2(new_n832_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT116), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n640_), .B1(new_n833_), .B2(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n815_), .B1(new_n826_), .B2(new_n837_), .ZN(new_n838_));
  AOI22_X1  g637(.A1(new_n628_), .A2(new_n816_), .B1(new_n630_), .B2(new_n819_), .ZN(new_n839_));
  AOI211_X1 g638(.A(new_n823_), .B(new_n638_), .C1(new_n839_), .C2(new_n818_), .ZN(new_n840_));
  AOI21_X1  g639(.A(KEYINPUT56), .B1(new_n821_), .B2(new_n637_), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n815_), .B(new_n837_), .C1(new_n840_), .C2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n706_), .B1(new_n838_), .B2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT119), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  XOR2_X1   g645(.A(KEYINPUT117), .B(KEYINPUT57), .Z(new_n847_));
  AND2_X1   g646(.A1(new_n836_), .A2(new_n833_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n641_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT115), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n821_), .A2(new_n850_), .A3(KEYINPUT56), .A4(new_n637_), .ZN(new_n851_));
  OAI21_X1  g650(.A(KEYINPUT114), .B1(new_n640_), .B2(new_n239_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT114), .ZN(new_n853_));
  OAI221_X1 g652(.A(new_n853_), .B1(new_n238_), .B2(new_n235_), .C1(new_n632_), .C2(new_n637_), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n851_), .A2(new_n852_), .A3(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n824_), .A2(KEYINPUT115), .A3(new_n825_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n849_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n847_), .B1(new_n857_), .B2(new_n657_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n657_), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n840_), .A2(new_n841_), .A3(new_n850_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n851_), .A2(new_n852_), .A3(new_n854_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  OAI211_X1 g661(.A(KEYINPUT57), .B(new_n859_), .C1(new_n862_), .C2(new_n849_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n837_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n815_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n842_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n867_), .A2(KEYINPUT119), .A3(new_n706_), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n846_), .A2(new_n858_), .A3(new_n863_), .A4(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n813_), .B1(new_n869_), .B2(new_n539_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n295_), .A2(new_n651_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n667_), .A2(new_n380_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n870_), .A2(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(G113gat), .B1(new_n874_), .B2(new_n656_), .ZN(new_n875_));
  AND2_X1   g674(.A1(new_n863_), .A2(new_n858_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n844_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n813_), .B1(new_n877_), .B2(new_n543_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n873_), .ZN(new_n879_));
  XOR2_X1   g678(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  OR2_X1    g680(.A1(new_n878_), .A2(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(KEYINPUT119), .B1(new_n867_), .B2(new_n706_), .ZN(new_n883_));
  AOI211_X1 g682(.A(new_n845_), .B(new_n705_), .C1(new_n866_), .C2(new_n842_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n660_), .B1(new_n876_), .B2(new_n885_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n879_), .B1(new_n886_), .B2(new_n813_), .ZN(new_n887_));
  AOI21_X1  g686(.A(KEYINPUT120), .B1(new_n887_), .B2(KEYINPUT59), .ZN(new_n888_));
  OAI211_X1 g687(.A(KEYINPUT120), .B(KEYINPUT59), .C1(new_n870_), .C2(new_n873_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n882_), .B1(new_n888_), .B2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(KEYINPUT122), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT122), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n893_), .B(new_n882_), .C1(new_n888_), .C2(new_n890_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n894_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n239_), .A2(new_n277_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n875_), .B1(new_n895_), .B2(new_n896_), .ZN(G1340gat));
  OAI21_X1  g696(.A(new_n279_), .B1(new_n661_), .B2(KEYINPUT60), .ZN(new_n898_));
  OAI211_X1 g697(.A(new_n874_), .B(new_n898_), .C1(KEYINPUT60), .C2(new_n279_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n690_), .B1(new_n878_), .B2(new_n881_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT120), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT59), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n874_), .B2(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n900_), .B1(new_n903_), .B2(new_n889_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n899_), .B1(new_n904_), .B2(new_n279_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(KEYINPUT123), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT123), .ZN(new_n907_));
  OAI211_X1 g706(.A(new_n907_), .B(new_n899_), .C1(new_n904_), .C2(new_n279_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n906_), .A2(new_n908_), .ZN(G1341gat));
  AOI21_X1  g708(.A(G127gat), .B1(new_n874_), .B2(new_n695_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n660_), .A2(G127gat), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n910_), .B1(new_n895_), .B2(new_n912_), .ZN(G1342gat));
  AOI21_X1  g712(.A(G134gat), .B1(new_n874_), .B2(new_n658_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n706_), .A2(G134gat), .ZN(new_n915_));
  XOR2_X1   g714(.A(new_n915_), .B(KEYINPUT124), .Z(new_n916_));
  AOI21_X1  g715(.A(new_n914_), .B1(new_n895_), .B2(new_n916_), .ZN(G1343gat));
  NOR2_X1   g716(.A1(new_n870_), .A2(new_n294_), .ZN(new_n918_));
  NOR3_X1   g717(.A1(new_n723_), .A2(new_n486_), .A3(new_n651_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n920_), .A2(new_n239_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(new_n314_), .ZN(G1344gat));
  NOR2_X1   g721(.A1(new_n920_), .A2(new_n661_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(new_n315_), .ZN(G1345gat));
  NOR2_X1   g723(.A1(new_n920_), .A2(new_n543_), .ZN(new_n925_));
  XOR2_X1   g724(.A(KEYINPUT61), .B(G155gat), .Z(new_n926_));
  XNOR2_X1  g725(.A(new_n925_), .B(new_n926_), .ZN(G1346gat));
  OAI21_X1  g726(.A(G162gat), .B1(new_n920_), .B2(new_n705_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n658_), .A2(new_n297_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n920_), .B2(new_n929_), .ZN(G1347gat));
  NAND3_X1  g729(.A1(new_n723_), .A2(new_n294_), .A3(new_n651_), .ZN(new_n931_));
  INV_X1    g730(.A(new_n931_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n695_), .B1(new_n876_), .B2(new_n844_), .ZN(new_n933_));
  OAI211_X1 g732(.A(new_n486_), .B(new_n932_), .C1(new_n933_), .C2(new_n813_), .ZN(new_n934_));
  OAI21_X1  g733(.A(G169gat), .B1(new_n934_), .B2(new_n239_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(KEYINPUT62), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n656_), .A2(new_n390_), .ZN(new_n937_));
  XOR2_X1   g736(.A(new_n937_), .B(KEYINPUT125), .Z(new_n938_));
  OAI21_X1  g737(.A(new_n936_), .B1(new_n934_), .B2(new_n938_), .ZN(G1348gat));
  INV_X1    g738(.A(new_n934_), .ZN(new_n940_));
  AOI21_X1  g739(.A(G176gat), .B1(new_n940_), .B2(new_n690_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n870_), .A2(new_n380_), .ZN(new_n942_));
  NOR3_X1   g741(.A1(new_n931_), .A2(new_n389_), .A3(new_n661_), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n941_), .B1(new_n942_), .B2(new_n943_), .ZN(G1349gat));
  NOR3_X1   g743(.A1(new_n934_), .A2(new_n261_), .A3(new_n539_), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n942_), .A2(new_n695_), .A3(new_n932_), .ZN(new_n946_));
  INV_X1    g745(.A(G183gat), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n945_), .B1(new_n946_), .B2(new_n947_), .ZN(G1350gat));
  OAI21_X1  g747(.A(G190gat), .B1(new_n934_), .B2(new_n705_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n658_), .A2(new_n262_), .ZN(new_n950_));
  XOR2_X1   g749(.A(new_n950_), .B(KEYINPUT126), .Z(new_n951_));
  OAI21_X1  g750(.A(new_n949_), .B1(new_n934_), .B2(new_n951_), .ZN(G1351gat));
  NAND3_X1  g751(.A1(new_n918_), .A2(new_n477_), .A3(new_n723_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n953_), .A2(new_n239_), .ZN(new_n954_));
  XNOR2_X1  g753(.A(new_n954_), .B(new_n329_), .ZN(G1352gat));
  NOR2_X1   g754(.A1(new_n953_), .A2(new_n661_), .ZN(new_n956_));
  NOR2_X1   g755(.A1(new_n956_), .A2(G204gat), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n957_), .B1(new_n342_), .B2(new_n956_), .ZN(G1353gat));
  NAND2_X1  g757(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n660_), .A2(new_n959_), .ZN(new_n960_));
  XNOR2_X1  g759(.A(new_n960_), .B(KEYINPUT127), .ZN(new_n961_));
  NOR2_X1   g760(.A1(new_n953_), .A2(new_n961_), .ZN(new_n962_));
  NOR2_X1   g761(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n963_));
  XNOR2_X1  g762(.A(new_n962_), .B(new_n963_), .ZN(G1354gat));
  OAI21_X1  g763(.A(G218gat), .B1(new_n953_), .B2(new_n705_), .ZN(new_n965_));
  INV_X1    g764(.A(G218gat), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n658_), .A2(new_n966_), .ZN(new_n967_));
  OAI21_X1  g766(.A(new_n965_), .B1(new_n953_), .B2(new_n967_), .ZN(G1355gat));
endmodule


