//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 0 1 0 1 0 1 1 1 0 1 1 0 1 0 0 1 0 0 0 1 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n711_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n843_,
    new_n844_, new_n845_, new_n847_, new_n848_, new_n849_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n866_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n902_, new_n903_, new_n904_, new_n906_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n914_, new_n915_;
  INV_X1    g000(.A(G141gat), .ZN(new_n202_));
  INV_X1    g001(.A(G148gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G141gat), .A2(G148gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  XOR2_X1   g006(.A(G155gat), .B(G162gat), .Z(new_n208_));
  INV_X1    g007(.A(KEYINPUT1), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n207_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT82), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT3), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n213_), .A2(new_n202_), .A3(new_n203_), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n215_));
  INV_X1    g014(.A(new_n205_), .ZN(new_n216_));
  OAI211_X1 g015(.A(new_n214_), .B(new_n215_), .C1(KEYINPUT2), .C2(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n208_), .B1(new_n212_), .B2(new_n217_), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n210_), .B1(new_n218_), .B2(KEYINPUT83), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT83), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n220_), .B(new_n208_), .C1(new_n212_), .C2(new_n217_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n219_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT79), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G127gat), .B(G134gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G113gat), .B(G120gat), .ZN(new_n225_));
  AND2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n224_), .A2(new_n225_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n223_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT79), .B1(new_n224_), .B2(new_n225_), .ZN(new_n229_));
  AND2_X1   g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n222_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT91), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G225gat), .A2(G233gat), .ZN(new_n233_));
  XOR2_X1   g032(.A(new_n233_), .B(KEYINPUT92), .Z(new_n234_));
  OAI211_X1 g033(.A(new_n219_), .B(new_n221_), .C1(new_n227_), .C2(new_n226_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT91), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n222_), .A2(new_n236_), .A3(new_n230_), .ZN(new_n237_));
  NAND4_X1  g036(.A1(new_n232_), .A2(new_n234_), .A3(new_n235_), .A4(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G1gat), .B(G29gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(G85gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT0), .B(G57gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n238_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n237_), .A2(new_n235_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n236_), .B1(new_n222_), .B2(new_n230_), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT4), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT4), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n231_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n243_), .B1(new_n249_), .B2(new_n233_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT90), .ZN(new_n251_));
  OAI21_X1  g050(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(G169gat), .ZN(new_n254_));
  INV_X1    g053(.A(G176gat), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n253_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G183gat), .A2(G190gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT23), .ZN(new_n258_));
  OR3_X1    g057(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n259_));
  AND3_X1   g058(.A1(new_n256_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT25), .B(G183gat), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  XOR2_X1   g061(.A(KEYINPUT26), .B(G190gat), .Z(new_n263_));
  OR2_X1    g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n260_), .A2(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n258_), .B1(G183gat), .B2(G190gat), .ZN(new_n266_));
  NOR2_X1   g065(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(G169gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n266_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n265_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G211gat), .B(G218gat), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT21), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(G197gat), .ZN(new_n274_));
  OAI21_X1  g073(.A(KEYINPUT85), .B1(new_n274_), .B2(G204gat), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT85), .ZN(new_n276_));
  INV_X1    g075(.A(G204gat), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n276_), .A2(new_n277_), .A3(G197gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n274_), .A2(G204gat), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n275_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n273_), .A2(new_n280_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n274_), .A2(G204gat), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n277_), .A2(G197gat), .ZN(new_n283_));
  OAI21_X1  g082(.A(KEYINPUT21), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n275_), .A2(new_n278_), .A3(new_n272_), .A4(new_n279_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT86), .ZN(new_n286_));
  OAI211_X1 g085(.A(new_n284_), .B(new_n271_), .C1(new_n285_), .C2(new_n286_), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n285_), .A2(new_n286_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n281_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n251_), .B1(new_n270_), .B2(new_n289_), .ZN(new_n290_));
  OR2_X1    g089(.A1(new_n287_), .A2(new_n288_), .ZN(new_n291_));
  AOI22_X1  g090(.A1(new_n260_), .A2(new_n264_), .B1(new_n266_), .B2(new_n268_), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n291_), .A2(new_n292_), .A3(KEYINPUT90), .A4(new_n281_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT20), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT26), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n295_), .A2(G190gat), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n261_), .B1(KEYINPUT78), .B2(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n297_), .B1(KEYINPUT78), .B2(new_n263_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n256_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n269_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n294_), .B1(new_n300_), .B2(new_n289_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G226gat), .A2(G233gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT19), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n290_), .A2(new_n293_), .A3(new_n301_), .A4(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n292_), .B1(new_n291_), .B2(new_n281_), .ZN(new_n306_));
  OAI21_X1  g105(.A(KEYINPUT20), .B1(new_n300_), .B2(new_n289_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n303_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n305_), .A2(new_n308_), .ZN(new_n309_));
  XOR2_X1   g108(.A(G8gat), .B(G36gat), .Z(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT18), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G64gat), .B(G92gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n309_), .A2(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n305_), .A2(new_n308_), .A3(new_n313_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n250_), .A2(new_n317_), .ZN(new_n318_));
  NAND4_X1  g117(.A1(new_n232_), .A2(new_n233_), .A3(new_n235_), .A4(new_n237_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(KEYINPUT93), .ZN(new_n320_));
  AND2_X1   g119(.A1(new_n237_), .A2(new_n235_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT93), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n321_), .A2(new_n322_), .A3(new_n233_), .A4(new_n232_), .ZN(new_n323_));
  AND2_X1   g122(.A1(new_n320_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n249_), .A2(new_n234_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n242_), .ZN(new_n326_));
  AND2_X1   g125(.A1(new_n326_), .A2(KEYINPUT33), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n324_), .A2(new_n325_), .A3(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n320_), .A2(new_n323_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n234_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n330_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n331_));
  NOR3_X1   g130(.A1(new_n329_), .A2(new_n331_), .A3(new_n242_), .ZN(new_n332_));
  OAI211_X1 g131(.A(new_n318_), .B(new_n328_), .C1(new_n332_), .C2(KEYINPUT33), .ZN(new_n333_));
  AND2_X1   g132(.A1(new_n313_), .A2(KEYINPUT32), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n309_), .A2(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n291_), .A2(KEYINPUT89), .A3(new_n281_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT89), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n289_), .A2(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n336_), .A2(new_n292_), .A3(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(new_n301_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(new_n303_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT94), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  OR2_X1    g142(.A1(new_n300_), .A2(new_n289_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n270_), .A2(new_n289_), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n344_), .A2(KEYINPUT20), .A3(new_n304_), .A4(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT95), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n306_), .A2(new_n307_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT95), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n348_), .A2(new_n349_), .A3(new_n304_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n347_), .A2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n340_), .A2(KEYINPUT94), .A3(new_n303_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n343_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n335_), .B1(new_n353_), .B2(new_n334_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n326_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n354_), .B1(new_n355_), .B2(new_n332_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n333_), .A2(new_n356_), .ZN(new_n357_));
  XOR2_X1   g156(.A(G78gat), .B(G106gat), .Z(new_n358_));
  INV_X1    g157(.A(G233gat), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n359_), .A2(KEYINPUT84), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n359_), .A2(KEYINPUT84), .ZN(new_n361_));
  OAI21_X1  g160(.A(G228gat), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n222_), .A2(KEYINPUT29), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT88), .ZN(new_n364_));
  AOI22_X1  g163(.A1(new_n363_), .A2(new_n364_), .B1(new_n336_), .B2(new_n338_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT29), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n366_), .B1(new_n219_), .B2(new_n221_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT88), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n362_), .B1(new_n365_), .B2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT87), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n363_), .A2(new_n370_), .A3(new_n289_), .A4(new_n362_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n289_), .A2(new_n362_), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT87), .B1(new_n367_), .B2(new_n372_), .ZN(new_n373_));
  AND2_X1   g172(.A1(new_n371_), .A2(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n358_), .B1(new_n369_), .B2(new_n374_), .ZN(new_n375_));
  OR3_X1    g174(.A1(new_n222_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT28), .B1(new_n222_), .B2(KEYINPUT29), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G22gat), .B(G50gat), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  AND3_X1   g178(.A1(new_n376_), .A2(new_n377_), .A3(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n379_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n363_), .A2(new_n364_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n336_), .A2(new_n338_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n383_), .A2(new_n384_), .A3(new_n368_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n362_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n358_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n371_), .A2(new_n373_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n387_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n390_));
  AND3_X1   g189(.A1(new_n375_), .A2(new_n382_), .A3(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n382_), .B1(new_n375_), .B2(new_n390_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n357_), .A2(new_n393_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n355_), .A2(new_n332_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n353_), .A2(new_n314_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT27), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n316_), .A2(KEYINPUT96), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT96), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n305_), .A2(new_n308_), .A3(new_n399_), .A4(new_n313_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n397_), .B1(new_n398_), .B2(new_n400_), .ZN(new_n401_));
  AOI22_X1  g200(.A1(new_n396_), .A2(new_n401_), .B1(new_n397_), .B2(new_n317_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n382_), .ZN(new_n403_));
  NOR3_X1   g202(.A1(new_n369_), .A2(new_n374_), .A3(new_n358_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n388_), .B1(new_n387_), .B2(new_n389_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n403_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n375_), .A2(new_n382_), .A3(new_n390_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n395_), .A2(new_n402_), .A3(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT97), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT97), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n395_), .A2(new_n402_), .A3(new_n408_), .A4(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n394_), .A2(new_n410_), .A3(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G71gat), .B(G99gat), .ZN(new_n414_));
  INV_X1    g213(.A(G43gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n300_), .B(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G227gat), .A2(G233gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(G15gat), .ZN(new_n419_));
  XOR2_X1   g218(.A(new_n419_), .B(KEYINPUT30), .Z(new_n420_));
  XNOR2_X1  g219(.A(new_n417_), .B(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n230_), .B(KEYINPUT31), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT80), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n422_), .A2(new_n423_), .ZN(new_n425_));
  NOR3_X1   g224(.A1(new_n421_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n426_), .B1(new_n424_), .B2(new_n421_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(KEYINPUT81), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n317_), .A2(new_n397_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n304_), .B1(new_n339_), .B2(new_n301_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n431_), .B(new_n342_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n313_), .B1(new_n432_), .B2(new_n351_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n398_), .A2(new_n400_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT27), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n430_), .B1(new_n433_), .B2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT98), .B1(new_n436_), .B2(new_n408_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT98), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n393_), .A2(new_n402_), .A3(new_n438_), .ZN(new_n439_));
  AND3_X1   g238(.A1(new_n437_), .A2(new_n439_), .A3(new_n427_), .ZN(new_n440_));
  AOI22_X1  g239(.A1(new_n413_), .A2(new_n429_), .B1(new_n440_), .B2(new_n395_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G15gat), .B(G22gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G1gat), .A2(G8gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(KEYINPUT14), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G1gat), .B(G8gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n445_), .B(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G29gat), .B(G36gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G43gat), .B(G50gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  XOR2_X1   g249(.A(new_n447_), .B(new_n450_), .Z(new_n451_));
  NAND2_X1  g250(.A1(G229gat), .A2(G233gat), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n450_), .B(KEYINPUT15), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(new_n447_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n447_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n453_), .B1(new_n456_), .B2(new_n450_), .ZN(new_n457_));
  AOI22_X1  g256(.A1(new_n451_), .A2(new_n453_), .B1(new_n455_), .B2(new_n457_), .ZN(new_n458_));
  XOR2_X1   g257(.A(G113gat), .B(G141gat), .Z(new_n459_));
  XNOR2_X1  g258(.A(G169gat), .B(G197gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n458_), .B(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n441_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT37), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G99gat), .A2(G106gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT6), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT6), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n468_), .A2(G99gat), .A3(G106gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n467_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT9), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n471_), .A2(G85gat), .A3(G92gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G85gat), .B(G92gat), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n470_), .B(new_n472_), .C1(new_n471_), .C2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT10), .B(G99gat), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT65), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(G106gat), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n474_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT66), .ZN(new_n480_));
  OAI22_X1  g279(.A1(new_n480_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(KEYINPUT66), .B(KEYINPUT7), .ZN(new_n482_));
  NOR2_X1   g281(.A1(G99gat), .A2(G106gat), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n481_), .B1(new_n482_), .B2(new_n484_), .ZN(new_n485_));
  AND3_X1   g284(.A1(new_n467_), .A2(new_n469_), .A3(KEYINPUT67), .ZN(new_n486_));
  AOI21_X1  g285(.A(KEYINPUT67), .B1(new_n467_), .B2(new_n469_), .ZN(new_n487_));
  NOR3_X1   g286(.A1(new_n485_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT8), .B1(new_n488_), .B2(new_n473_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n470_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n485_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n473_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT8), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  OR2_X1    g293(.A1(new_n491_), .A2(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n479_), .B1(new_n489_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(new_n450_), .ZN(new_n497_));
  AND2_X1   g296(.A1(new_n470_), .A2(new_n472_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n492_), .A2(KEYINPUT9), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n475_), .B(KEYINPUT65), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n498_), .B(new_n499_), .C1(new_n500_), .C2(G106gat), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT67), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n470_), .A2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n467_), .A2(new_n469_), .A3(KEYINPUT67), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n480_), .A2(KEYINPUT7), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT7), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n506_), .A2(KEYINPUT66), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n483_), .B1(new_n505_), .B2(new_n507_), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n503_), .A2(new_n504_), .A3(new_n508_), .A4(new_n481_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n493_), .B1(new_n509_), .B2(new_n492_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n491_), .A2(new_n494_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n501_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(new_n454_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G232gat), .A2(G233gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT34), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT35), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n497_), .A2(new_n513_), .A3(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT75), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT73), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT73), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n497_), .A2(new_n522_), .A3(new_n513_), .A4(new_n518_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n516_), .A2(new_n517_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n521_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  OAI221_X1 g324(.A(KEYINPUT73), .B1(new_n517_), .B2(new_n516_), .C1(new_n519_), .C2(new_n520_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G190gat), .B(G218gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT74), .ZN(new_n528_));
  XOR2_X1   g327(.A(G134gat), .B(G162gat), .Z(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n530_), .B(KEYINPUT36), .Z(new_n531_));
  NAND3_X1  g330(.A1(new_n525_), .A2(new_n526_), .A3(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT76), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n465_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n532_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n530_), .A2(KEYINPUT36), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n537_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n534_), .B1(new_n535_), .B2(new_n538_), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n525_), .A2(new_n526_), .ZN(new_n540_));
  OAI221_X1 g339(.A(new_n532_), .B1(new_n533_), .B2(new_n465_), .C1(new_n540_), .C2(new_n537_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT12), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G57gat), .B(G64gat), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(KEYINPUT11), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT68), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT11), .ZN(new_n548_));
  INV_X1    g347(.A(G57gat), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n549_), .A2(G64gat), .ZN(new_n550_));
  INV_X1    g349(.A(G64gat), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n551_), .A2(G57gat), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n548_), .B1(new_n550_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(G71gat), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(G78gat), .ZN(new_n555_));
  INV_X1    g354(.A(G78gat), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(G71gat), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n547_), .B1(new_n553_), .B2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n551_), .A2(G57gat), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n549_), .A2(G64gat), .ZN(new_n561_));
  AOI21_X1  g360(.A(KEYINPUT11), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G71gat), .B(G78gat), .ZN(new_n563_));
  NOR3_X1   g362(.A1(new_n562_), .A2(KEYINPUT68), .A3(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n546_), .B1(new_n559_), .B2(new_n564_), .ZN(new_n565_));
  OAI21_X1  g364(.A(KEYINPUT68), .B1(new_n562_), .B2(new_n563_), .ZN(new_n566_));
  OAI211_X1 g365(.A(new_n558_), .B(new_n547_), .C1(new_n545_), .C2(KEYINPUT11), .ZN(new_n567_));
  INV_X1    g366(.A(new_n546_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n566_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n565_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n544_), .B1(new_n496_), .B2(new_n571_), .ZN(new_n572_));
  AND3_X1   g371(.A1(new_n566_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n568_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT69), .ZN(new_n575_));
  NOR3_X1   g374(.A1(new_n573_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(KEYINPUT69), .B1(new_n565_), .B2(new_n569_), .ZN(new_n577_));
  OAI211_X1 g376(.A(KEYINPUT12), .B(new_n512_), .C1(new_n576_), .C2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G230gat), .A2(G233gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT64), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n496_), .A2(new_n571_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n572_), .A2(new_n578_), .A3(new_n581_), .A4(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n496_), .A2(new_n571_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n512_), .A2(new_n570_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n580_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  XOR2_X1   g385(.A(G120gat), .B(G148gat), .Z(new_n587_));
  XNOR2_X1  g386(.A(G176gat), .B(G204gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n583_), .A2(new_n586_), .A3(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n591_), .B(KEYINPUT71), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n594_), .B1(new_n583_), .B2(new_n586_), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(KEYINPUT72), .B(KEYINPUT13), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT72), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n596_), .B1(new_n599_), .B2(KEYINPUT13), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(G231gat), .A2(G233gat), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n447_), .B(new_n603_), .Z(new_n604_));
  OR2_X1    g403(.A1(new_n604_), .A2(new_n571_), .ZN(new_n605_));
  XOR2_X1   g404(.A(G127gat), .B(G155gat), .Z(new_n606_));
  XNOR2_X1  g405(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G183gat), .B(G211gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(KEYINPUT17), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n604_), .A2(new_n571_), .ZN(new_n612_));
  OR2_X1    g411(.A1(new_n610_), .A2(KEYINPUT17), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n605_), .A2(new_n611_), .A3(new_n612_), .A4(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n575_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n565_), .A2(KEYINPUT69), .A3(new_n569_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n611_), .B1(new_n617_), .B2(new_n604_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n618_), .B1(new_n617_), .B2(new_n604_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n614_), .A2(new_n619_), .ZN(new_n620_));
  NOR3_X1   g419(.A1(new_n543_), .A2(new_n602_), .A3(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n464_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n395_), .ZN(new_n623_));
  OR2_X1    g422(.A1(new_n623_), .A2(KEYINPUT99), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(KEYINPUT99), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NOR3_X1   g426(.A1(new_n622_), .A2(G1gat), .A3(new_n627_), .ZN(new_n628_));
  XOR2_X1   g427(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n629_));
  OR2_X1    g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n535_), .A2(new_n538_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n441_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n620_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n602_), .A2(new_n463_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n632_), .A2(new_n633_), .A3(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(G1gat), .B1(new_n635_), .B2(new_n395_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n628_), .A2(new_n629_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n630_), .A2(new_n636_), .A3(new_n637_), .ZN(G1324gat));
  NOR3_X1   g437(.A1(new_n622_), .A2(G8gat), .A3(new_n402_), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n639_), .B(KEYINPUT101), .Z(new_n640_));
  OAI21_X1  g439(.A(G8gat), .B1(new_n635_), .B2(new_n402_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT39), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n642_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g443(.A(G15gat), .B1(new_n635_), .B2(new_n429_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT41), .ZN(new_n646_));
  NOR3_X1   g445(.A1(new_n622_), .A2(G15gat), .A3(new_n429_), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n646_), .A2(new_n647_), .ZN(G1326gat));
  XNOR2_X1  g447(.A(new_n408_), .B(KEYINPUT102), .ZN(new_n649_));
  OAI21_X1  g448(.A(G22gat), .B1(new_n635_), .B2(new_n649_), .ZN(new_n650_));
  XOR2_X1   g449(.A(KEYINPUT103), .B(KEYINPUT42), .Z(new_n651_));
  XNOR2_X1  g450(.A(new_n650_), .B(new_n651_), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n649_), .A2(G22gat), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n652_), .B1(new_n622_), .B2(new_n653_), .ZN(G1327gat));
  NAND2_X1  g453(.A1(new_n631_), .A2(new_n620_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n602_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n464_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(G29gat), .B1(new_n658_), .B2(new_n623_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(KEYINPUT104), .A2(KEYINPUT43), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(KEYINPUT104), .A2(KEYINPUT43), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n664_), .B1(new_n441_), .B2(new_n542_), .ZN(new_n665_));
  AOI22_X1  g464(.A1(new_n393_), .A2(new_n357_), .B1(new_n409_), .B2(KEYINPUT97), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n428_), .B1(new_n666_), .B2(new_n412_), .ZN(new_n667_));
  AND4_X1   g466(.A1(new_n395_), .A2(new_n437_), .A3(new_n439_), .A4(new_n427_), .ZN(new_n668_));
  OAI211_X1 g467(.A(new_n543_), .B(new_n660_), .C1(new_n667_), .C2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n665_), .A2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n634_), .A2(new_n620_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n670_), .A2(KEYINPUT44), .A3(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT105), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n671_), .B1(new_n665_), .B2(new_n669_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n676_), .A2(KEYINPUT105), .A3(KEYINPUT44), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n413_), .A2(new_n429_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n440_), .A2(new_n395_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n663_), .B1(new_n681_), .B2(new_n543_), .ZN(new_n682_));
  AOI211_X1 g481(.A(new_n542_), .B(new_n661_), .C1(new_n679_), .C2(new_n680_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n672_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  AOI22_X1  g483(.A1(new_n675_), .A2(new_n677_), .B1(new_n678_), .B2(new_n684_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n626_), .A2(G29gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n659_), .B1(new_n685_), .B2(new_n686_), .ZN(G1328gat));
  NOR3_X1   g486(.A1(new_n657_), .A2(G36gat), .A3(new_n402_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n688_), .B(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n436_), .B1(new_n676_), .B2(KEYINPUT44), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n691_), .B1(new_n675_), .B2(new_n677_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT106), .ZN(new_n693_));
  INV_X1    g492(.A(G36gat), .ZN(new_n694_));
  NOR3_X1   g493(.A1(new_n692_), .A2(new_n693_), .A3(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n402_), .B1(new_n684_), .B2(new_n678_), .ZN(new_n696_));
  AND4_X1   g495(.A1(KEYINPUT105), .A2(new_n670_), .A3(KEYINPUT44), .A4(new_n672_), .ZN(new_n697_));
  AOI21_X1  g496(.A(KEYINPUT105), .B1(new_n676_), .B2(KEYINPUT44), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n696_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(KEYINPUT106), .B1(new_n699_), .B2(G36gat), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n690_), .B1(new_n695_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT46), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  OAI211_X1 g502(.A(KEYINPUT46), .B(new_n690_), .C1(new_n695_), .C2(new_n700_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(G1329gat));
  NAND3_X1  g504(.A1(new_n685_), .A2(G43gat), .A3(new_n427_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n415_), .B1(new_n657_), .B2(new_n429_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n708_), .B(new_n709_), .ZN(G1330gat));
  INV_X1    g509(.A(new_n649_), .ZN(new_n711_));
  AOI21_X1  g510(.A(G50gat), .B1(new_n658_), .B2(new_n711_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n408_), .A2(G50gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n685_), .B2(new_n713_), .ZN(G1331gat));
  NOR2_X1   g513(.A1(new_n441_), .A2(new_n462_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n543_), .A2(new_n620_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n715_), .A2(new_n602_), .A3(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(G57gat), .B1(new_n718_), .B2(new_n626_), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n632_), .A2(new_n463_), .A3(new_n602_), .A4(new_n633_), .ZN(new_n720_));
  XOR2_X1   g519(.A(KEYINPUT109), .B(G57gat), .Z(new_n721_));
  NOR3_X1   g520(.A1(new_n720_), .A2(new_n395_), .A3(new_n721_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n719_), .A2(new_n722_), .ZN(G1332gat));
  OAI21_X1  g522(.A(G64gat), .B1(new_n720_), .B2(new_n402_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT48), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n718_), .A2(new_n551_), .A3(new_n436_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1333gat));
  OAI21_X1  g526(.A(G71gat), .B1(new_n720_), .B2(new_n429_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT49), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n718_), .A2(new_n554_), .A3(new_n428_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1334gat));
  OAI21_X1  g530(.A(G78gat), .B1(new_n720_), .B2(new_n649_), .ZN(new_n732_));
  XOR2_X1   g531(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n733_));
  XNOR2_X1  g532(.A(new_n732_), .B(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n718_), .A2(new_n556_), .A3(new_n711_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(G1335gat));
  NOR3_X1   g535(.A1(new_n601_), .A2(new_n462_), .A3(new_n633_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n670_), .A2(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(G85gat), .B1(new_n738_), .B2(new_n395_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n601_), .A2(new_n655_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n715_), .A2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(G85gat), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n626_), .A2(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n739_), .B1(new_n741_), .B2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT111), .ZN(G1336gat));
  OAI21_X1  g544(.A(G92gat), .B1(new_n738_), .B2(new_n402_), .ZN(new_n746_));
  OR3_X1    g545(.A1(new_n741_), .A2(G92gat), .A3(new_n402_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(G1337gat));
  OAI21_X1  g547(.A(G99gat), .B1(new_n738_), .B2(new_n429_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n741_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n750_), .A2(new_n427_), .A3(new_n477_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n749_), .A2(new_n751_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(KEYINPUT112), .B(KEYINPUT51), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n752_), .B(new_n753_), .ZN(G1338gat));
  NAND3_X1  g553(.A1(new_n750_), .A2(new_n478_), .A3(new_n408_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n670_), .A2(new_n408_), .A3(new_n737_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n756_), .A2(G106gat), .A3(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n757_), .B1(new_n756_), .B2(G106gat), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n755_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g560(.A1(new_n626_), .A2(new_n440_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n461_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n452_), .B1(new_n456_), .B2(new_n450_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n455_), .A2(new_n764_), .ZN(new_n765_));
  AOI22_X1  g564(.A1(new_n458_), .A2(new_n461_), .B1(new_n763_), .B2(new_n765_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n766_), .B1(new_n593_), .B2(new_n595_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT116), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n462_), .A2(new_n592_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n594_), .ZN(new_n770_));
  AND4_X1   g569(.A1(new_n581_), .A2(new_n572_), .A3(new_n582_), .A4(new_n578_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n572_), .A2(new_n578_), .A3(new_n582_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(new_n580_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n771_), .B1(KEYINPUT55), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT55), .ZN(new_n775_));
  NOR3_X1   g574(.A1(new_n772_), .A2(new_n775_), .A3(new_n580_), .ZN(new_n776_));
  OAI211_X1 g575(.A(KEYINPUT56), .B(new_n770_), .C1(new_n774_), .C2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT115), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n769_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n770_), .B1(new_n774_), .B2(new_n776_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT56), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n783_), .A2(KEYINPUT115), .A3(new_n777_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n768_), .B1(new_n780_), .B2(new_n784_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n785_), .A2(new_n631_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n592_), .A2(new_n766_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n783_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n787_), .B1(new_n788_), .B2(new_n778_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT58), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n542_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  OAI211_X1 g590(.A(KEYINPUT58), .B(new_n787_), .C1(new_n788_), .C2(new_n778_), .ZN(new_n792_));
  AOI22_X1  g591(.A1(new_n786_), .A2(KEYINPUT57), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT118), .ZN(new_n794_));
  INV_X1    g593(.A(new_n768_), .ZN(new_n795_));
  AND3_X1   g594(.A1(new_n783_), .A2(KEYINPUT115), .A3(new_n777_), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n462_), .B(new_n592_), .C1(new_n777_), .C2(KEYINPUT115), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n795_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n631_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  XOR2_X1   g599(.A(KEYINPUT117), .B(KEYINPUT57), .Z(new_n801_));
  AOI21_X1  g600(.A(new_n794_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n794_), .B(new_n801_), .C1(new_n785_), .C2(new_n631_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n793_), .B1(new_n802_), .B2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT119), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT119), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n793_), .B(new_n807_), .C1(new_n802_), .C2(new_n804_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n806_), .A2(new_n620_), .A3(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT54), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n716_), .A2(new_n810_), .A3(new_n463_), .A4(new_n601_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(KEYINPUT114), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n621_), .A2(new_n463_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT54), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT114), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n621_), .A2(new_n815_), .A3(new_n810_), .A4(new_n463_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n812_), .A2(new_n814_), .A3(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n762_), .B1(new_n809_), .B2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n800_), .A2(new_n801_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n633_), .B1(new_n793_), .B2(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n817_), .B1(new_n821_), .B2(KEYINPUT120), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n821_), .A2(KEYINPUT120), .ZN(new_n823_));
  OR2_X1    g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n762_), .A2(KEYINPUT59), .ZN(new_n825_));
  AOI22_X1  g624(.A1(new_n819_), .A2(KEYINPUT59), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n462_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(G113gat), .ZN(new_n828_));
  OR2_X1    g627(.A1(new_n463_), .A2(G113gat), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n828_), .B1(new_n819_), .B2(new_n829_), .ZN(G1340gat));
  OAI21_X1  g629(.A(new_n825_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT59), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n602_), .B(new_n831_), .C1(new_n818_), .C2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(G120gat), .ZN(new_n834_));
  INV_X1    g633(.A(G120gat), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n835_), .B1(new_n601_), .B2(KEYINPUT60), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n818_), .B(new_n836_), .C1(KEYINPUT60), .C2(new_n835_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n834_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT121), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n834_), .A2(KEYINPUT121), .A3(new_n837_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(G1341gat));
  NAND2_X1  g641(.A1(new_n826_), .A2(new_n633_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(G127gat), .ZN(new_n844_));
  OR2_X1    g643(.A1(new_n620_), .A2(G127gat), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n844_), .B1(new_n819_), .B2(new_n845_), .ZN(G1342gat));
  NAND2_X1  g645(.A1(new_n826_), .A2(new_n543_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(G134gat), .ZN(new_n848_));
  OR2_X1    g647(.A1(new_n799_), .A2(G134gat), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n848_), .B1(new_n819_), .B2(new_n849_), .ZN(G1343gat));
  NAND2_X1  g649(.A1(new_n809_), .A2(new_n817_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT122), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n428_), .A2(new_n393_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n627_), .A2(new_n436_), .A3(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n851_), .A2(new_n852_), .A3(new_n855_), .ZN(new_n856_));
  AND3_X1   g655(.A1(new_n812_), .A2(new_n814_), .A3(new_n816_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n633_), .B1(new_n805_), .B2(KEYINPUT119), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n857_), .B1(new_n858_), .B2(new_n808_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n855_), .ZN(new_n860_));
  OAI21_X1  g659(.A(KEYINPUT122), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n856_), .A2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n462_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(KEYINPUT123), .B(G141gat), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n863_), .B(new_n864_), .ZN(G1344gat));
  NAND2_X1  g664(.A1(new_n862_), .A2(new_n602_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g666(.A1(new_n862_), .A2(new_n633_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(KEYINPUT61), .B(G155gat), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n868_), .B(new_n869_), .ZN(G1346gat));
  INV_X1    g669(.A(G162gat), .ZN(new_n871_));
  AOI211_X1 g670(.A(new_n871_), .B(new_n542_), .C1(new_n856_), .C2(new_n861_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n862_), .A2(new_n631_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT124), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n873_), .A2(new_n874_), .A3(new_n871_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n799_), .B1(new_n856_), .B2(new_n861_), .ZN(new_n876_));
  OAI21_X1  g675(.A(KEYINPUT124), .B1(new_n876_), .B2(G162gat), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n872_), .B1(new_n875_), .B2(new_n877_), .ZN(G1347gat));
  NOR3_X1   g677(.A1(new_n626_), .A2(new_n402_), .A3(new_n429_), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n824_), .A2(new_n462_), .A3(new_n649_), .A4(new_n879_), .ZN(new_n880_));
  OAI21_X1  g679(.A(KEYINPUT62), .B1(new_n880_), .B2(KEYINPUT22), .ZN(new_n881_));
  OAI21_X1  g680(.A(G169gat), .B1(new_n880_), .B2(KEYINPUT62), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n883_), .B1(new_n254_), .B2(new_n881_), .ZN(G1348gat));
  AND3_X1   g683(.A1(new_n824_), .A2(new_n649_), .A3(new_n879_), .ZN(new_n885_));
  AOI21_X1  g684(.A(G176gat), .B1(new_n885_), .B2(new_n602_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n859_), .A2(new_n408_), .ZN(new_n887_));
  AND3_X1   g686(.A1(new_n879_), .A2(G176gat), .A3(new_n602_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n886_), .B1(new_n887_), .B2(new_n888_), .ZN(G1349gat));
  AND2_X1   g688(.A1(new_n879_), .A2(new_n633_), .ZN(new_n890_));
  AND4_X1   g689(.A1(new_n262_), .A2(new_n824_), .A3(new_n649_), .A4(new_n890_), .ZN(new_n891_));
  AND2_X1   g690(.A1(new_n887_), .A2(new_n890_), .ZN(new_n892_));
  OR2_X1    g691(.A1(new_n892_), .A2(KEYINPUT125), .ZN(new_n893_));
  AOI21_X1  g692(.A(G183gat), .B1(new_n892_), .B2(KEYINPUT125), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n891_), .B1(new_n893_), .B2(new_n894_), .ZN(G1350gat));
  NAND2_X1  g694(.A1(new_n885_), .A2(new_n543_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(G190gat), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n799_), .A2(new_n263_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(KEYINPUT126), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n885_), .A2(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n897_), .A2(new_n900_), .ZN(G1351gat));
  NOR4_X1   g700(.A1(new_n859_), .A2(new_n623_), .A3(new_n402_), .A4(new_n854_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(new_n462_), .ZN(new_n903_));
  XOR2_X1   g702(.A(KEYINPUT127), .B(G197gat), .Z(new_n904_));
  XNOR2_X1  g703(.A(new_n903_), .B(new_n904_), .ZN(G1352gat));
  NAND2_X1  g704(.A1(new_n902_), .A2(new_n602_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g706(.A1(new_n902_), .A2(new_n633_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(KEYINPUT63), .B(G211gat), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n910_), .B1(new_n908_), .B2(new_n911_), .ZN(G1354gat));
  INV_X1    g711(.A(G218gat), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n902_), .A2(new_n913_), .A3(new_n631_), .ZN(new_n914_));
  AND2_X1   g713(.A1(new_n902_), .A2(new_n543_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n914_), .B1(new_n915_), .B2(new_n913_), .ZN(G1355gat));
endmodule


