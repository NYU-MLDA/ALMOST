//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 1 1 1 1 1 0 1 1 0 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 0 1 0 0 1 1 0 0 1 0 1 1 1 0 0 0 0 0 1 0 1 0 1 0 1 0 1 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n599_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n853_, new_n854_, new_n855_, new_n856_, new_n858_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n896_, new_n897_, new_n898_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_;
  XNOR2_X1  g000(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G71gat), .B(G99gat), .ZN(new_n204_));
  INV_X1    g003(.A(G43gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT30), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G227gat), .A2(G233gat), .ZN(new_n208_));
  INV_X1    g007(.A(G15gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n207_), .B(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT23), .ZN(new_n213_));
  OR3_X1    g012(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n214_));
  AND2_X1   g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT25), .B(G183gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT26), .B(G190gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT76), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n215_), .A2(new_n218_), .A3(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT79), .B(G176gat), .ZN(new_n225_));
  INV_X1    g024(.A(G169gat), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n225_), .B1(KEYINPUT22), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT22), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n226_), .A2(KEYINPUT77), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT77), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(G169gat), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n228_), .B1(new_n229_), .B2(new_n231_), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n232_), .A2(KEYINPUT78), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(KEYINPUT78), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n227_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n213_), .B1(G183gat), .B2(G190gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(new_n220_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n224_), .B1(new_n235_), .B2(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(KEYINPUT82), .B1(new_n211_), .B2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n210_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n207_), .B(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n238_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  OAI21_X1  g042(.A(KEYINPUT83), .B1(new_n239_), .B2(new_n243_), .ZN(new_n244_));
  XOR2_X1   g043(.A(G127gat), .B(G134gat), .Z(new_n245_));
  XOR2_X1   g044(.A(G113gat), .B(G120gat), .Z(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT80), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n245_), .A2(new_n246_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n211_), .A2(new_n238_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n241_), .A2(new_n242_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT83), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n253_), .A2(new_n254_), .A3(KEYINPUT82), .A4(new_n255_), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n244_), .A2(new_n252_), .A3(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n252_), .B1(new_n244_), .B2(new_n256_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n203_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n244_), .A2(new_n256_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(new_n251_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n244_), .A2(new_n252_), .A3(new_n256_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n261_), .A2(new_n202_), .A3(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n259_), .A2(new_n263_), .ZN(new_n264_));
  XOR2_X1   g063(.A(G197gat), .B(G204gat), .Z(new_n265_));
  OR2_X1    g064(.A1(new_n265_), .A2(KEYINPUT21), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(KEYINPUT21), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G211gat), .B(G218gat), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n266_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n269_));
  OR2_X1    g068(.A1(new_n267_), .A2(new_n268_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G155gat), .A2(G162gat), .ZN(new_n272_));
  NOR2_X1   g071(.A1(G155gat), .A2(G162gat), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  OR3_X1    g073(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n275_));
  OAI21_X1  g074(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT85), .ZN(new_n277_));
  AOI22_X1  g076(.A1(new_n277_), .A2(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n277_), .A2(KEYINPUT2), .ZN(new_n279_));
  OAI211_X1 g078(.A(new_n275_), .B(new_n276_), .C1(new_n278_), .C2(new_n279_), .ZN(new_n280_));
  AND2_X1   g079(.A1(new_n278_), .A2(new_n279_), .ZN(new_n281_));
  OAI211_X1 g080(.A(new_n272_), .B(new_n274_), .C1(new_n280_), .C2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n272_), .A2(KEYINPUT1), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT84), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n272_), .A2(KEYINPUT1), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n272_), .A2(KEYINPUT84), .A3(KEYINPUT1), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n285_), .A2(new_n286_), .A3(new_n287_), .A4(new_n274_), .ZN(new_n288_));
  OR2_X1    g087(.A1(G141gat), .A2(G148gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G141gat), .A2(G148gat), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n288_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  AND2_X1   g090(.A1(new_n282_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT29), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n271_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G228gat), .A2(G233gat), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n294_), .B(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G78gat), .B(G106gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n294_), .B(new_n295_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n298_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n299_), .A2(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(KEYINPUT87), .B1(new_n297_), .B2(new_n298_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n282_), .A2(new_n291_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n306_));
  OR3_X1    g105(.A1(new_n305_), .A2(KEYINPUT29), .A3(new_n306_), .ZN(new_n307_));
  XOR2_X1   g106(.A(G22gat), .B(G50gat), .Z(new_n308_));
  OAI21_X1  g107(.A(new_n306_), .B1(new_n305_), .B2(KEYINPUT29), .ZN(new_n309_));
  AND3_X1   g108(.A1(new_n307_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n308_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n303_), .B1(new_n304_), .B2(new_n313_), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n299_), .A2(new_n302_), .A3(new_n312_), .A4(KEYINPUT87), .ZN(new_n315_));
  AND2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT22), .B(G169gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n225_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(new_n220_), .ZN(new_n319_));
  OR2_X1    g118(.A1(new_n319_), .A2(KEYINPUT90), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(KEYINPUT90), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n320_), .A2(new_n236_), .A3(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT89), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n217_), .B(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(new_n216_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n222_), .A2(new_n219_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n325_), .A2(new_n215_), .A3(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n322_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(new_n271_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n271_), .ZN(new_n330_));
  OAI211_X1 g129(.A(new_n330_), .B(new_n224_), .C1(new_n235_), .C2(new_n237_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n329_), .A2(new_n331_), .A3(KEYINPUT20), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G226gat), .A2(G233gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n332_), .A2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G8gat), .B(G36gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT18), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G64gat), .B(G92gat), .ZN(new_n340_));
  XOR2_X1   g139(.A(new_n339_), .B(new_n340_), .Z(new_n341_));
  NAND3_X1  g140(.A1(new_n330_), .A2(new_n322_), .A3(new_n327_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n238_), .A2(new_n271_), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n342_), .A2(new_n343_), .A3(KEYINPUT20), .A4(new_n335_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n337_), .A2(new_n341_), .A3(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n341_), .B1(new_n337_), .B2(new_n344_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G225gat), .A2(G233gat), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT4), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n252_), .A2(new_n305_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n305_), .B1(new_n250_), .B2(new_n247_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n351_), .B1(new_n352_), .B2(new_n354_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n251_), .A2(new_n292_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n356_), .A2(KEYINPUT4), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n350_), .B1(new_n355_), .B2(new_n357_), .ZN(new_n358_));
  XOR2_X1   g157(.A(G1gat), .B(G29gat), .Z(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT91), .B(G85gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT0), .B(G57gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n352_), .A2(new_n354_), .A3(KEYINPUT92), .A4(new_n349_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n352_), .A2(new_n354_), .A3(new_n349_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT92), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n358_), .A2(new_n363_), .A3(new_n364_), .A4(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT33), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  AND2_X1   g169(.A1(new_n367_), .A2(new_n364_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n371_), .A2(KEYINPUT33), .A3(new_n363_), .A4(new_n358_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n349_), .B1(new_n355_), .B2(new_n357_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n363_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n352_), .A2(new_n350_), .A3(new_n354_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n373_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n348_), .A2(new_n370_), .A3(new_n372_), .A4(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n367_), .A2(new_n364_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n352_), .A2(new_n351_), .ZN(new_n379_));
  OAI21_X1  g178(.A(KEYINPUT4), .B1(new_n356_), .B2(new_n353_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n349_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n374_), .B1(new_n378_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(new_n368_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n342_), .A2(new_n343_), .A3(KEYINPUT20), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(new_n336_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n385_), .B1(new_n332_), .B2(new_n336_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n386_), .A2(KEYINPUT32), .A3(new_n341_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n341_), .A2(KEYINPUT32), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n337_), .A2(new_n344_), .A3(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n383_), .A2(new_n387_), .A3(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n316_), .B1(new_n377_), .B2(new_n390_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n314_), .A2(new_n368_), .A3(new_n382_), .A4(new_n315_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n345_), .A2(KEYINPUT93), .ZN(new_n393_));
  INV_X1    g192(.A(new_n341_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n386_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT93), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n337_), .A2(new_n396_), .A3(new_n341_), .A4(new_n344_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n393_), .A2(new_n395_), .A3(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT27), .ZN(new_n399_));
  OR3_X1    g198(.A1(new_n346_), .A2(new_n347_), .A3(KEYINPUT27), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n392_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n264_), .B1(new_n391_), .B2(new_n401_), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n259_), .A2(new_n263_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n383_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n314_), .A2(new_n315_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n399_), .A2(new_n400_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n403_), .A2(new_n404_), .A3(new_n405_), .A4(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n402_), .A2(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G29gat), .B(G36gat), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  XOR2_X1   g209(.A(G43gat), .B(G50gat), .Z(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G43gat), .B(G50gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n409_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(KEYINPUT68), .B(KEYINPUT15), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n415_), .B(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G15gat), .B(G22gat), .ZN(new_n418_));
  INV_X1    g217(.A(G1gat), .ZN(new_n419_));
  INV_X1    g218(.A(G8gat), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT14), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n418_), .A2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G1gat), .B(G8gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n417_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n424_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(new_n415_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G229gat), .A2(G233gat), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n425_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n424_), .B(new_n415_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT75), .ZN(new_n431_));
  NOR3_X1   g230(.A1(new_n430_), .A2(new_n431_), .A3(new_n428_), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n412_), .A2(new_n414_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n424_), .B(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n428_), .ZN(new_n435_));
  AOI21_X1  g234(.A(KEYINPUT75), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n429_), .B1(new_n432_), .B2(new_n436_), .ZN(new_n437_));
  XOR2_X1   g236(.A(G169gat), .B(G197gat), .Z(new_n438_));
  XNOR2_X1  g237(.A(G113gat), .B(G141gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n438_), .B(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n437_), .A2(new_n441_), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n429_), .B(new_n440_), .C1(new_n432_), .C2(new_n436_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT74), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G57gat), .B(G64gat), .ZN(new_n446_));
  OR2_X1    g245(.A1(new_n446_), .A2(KEYINPUT11), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(KEYINPUT11), .ZN(new_n448_));
  XOR2_X1   g247(.A(G71gat), .B(G78gat), .Z(new_n449_));
  NAND3_X1  g248(.A1(new_n447_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  OR2_X1    g249(.A1(new_n448_), .A2(new_n449_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G231gat), .A2(G233gat), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n424_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n424_), .A2(new_n454_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n452_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n457_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n452_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n459_), .A2(new_n460_), .A3(new_n455_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n458_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT70), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G127gat), .B(G155gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(KEYINPUT16), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G183gat), .B(G211gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n466_), .B(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(KEYINPUT71), .B(KEYINPUT17), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT72), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n470_), .B(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n458_), .A2(new_n461_), .A3(KEYINPUT70), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n464_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n474_));
  XOR2_X1   g273(.A(new_n468_), .B(KEYINPUT17), .Z(new_n475_));
  NAND3_X1  g274(.A1(new_n475_), .A2(new_n461_), .A3(new_n458_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT73), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n474_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n477_), .B1(new_n474_), .B2(new_n476_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n445_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n480_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n482_), .A2(KEYINPUT74), .A3(new_n478_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n481_), .A2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT67), .B(KEYINPUT34), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G232gat), .A2(G233gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n485_), .B(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT35), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT7), .ZN(new_n489_));
  INV_X1    g288(.A(G99gat), .ZN(new_n490_));
  INV_X1    g289(.A(G106gat), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n489_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT64), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G99gat), .A2(G106gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(KEYINPUT6), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT6), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n497_), .A2(G99gat), .A3(G106gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  OAI21_X1  g298(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n489_), .A2(new_n490_), .A3(new_n491_), .A4(KEYINPUT64), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n494_), .A2(new_n499_), .A3(new_n500_), .A4(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(G85gat), .ZN(new_n503_));
  INV_X1    g302(.A(G92gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G85gat), .A2(G92gat), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n502_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT8), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n502_), .A2(KEYINPUT8), .A3(new_n507_), .ZN(new_n511_));
  OR2_X1    g310(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n512_), .A2(new_n491_), .A3(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n505_), .A2(KEYINPUT9), .A3(new_n506_), .ZN(new_n515_));
  OR2_X1    g314(.A1(new_n506_), .A2(KEYINPUT9), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n499_), .A2(new_n514_), .A3(new_n515_), .A4(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n510_), .A2(new_n511_), .A3(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n417_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT69), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n488_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n519_), .B1(new_n433_), .B2(new_n518_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G190gat), .B(G218gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G134gat), .B(G162gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  AOI22_X1  g325(.A1(new_n522_), .A2(new_n523_), .B1(KEYINPUT36), .B2(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n487_), .A2(KEYINPUT35), .ZN(new_n528_));
  OAI221_X1 g327(.A(new_n519_), .B1(new_n433_), .B2(new_n518_), .C1(new_n521_), .C2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(new_n529_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n526_), .A2(KEYINPUT36), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n527_), .B(new_n529_), .C1(KEYINPUT36), .C2(new_n526_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n532_), .A2(KEYINPUT37), .A3(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n532_), .A2(new_n533_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT37), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n484_), .A2(new_n534_), .A3(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G230gat), .A2(G233gat), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n502_), .A2(KEYINPUT8), .A3(new_n507_), .ZN(new_n541_));
  AOI21_X1  g340(.A(KEYINPUT8), .B1(new_n502_), .B2(new_n507_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n517_), .ZN(new_n543_));
  NOR3_X1   g342(.A1(new_n541_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n540_), .B1(new_n544_), .B2(new_n452_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n543_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n546_));
  AOI211_X1 g345(.A(KEYINPUT12), .B(new_n452_), .C1(new_n546_), .C2(new_n511_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT12), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n548_), .B1(new_n518_), .B2(new_n460_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n545_), .B1(new_n547_), .B2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(KEYINPUT65), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n518_), .A2(new_n460_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n546_), .A2(new_n452_), .A3(new_n511_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(new_n540_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT65), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n556_), .B(new_n545_), .C1(new_n547_), .C2(new_n549_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n551_), .A2(new_n555_), .A3(new_n557_), .ZN(new_n558_));
  XOR2_X1   g357(.A(G120gat), .B(G148gat), .Z(new_n559_));
  XNOR2_X1  g358(.A(KEYINPUT66), .B(KEYINPUT5), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G176gat), .B(G204gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n558_), .A2(new_n564_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n551_), .A2(new_n555_), .A3(new_n557_), .A4(new_n563_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  OR2_X1    g366(.A1(new_n567_), .A2(KEYINPUT13), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(KEYINPUT13), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n538_), .A2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n408_), .A2(new_n444_), .A3(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT94), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n383_), .B(KEYINPUT95), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n575_), .A2(G1gat), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n573_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT38), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n573_), .A2(KEYINPUT38), .A3(new_n576_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n479_), .A2(new_n480_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n444_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n570_), .A2(new_n582_), .ZN(new_n583_));
  AND4_X1   g382(.A1(new_n408_), .A2(new_n581_), .A3(new_n535_), .A4(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(new_n383_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(G1gat), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n579_), .A2(new_n580_), .A3(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT96), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(G1324gat));
  INV_X1    g388(.A(new_n406_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n573_), .A2(new_n420_), .A3(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n584_), .A2(new_n590_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(KEYINPUT97), .A2(KEYINPUT39), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n420_), .B1(KEYINPUT97), .B2(KEYINPUT39), .ZN(new_n594_));
  AND3_X1   g393(.A1(new_n592_), .A2(new_n593_), .A3(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n593_), .B1(new_n592_), .B2(new_n594_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n591_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  XOR2_X1   g396(.A(new_n597_), .B(KEYINPUT40), .Z(G1325gat));
  NAND2_X1  g397(.A1(new_n584_), .A2(new_n403_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(G15gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(KEYINPUT98), .B(KEYINPUT41), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n601_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n573_), .A2(new_n209_), .A3(new_n403_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n602_), .A2(new_n603_), .A3(new_n604_), .ZN(G1326gat));
  INV_X1    g404(.A(G22gat), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n606_), .B1(new_n584_), .B2(new_n316_), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n607_), .B(KEYINPUT42), .Z(new_n608_));
  NOR2_X1   g407(.A1(new_n405_), .A2(G22gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT99), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n573_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n608_), .A2(new_n611_), .ZN(G1327gat));
  INV_X1    g411(.A(new_n484_), .ZN(new_n613_));
  OAI211_X1 g412(.A(new_n583_), .B(new_n613_), .C1(KEYINPUT102), .C2(KEYINPUT44), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n537_), .A2(new_n534_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n377_), .A2(new_n390_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(new_n405_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n392_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n406_), .A2(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n403_), .B1(new_n618_), .B2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n406_), .A2(new_n405_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n259_), .A2(new_n263_), .A3(new_n404_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n616_), .B1(new_n621_), .B2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT100), .ZN(new_n626_));
  AOI21_X1  g425(.A(KEYINPUT43), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n616_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n628_), .B1(new_n402_), .B2(new_n407_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT43), .ZN(new_n630_));
  NOR3_X1   g429(.A1(new_n629_), .A2(KEYINPUT100), .A3(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n615_), .B1(new_n627_), .B2(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(KEYINPUT102), .B1(KEYINPUT101), .B2(KEYINPUT44), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n625_), .A2(new_n626_), .A3(KEYINPUT43), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n630_), .B1(new_n629_), .B2(KEYINPUT100), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n638_), .A2(new_n615_), .A3(new_n633_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n575_), .B1(new_n635_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(G29gat), .ZN(new_n641_));
  INV_X1    g440(.A(new_n535_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n613_), .A2(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n643_), .A2(new_n570_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n408_), .A2(new_n444_), .A3(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT103), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n408_), .A2(KEYINPUT103), .A3(new_n444_), .A4(new_n644_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n383_), .A2(new_n641_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT104), .ZN(new_n651_));
  OAI22_X1  g450(.A1(new_n640_), .A2(new_n641_), .B1(new_n649_), .B2(new_n651_), .ZN(G1328gat));
  NOR2_X1   g451(.A1(new_n406_), .A2(G36gat), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  OR3_X1    g453(.A1(new_n649_), .A2(KEYINPUT45), .A3(new_n654_), .ZN(new_n655_));
  OAI21_X1  g454(.A(KEYINPUT45), .B1(new_n649_), .B2(new_n654_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n406_), .B1(new_n635_), .B2(new_n639_), .ZN(new_n658_));
  INV_X1    g457(.A(G36gat), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n657_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT46), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  OAI211_X1 g461(.A(new_n657_), .B(KEYINPUT46), .C1(new_n658_), .C2(new_n659_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1329gat));
  INV_X1    g463(.A(new_n649_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n665_), .A2(new_n205_), .A3(new_n403_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n264_), .B1(new_n635_), .B2(new_n639_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n666_), .B1(new_n667_), .B2(new_n205_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT47), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  OAI211_X1 g469(.A(KEYINPUT47), .B(new_n666_), .C1(new_n667_), .C2(new_n205_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(G1330gat));
  INV_X1    g471(.A(KEYINPUT105), .ZN(new_n673_));
  INV_X1    g472(.A(G50gat), .ZN(new_n674_));
  AOI211_X1 g473(.A(new_n674_), .B(new_n405_), .C1(new_n635_), .C2(new_n639_), .ZN(new_n675_));
  AOI21_X1  g474(.A(G50gat), .B1(new_n665_), .B2(new_n316_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n673_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n635_), .A2(new_n639_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n405_), .A2(new_n674_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n676_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(KEYINPUT105), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n677_), .A2(new_n681_), .ZN(G1331gat));
  NAND2_X1  g481(.A1(new_n408_), .A2(new_n535_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n570_), .ZN(new_n685_));
  NOR3_X1   g484(.A1(new_n685_), .A2(new_n444_), .A3(new_n613_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(new_n687_));
  OAI21_X1  g486(.A(G57gat), .B1(new_n687_), .B2(new_n404_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n685_), .A2(new_n444_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n408_), .A2(new_n689_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n690_), .A2(new_n538_), .ZN(new_n691_));
  INV_X1    g490(.A(G57gat), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n691_), .A2(new_n692_), .A3(new_n574_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n688_), .A2(new_n693_), .ZN(G1332gat));
  INV_X1    g493(.A(G64gat), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n691_), .A2(new_n695_), .A3(new_n590_), .ZN(new_n696_));
  OAI21_X1  g495(.A(G64gat), .B1(new_n687_), .B2(new_n406_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n697_), .A2(KEYINPUT48), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n697_), .A2(KEYINPUT48), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n696_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT106), .ZN(G1333gat));
  OAI21_X1  g500(.A(G71gat), .B1(new_n687_), .B2(new_n264_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT49), .ZN(new_n703_));
  INV_X1    g502(.A(G71gat), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n691_), .A2(new_n704_), .A3(new_n403_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(G1334gat));
  INV_X1    g505(.A(G78gat), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n691_), .A2(new_n707_), .A3(new_n316_), .ZN(new_n708_));
  OAI21_X1  g507(.A(G78gat), .B1(new_n687_), .B2(new_n405_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n709_), .A2(KEYINPUT50), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(KEYINPUT50), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n708_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT107), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n712_), .B(new_n713_), .ZN(G1335gat));
  NOR2_X1   g513(.A1(new_n690_), .A2(new_n643_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n715_), .A2(new_n503_), .A3(new_n574_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n638_), .A2(KEYINPUT108), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n689_), .A2(new_n613_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT108), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n636_), .A2(new_n637_), .A3(new_n720_), .ZN(new_n721_));
  AND4_X1   g520(.A1(new_n383_), .A2(new_n717_), .A3(new_n719_), .A4(new_n721_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n716_), .B1(new_n722_), .B2(new_n503_), .ZN(G1336gat));
  NAND2_X1  g522(.A1(new_n590_), .A2(G92gat), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT109), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n717_), .A2(new_n719_), .A3(new_n721_), .A4(new_n725_), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n690_), .A2(new_n406_), .A3(new_n643_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n726_), .B1(G92gat), .B2(new_n727_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT110), .ZN(G1337gat));
  NAND3_X1  g528(.A1(new_n717_), .A2(new_n719_), .A3(new_n721_), .ZN(new_n730_));
  OAI21_X1  g529(.A(G99gat), .B1(new_n730_), .B2(new_n264_), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n715_), .A2(new_n403_), .A3(new_n512_), .A4(new_n513_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(KEYINPUT51), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT51), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n731_), .A2(new_n735_), .A3(new_n732_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(G1338gat));
  NAND3_X1  g536(.A1(new_n715_), .A2(new_n491_), .A3(new_n316_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT52), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n718_), .A2(new_n405_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n638_), .A2(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n739_), .B1(new_n741_), .B2(G106gat), .ZN(new_n742_));
  AOI211_X1 g541(.A(KEYINPUT52), .B(new_n491_), .C1(new_n638_), .C2(new_n740_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n738_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g544(.A1(new_n403_), .A2(new_n574_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n746_), .A2(new_n622_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n748_), .A2(KEYINPUT59), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n444_), .A2(new_n566_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT111), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT55), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n551_), .A2(new_n752_), .A3(new_n557_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n553_), .A2(new_n539_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n552_), .A2(KEYINPUT12), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n518_), .A2(new_n548_), .A3(new_n460_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n754_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n553_), .B1(new_n547_), .B2(new_n549_), .ZN(new_n758_));
  AOI22_X1  g557(.A1(new_n757_), .A2(KEYINPUT55), .B1(new_n758_), .B2(new_n540_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n753_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT113), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT56), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(KEYINPUT112), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n760_), .A2(new_n761_), .A3(new_n564_), .A4(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n563_), .B1(new_n753_), .B2(new_n759_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n764_), .B1(new_n765_), .B2(new_n763_), .ZN(new_n766_));
  AOI211_X1 g565(.A(new_n762_), .B(new_n563_), .C1(new_n753_), .C2(new_n759_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n767_), .A2(new_n761_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n751_), .B1(new_n766_), .B2(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n441_), .B1(new_n430_), .B2(new_n435_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT114), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT114), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n772_), .B(new_n441_), .C1(new_n430_), .C2(new_n435_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n425_), .A2(new_n427_), .A3(new_n435_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n771_), .A2(new_n773_), .A3(new_n774_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n775_), .A2(new_n443_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n567_), .A2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n769_), .A2(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(KEYINPUT57), .B1(new_n778_), .B2(new_n535_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT57), .ZN(new_n780_));
  AOI211_X1 g579(.A(new_n780_), .B(new_n642_), .C1(new_n769_), .C2(new_n777_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n779_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT58), .ZN(new_n783_));
  AOI21_X1  g582(.A(KEYINPUT56), .B1(new_n760_), .B2(new_n564_), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n784_), .A2(new_n767_), .A3(KEYINPUT115), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n760_), .A2(new_n564_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n786_), .A2(KEYINPUT115), .A3(new_n762_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n776_), .A2(new_n566_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n783_), .B1(new_n785_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT116), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(new_n792_), .A3(new_n616_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n786_), .A2(new_n762_), .ZN(new_n794_));
  AOI21_X1  g593(.A(KEYINPUT115), .B1(new_n765_), .B2(KEYINPUT56), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n788_), .B1(new_n784_), .B2(KEYINPUT115), .ZN(new_n797_));
  AOI21_X1  g596(.A(KEYINPUT58), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(KEYINPUT116), .B1(new_n798_), .B2(new_n628_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n796_), .A2(new_n797_), .A3(KEYINPUT58), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n793_), .A2(new_n799_), .A3(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n484_), .B1(new_n782_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT119), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT54), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(new_n571_), .B2(new_n582_), .ZN(new_n805_));
  NOR4_X1   g604(.A1(new_n538_), .A2(new_n570_), .A3(KEYINPUT54), .A4(new_n444_), .ZN(new_n806_));
  OAI22_X1  g605(.A1(new_n802_), .A2(new_n803_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  OR2_X1    g606(.A1(new_n765_), .A2(new_n763_), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n808_), .B(new_n764_), .C1(new_n761_), .C2(new_n767_), .ZN(new_n809_));
  AOI22_X1  g608(.A1(new_n809_), .A2(new_n751_), .B1(new_n567_), .B2(new_n776_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n780_), .B1(new_n810_), .B2(new_n642_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n778_), .A2(KEYINPUT57), .A3(new_n535_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n801_), .A2(new_n811_), .A3(new_n812_), .ZN(new_n813_));
  AND3_X1   g612(.A1(new_n813_), .A2(new_n803_), .A3(new_n613_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n749_), .B1(new_n807_), .B2(new_n814_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n805_), .A2(new_n806_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n581_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n816_), .B1(new_n813_), .B2(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(KEYINPUT59), .B1(new_n818_), .B2(new_n748_), .ZN(new_n819_));
  INV_X1    g618(.A(G113gat), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n582_), .A2(new_n820_), .ZN(new_n821_));
  AND3_X1   g620(.A1(new_n815_), .A2(new_n819_), .A3(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT117), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(new_n818_), .B2(new_n748_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n581_), .B1(new_n782_), .B2(new_n801_), .ZN(new_n825_));
  OAI211_X1 g624(.A(KEYINPUT117), .B(new_n747_), .C1(new_n825_), .C2(new_n816_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n824_), .A2(new_n444_), .A3(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n820_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT118), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT118), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n827_), .A2(new_n830_), .A3(new_n820_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n822_), .B1(new_n829_), .B2(new_n831_), .ZN(G1340gat));
  NAND3_X1  g631(.A1(new_n815_), .A2(new_n570_), .A3(new_n819_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(G120gat), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT60), .ZN(new_n835_));
  AOI21_X1  g634(.A(G120gat), .B1(new_n570_), .B2(new_n835_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n836_), .B(KEYINPUT120), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n837_), .B1(new_n835_), .B2(G120gat), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n824_), .A2(new_n826_), .A3(new_n838_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n839_), .A2(KEYINPUT121), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n839_), .A2(KEYINPUT121), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n834_), .B1(new_n840_), .B2(new_n841_), .ZN(G1341gat));
  NAND3_X1  g641(.A1(new_n815_), .A2(new_n581_), .A3(new_n819_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(G127gat), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n613_), .A2(G127gat), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n824_), .A2(new_n826_), .A3(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n846_), .ZN(G1342gat));
  NAND3_X1  g646(.A1(new_n815_), .A2(new_n616_), .A3(new_n819_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(G134gat), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n535_), .A2(G134gat), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n824_), .A2(new_n826_), .A3(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n851_), .ZN(G1343gat));
  NAND4_X1  g651(.A1(new_n574_), .A2(new_n264_), .A3(new_n406_), .A4(new_n316_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(KEYINPUT122), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n818_), .A2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n444_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n570_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g658(.A(KEYINPUT61), .B(G155gat), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT123), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n855_), .A2(new_n862_), .A3(new_n484_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n862_), .B1(new_n855_), .B2(new_n484_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n861_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n865_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n867_), .A2(new_n863_), .A3(new_n860_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n868_), .ZN(G1346gat));
  INV_X1    g668(.A(G162gat), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n855_), .A2(new_n870_), .A3(new_n642_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n855_), .A2(new_n616_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n871_), .B1(new_n873_), .B2(new_n870_), .ZN(G1347gat));
  NOR4_X1   g673(.A1(new_n574_), .A2(new_n264_), .A3(new_n406_), .A4(new_n316_), .ZN(new_n875_));
  OAI211_X1 g674(.A(new_n444_), .B(new_n875_), .C1(new_n807_), .C2(new_n814_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(G169gat), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT62), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  OR2_X1    g678(.A1(new_n807_), .A2(new_n814_), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n880_), .A2(new_n317_), .A3(new_n444_), .A4(new_n875_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n876_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n879_), .A2(new_n881_), .A3(new_n882_), .ZN(G1348gat));
  NAND2_X1  g682(.A1(new_n570_), .A2(G176gat), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n875_), .B(new_n885_), .C1(new_n825_), .C2(new_n816_), .ZN(new_n886_));
  XOR2_X1   g685(.A(new_n886_), .B(KEYINPUT124), .Z(new_n887_));
  NAND3_X1  g686(.A1(new_n880_), .A2(new_n570_), .A3(new_n875_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n887_), .B1(new_n225_), .B2(new_n888_), .ZN(G1349gat));
  AND2_X1   g688(.A1(new_n880_), .A2(new_n875_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n817_), .A2(new_n216_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n818_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n892_), .A2(new_n484_), .A3(new_n875_), .ZN(new_n893_));
  INV_X1    g692(.A(G183gat), .ZN(new_n894_));
  AOI22_X1  g693(.A1(new_n890_), .A2(new_n891_), .B1(new_n893_), .B2(new_n894_), .ZN(G1350gat));
  NAND3_X1  g694(.A1(new_n880_), .A2(new_n616_), .A3(new_n875_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(G190gat), .ZN(new_n897_));
  NAND4_X1  g696(.A1(new_n880_), .A2(new_n324_), .A3(new_n642_), .A4(new_n875_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(G1351gat));
  NOR3_X1   g698(.A1(new_n403_), .A2(new_n392_), .A3(new_n406_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n818_), .A2(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(new_n444_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n903_), .ZN(new_n904_));
  AOI21_X1  g703(.A(KEYINPUT125), .B1(new_n904_), .B2(G197gat), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n904_), .A2(G197gat), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT125), .ZN(new_n907_));
  INV_X1    g706(.A(G197gat), .ZN(new_n908_));
  NOR3_X1   g707(.A1(new_n903_), .A2(new_n907_), .A3(new_n908_), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n905_), .A2(new_n906_), .A3(new_n909_), .ZN(G1352gat));
  NAND2_X1  g709(.A1(new_n902_), .A2(new_n570_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g711(.A(new_n817_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n902_), .A2(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT127), .ZN(new_n915_));
  NOR2_X1   g714(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(KEYINPUT126), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n914_), .B1(new_n915_), .B2(new_n917_), .ZN(new_n918_));
  XOR2_X1   g717(.A(new_n917_), .B(KEYINPUT127), .Z(new_n919_));
  AOI21_X1  g718(.A(new_n918_), .B1(new_n914_), .B2(new_n919_), .ZN(G1354gat));
  INV_X1    g719(.A(new_n902_), .ZN(new_n921_));
  OAI21_X1  g720(.A(G218gat), .B1(new_n921_), .B2(new_n628_), .ZN(new_n922_));
  OR2_X1    g721(.A1(new_n535_), .A2(G218gat), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n922_), .B1(new_n921_), .B2(new_n923_), .ZN(G1355gat));
endmodule


