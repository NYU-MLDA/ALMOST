//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 1 0 0 1 1 1 0 0 1 0 1 0 0 0 0 1 0 1 0 1 1 1 0 1 0 1 0 0 0 1 1 0 0 0 1 0 1 0 0 1 0 0 0 1 0 0 0 0 1 1 1 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n715_, new_n716_,
    new_n717_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n726_, new_n727_, new_n728_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n835_, new_n836_, new_n838_,
    new_n839_, new_n841_, new_n842_, new_n843_, new_n844_, new_n846_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n857_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n892_, new_n893_, new_n894_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_;
  XOR2_X1   g000(.A(G71gat), .B(G99gat), .Z(new_n202_));
  NAND2_X1  g001(.A1(G227gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(G15gat), .B(G43gat), .Z(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT23), .ZN(new_n208_));
  INV_X1    g007(.A(G169gat), .ZN(new_n209_));
  INV_X1    g008(.A(G176gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT82), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT82), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n216_), .A2(KEYINPUT24), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT25), .B(G183gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT26), .B(G190gat), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n217_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT24), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n222_), .B1(new_n213_), .B2(new_n215_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n223_), .A2(KEYINPUT83), .A3(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(KEYINPUT83), .B1(new_n223_), .B2(new_n224_), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n208_), .B(new_n221_), .C1(new_n226_), .C2(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n208_), .B1(G183gat), .B2(G190gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT22), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n210_), .B1(new_n230_), .B2(KEYINPUT84), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(G169gat), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n214_), .B1(KEYINPUT84), .B2(new_n230_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n229_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n228_), .A2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT30), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n206_), .B1(new_n237_), .B2(KEYINPUT85), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT31), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G127gat), .B(G134gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G113gat), .B(G120gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n239_), .A2(new_n242_), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n238_), .A2(KEYINPUT31), .ZN(new_n244_));
  INV_X1    g043(.A(new_n242_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n238_), .A2(KEYINPUT31), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n244_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n243_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT85), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n236_), .A2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n248_), .B(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G155gat), .A2(G162gat), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT86), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(KEYINPUT86), .B1(G155gat), .B2(G162gat), .ZN(new_n255_));
  OR2_X1    g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(KEYINPUT88), .B1(new_n256_), .B2(KEYINPUT1), .ZN(new_n257_));
  OR4_X1    g056(.A1(KEYINPUT88), .A2(new_n254_), .A3(KEYINPUT1), .A4(new_n255_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n256_), .A2(KEYINPUT87), .A3(KEYINPUT1), .ZN(new_n259_));
  NOR2_X1   g058(.A1(G155gat), .A2(G162gat), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT1), .B1(new_n254_), .B2(new_n255_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT87), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n260_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n257_), .A2(new_n258_), .A3(new_n259_), .A4(new_n263_), .ZN(new_n264_));
  XOR2_X1   g063(.A(G141gat), .B(G148gat), .Z(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  OR3_X1    g065(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT2), .ZN(new_n268_));
  INV_X1    g067(.A(G141gat), .ZN(new_n269_));
  INV_X1    g068(.A(G148gat), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n268_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n267_), .A2(new_n271_), .A3(new_n272_), .A4(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n260_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n274_), .A2(new_n256_), .A3(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n266_), .A2(new_n276_), .ZN(new_n277_));
  XOR2_X1   g076(.A(KEYINPUT92), .B(KEYINPUT29), .Z(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT93), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G211gat), .B(G218gat), .ZN(new_n282_));
  INV_X1    g081(.A(G197gat), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n283_), .A2(G204gat), .ZN(new_n284_));
  OAI211_X1 g083(.A(new_n282_), .B(KEYINPUT21), .C1(KEYINPUT91), .C2(new_n284_), .ZN(new_n285_));
  XOR2_X1   g084(.A(G197gat), .B(G204gat), .Z(new_n286_));
  OR2_X1    g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n285_), .B(new_n286_), .C1(KEYINPUT21), .C2(new_n282_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n277_), .A2(KEYINPUT93), .A3(new_n278_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n281_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(G233gat), .ZN(new_n292_));
  NOR2_X1   g091(.A1(KEYINPUT90), .A2(G228gat), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(KEYINPUT90), .A2(G228gat), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n292_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n291_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n277_), .A2(KEYINPUT89), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT89), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n266_), .A2(new_n299_), .A3(new_n276_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n298_), .A2(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n296_), .B1(new_n301_), .B2(KEYINPUT29), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(new_n289_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G78gat), .B(G106gat), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  AND3_X1   g104(.A1(new_n297_), .A2(new_n303_), .A3(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n301_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT29), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  XOR2_X1   g108(.A(G22gat), .B(G50gat), .Z(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT28), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n309_), .B(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n305_), .B1(new_n303_), .B2(new_n297_), .ZN(new_n313_));
  OR3_X1    g112(.A1(new_n306_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n312_), .B1(new_n306_), .B2(new_n313_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT95), .ZN(new_n317_));
  INV_X1    g116(.A(new_n234_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n208_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n216_), .A2(KEYINPUT24), .A3(new_n224_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT83), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n319_), .B1(new_n322_), .B2(new_n225_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n318_), .B1(new_n323_), .B2(new_n221_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n289_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n317_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT20), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n208_), .B(KEYINPUT94), .C1(KEYINPUT24), .C2(new_n211_), .ZN(new_n328_));
  AND2_X1   g127(.A1(new_n328_), .A2(new_n320_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n208_), .B1(KEYINPUT24), .B2(new_n211_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT94), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n220_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT22), .B(G169gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(new_n210_), .ZN(new_n334_));
  AND2_X1   g133(.A1(new_n334_), .A2(new_n224_), .ZN(new_n335_));
  AOI22_X1  g134(.A1(new_n329_), .A2(new_n332_), .B1(new_n229_), .B2(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n327_), .B1(new_n336_), .B2(new_n325_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n235_), .A2(KEYINPUT95), .A3(new_n289_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n326_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G226gat), .A2(G233gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(KEYINPUT19), .ZN(new_n341_));
  OR2_X1    g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G8gat), .B(G36gat), .ZN(new_n343_));
  INV_X1    g142(.A(G92gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT18), .B(G64gat), .ZN(new_n346_));
  XOR2_X1   g145(.A(new_n345_), .B(new_n346_), .Z(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(KEYINPUT32), .ZN(new_n349_));
  INV_X1    g148(.A(new_n336_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n327_), .B1(new_n350_), .B2(new_n289_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n324_), .A2(new_n325_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(new_n341_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n342_), .A2(new_n349_), .A3(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n341_), .ZN(new_n356_));
  AND3_X1   g155(.A1(new_n351_), .A2(new_n356_), .A3(new_n352_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n357_), .B1(new_n339_), .B2(new_n341_), .ZN(new_n358_));
  OR2_X1    g157(.A1(new_n358_), .A2(new_n349_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G225gat), .A2(G233gat), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT4), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n299_), .B1(new_n266_), .B2(new_n276_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n276_), .ZN(new_n364_));
  AOI211_X1 g163(.A(KEYINPUT89), .B(new_n364_), .C1(new_n264_), .C2(new_n265_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n245_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n266_), .A2(new_n276_), .A3(new_n242_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n362_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(KEYINPUT4), .B1(new_n301_), .B2(new_n245_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n361_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT96), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  OAI211_X1 g171(.A(KEYINPUT96), .B(new_n361_), .C1(new_n368_), .C2(new_n369_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G1gat), .B(G29gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(G85gat), .ZN(new_n376_));
  XOR2_X1   g175(.A(KEYINPUT0), .B(G57gat), .Z(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n366_), .A2(new_n367_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n379_), .A2(new_n361_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT97), .ZN(new_n381_));
  AND3_X1   g180(.A1(new_n374_), .A2(new_n378_), .A3(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n378_), .B1(new_n374_), .B2(new_n381_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n355_), .B(new_n359_), .C1(new_n382_), .C2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n374_), .A2(new_n378_), .A3(new_n381_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT33), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n342_), .A2(new_n354_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(new_n347_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n342_), .A2(new_n348_), .A3(new_n354_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n366_), .A2(new_n361_), .A3(new_n367_), .ZN(new_n392_));
  OR2_X1    g191(.A1(new_n368_), .A2(new_n369_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n378_), .B1(new_n393_), .B2(new_n360_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n391_), .B1(new_n392_), .B2(new_n394_), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n374_), .A2(KEYINPUT33), .A3(new_n381_), .A4(new_n378_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n387_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n316_), .B1(new_n384_), .B2(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n382_), .A2(new_n383_), .ZN(new_n399_));
  OAI21_X1  g198(.A(KEYINPUT98), .B1(new_n358_), .B2(new_n348_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT98), .ZN(new_n401_));
  AND2_X1   g200(.A1(new_n339_), .A2(new_n341_), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n401_), .B(new_n347_), .C1(new_n402_), .C2(new_n357_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n400_), .A2(new_n390_), .A3(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(KEYINPUT27), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT27), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n389_), .A2(new_n406_), .A3(new_n390_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n405_), .A2(new_n407_), .ZN(new_n408_));
  AND3_X1   g207(.A1(new_n399_), .A2(new_n316_), .A3(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n251_), .B1(new_n398_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n250_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n248_), .B(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n316_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n412_), .A2(new_n399_), .A3(new_n413_), .A4(new_n408_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n410_), .A2(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G190gat), .B(G218gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G134gat), .B(G162gat), .ZN(new_n417_));
  XOR2_X1   g216(.A(new_n416_), .B(new_n417_), .Z(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(KEYINPUT36), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT35), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G29gat), .B(G36gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(G50gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT74), .B(G43gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  XOR2_X1   g223(.A(G85gat), .B(G92gat), .Z(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(KEYINPUT9), .ZN(new_n426_));
  XOR2_X1   g225(.A(KEYINPUT10), .B(G99gat), .Z(new_n427_));
  INV_X1    g226(.A(G106gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G99gat), .A2(G106gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT6), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT6), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n432_), .A2(G99gat), .A3(G106gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n431_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(G85gat), .ZN(new_n435_));
  OR3_X1    g234(.A1(new_n435_), .A2(new_n344_), .A3(KEYINPUT9), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n426_), .A2(new_n429_), .A3(new_n434_), .A4(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT8), .ZN(new_n438_));
  AND3_X1   g237(.A1(new_n431_), .A2(new_n433_), .A3(KEYINPUT66), .ZN(new_n439_));
  AOI21_X1  g238(.A(KEYINPUT66), .B1(new_n431_), .B2(new_n433_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(G99gat), .A2(G106gat), .ZN(new_n442_));
  AND2_X1   g241(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n443_));
  NOR2_X1   g242(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n442_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT67), .ZN(new_n446_));
  OAI22_X1  g245(.A1(KEYINPUT64), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n447_));
  AND3_X1   g246(.A1(new_n445_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n446_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n441_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n438_), .B1(new_n450_), .B2(new_n425_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n445_), .A2(new_n434_), .A3(new_n447_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n452_), .A2(new_n438_), .A3(new_n425_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT65), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT65), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n452_), .A2(new_n455_), .A3(new_n438_), .A4(new_n425_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n454_), .A2(new_n456_), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n424_), .B(new_n437_), .C1(new_n451_), .C2(new_n457_), .ZN(new_n458_));
  AND2_X1   g257(.A1(new_n422_), .A2(new_n423_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n422_), .A2(new_n423_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT15), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT15), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n424_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n437_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n450_), .A2(new_n425_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT8), .ZN(new_n468_));
  AND2_X1   g267(.A1(new_n454_), .A2(new_n456_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n466_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  OAI211_X1 g269(.A(new_n420_), .B(new_n458_), .C1(new_n465_), .C2(new_n470_), .ZN(new_n471_));
  XOR2_X1   g270(.A(KEYINPUT73), .B(KEYINPUT34), .Z(new_n472_));
  NAND2_X1  g271(.A1(G232gat), .A2(G233gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n471_), .A2(new_n474_), .ZN(new_n475_));
  AND2_X1   g274(.A1(new_n462_), .A2(new_n464_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n437_), .B1(new_n451_), .B2(new_n457_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n478_), .A2(KEYINPUT75), .A3(new_n458_), .ZN(new_n479_));
  OR2_X1    g278(.A1(new_n474_), .A2(KEYINPUT35), .ZN(new_n480_));
  AND3_X1   g279(.A1(new_n475_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n479_), .B1(new_n475_), .B2(new_n480_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n419_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n475_), .A2(new_n480_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n479_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n418_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n487_), .A2(KEYINPUT36), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n475_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n486_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  AOI211_X1 g289(.A(KEYINPUT76), .B(KEYINPUT37), .C1(new_n483_), .C2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(KEYINPUT76), .A2(KEYINPUT37), .ZN(new_n492_));
  NOR2_X1   g291(.A1(KEYINPUT76), .A2(KEYINPUT37), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  AND4_X1   g293(.A1(new_n490_), .A2(new_n483_), .A3(new_n492_), .A4(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n491_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(G57gat), .ZN(new_n498_));
  INV_X1    g297(.A(G64gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT11), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G57gat), .A2(G64gat), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n500_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT68), .ZN(new_n504_));
  INV_X1    g303(.A(G78gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(G71gat), .ZN(new_n506_));
  INV_X1    g305(.A(G71gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(G78gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  AND3_X1   g308(.A1(new_n503_), .A2(new_n504_), .A3(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n504_), .B1(new_n503_), .B2(new_n509_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n501_), .B1(new_n500_), .B2(new_n502_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NOR3_X1   g312(.A1(new_n510_), .A2(new_n511_), .A3(new_n513_), .ZN(new_n514_));
  AND2_X1   g313(.A1(G57gat), .A2(G64gat), .ZN(new_n515_));
  NOR2_X1   g314(.A1(G57gat), .A2(G64gat), .ZN(new_n516_));
  NOR3_X1   g315(.A1(new_n515_), .A2(new_n516_), .A3(KEYINPUT11), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G71gat), .B(G78gat), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT68), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n503_), .A2(new_n504_), .A3(new_n509_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n512_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n514_), .A2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G15gat), .B(G22gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G1gat), .A2(G8gat), .ZN(new_n524_));
  AND3_X1   g323(.A1(new_n524_), .A2(KEYINPUT77), .A3(KEYINPUT14), .ZN(new_n525_));
  AOI21_X1  g324(.A(KEYINPUT77), .B1(new_n524_), .B2(KEYINPUT14), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n523_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  XOR2_X1   g326(.A(G1gat), .B(G8gat), .Z(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n522_), .B(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G231gat), .A2(G233gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT69), .ZN(new_n534_));
  XOR2_X1   g333(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n535_));
  XNOR2_X1  g334(.A(G127gat), .B(G155gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  XOR2_X1   g336(.A(G183gat), .B(G211gat), .Z(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT17), .ZN(new_n540_));
  OR2_X1    g339(.A1(new_n539_), .A2(KEYINPUT17), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n534_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n540_), .B(KEYINPUT79), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n533_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n497_), .A2(new_n545_), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n415_), .A2(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n461_), .A2(new_n530_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n548_), .B1(new_n476_), .B2(new_n530_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G229gat), .A2(G233gat), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n548_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n461_), .A2(new_n530_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n550_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n551_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G113gat), .B(G141gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G169gat), .B(G197gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n558_), .A2(KEYINPUT81), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT81), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n564_), .B1(new_n557_), .B2(new_n561_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n558_), .A2(KEYINPUT80), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT80), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n557_), .A2(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n567_), .A2(new_n561_), .A3(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n566_), .A2(new_n570_), .ZN(new_n571_));
  AND3_X1   g370(.A1(new_n477_), .A2(KEYINPUT12), .A3(new_n522_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n513_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n519_), .A2(new_n512_), .A3(new_n520_), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n573_), .A2(KEYINPUT69), .A3(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(KEYINPUT69), .B1(new_n573_), .B2(new_n574_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(KEYINPUT12), .B1(new_n477_), .B2(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n572_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G230gat), .A2(G233gat), .ZN(new_n580_));
  OAI211_X1 g379(.A(KEYINPUT70), .B(new_n580_), .C1(new_n477_), .C2(new_n577_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n425_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n445_), .A2(new_n447_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(KEYINPUT67), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n445_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n583_), .B1(new_n587_), .B2(new_n441_), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n454_), .B(new_n456_), .C1(new_n588_), .C2(new_n438_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT69), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n590_), .B1(new_n514_), .B2(new_n521_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n573_), .A2(KEYINPUT69), .A3(new_n574_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n589_), .A2(new_n437_), .A3(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(KEYINPUT70), .B1(new_n594_), .B2(new_n580_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n579_), .B1(new_n582_), .B2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n594_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n593_), .B1(new_n589_), .B2(new_n437_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n596_), .B1(new_n580_), .B2(new_n599_), .ZN(new_n600_));
  XOR2_X1   g399(.A(G176gat), .B(G204gat), .Z(new_n601_));
  XNOR2_X1  g400(.A(G120gat), .B(G148gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  OR2_X1    g404(.A1(new_n605_), .A2(KEYINPUT71), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n600_), .B(new_n606_), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n607_), .A2(KEYINPUT13), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(KEYINPUT13), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n547_), .A2(new_n571_), .A3(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(G1gat), .ZN(new_n613_));
  INV_X1    g412(.A(new_n399_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n612_), .A2(new_n613_), .A3(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT38), .ZN(new_n616_));
  INV_X1    g415(.A(new_n571_), .ZN(new_n617_));
  NOR3_X1   g416(.A1(new_n610_), .A2(new_n617_), .A3(new_n545_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT99), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n483_), .A2(new_n490_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n620_), .B1(new_n410_), .B2(new_n414_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n622_), .B(KEYINPUT100), .Z(new_n623_));
  OAI21_X1  g422(.A(G1gat), .B1(new_n623_), .B2(new_n399_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n616_), .A2(new_n624_), .ZN(G1324gat));
  INV_X1    g424(.A(G8gat), .ZN(new_n626_));
  INV_X1    g425(.A(new_n408_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n626_), .B1(new_n622_), .B2(new_n627_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n628_), .B(KEYINPUT39), .Z(new_n629_));
  NAND3_X1  g428(.A1(new_n612_), .A2(new_n626_), .A3(new_n627_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g431(.A(G15gat), .B1(new_n623_), .B2(new_n251_), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n633_), .B(KEYINPUT41), .Z(new_n634_));
  INV_X1    g433(.A(G15gat), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n612_), .A2(new_n635_), .A3(new_n412_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n634_), .A2(new_n636_), .ZN(G1326gat));
  OAI21_X1  g436(.A(G22gat), .B1(new_n623_), .B2(new_n413_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT42), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n413_), .A2(G22gat), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT101), .Z(new_n641_));
  NAND2_X1  g440(.A1(new_n612_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n639_), .A2(new_n642_), .ZN(G1327gat));
  INV_X1    g442(.A(new_n620_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n644_), .B1(new_n410_), .B2(new_n414_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n545_), .ZN(new_n646_));
  NOR3_X1   g445(.A1(new_n610_), .A2(new_n617_), .A3(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n648_), .A2(G29gat), .A3(new_n399_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n415_), .A2(new_n497_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT102), .ZN(new_n652_));
  AOI21_X1  g451(.A(KEYINPUT43), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n496_), .B1(new_n410_), .B2(new_n414_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT43), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n654_), .A2(KEYINPUT102), .A3(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n647_), .B1(new_n653_), .B2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(KEYINPUT103), .A2(KEYINPUT44), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT103), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT44), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n657_), .A2(new_n658_), .A3(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n651_), .A2(new_n652_), .A3(KEYINPUT43), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n655_), .B1(new_n654_), .B2(KEYINPUT102), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n665_), .A2(new_n659_), .A3(new_n660_), .A4(new_n647_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n399_), .B1(new_n662_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(G29gat), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n650_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT104), .ZN(G1328gat));
  NOR3_X1   g469(.A1(new_n648_), .A2(G36gat), .A3(new_n408_), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n671_), .B(KEYINPUT45), .Z(new_n672_));
  AOI21_X1  g471(.A(new_n408_), .B1(new_n662_), .B2(new_n666_), .ZN(new_n673_));
  INV_X1    g472(.A(G36gat), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n672_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT105), .ZN(new_n676_));
  XNOR2_X1  g475(.A(KEYINPUT106), .B(KEYINPUT46), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n675_), .A2(new_n676_), .A3(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n677_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n678_), .A2(new_n679_), .ZN(G1329gat));
  INV_X1    g479(.A(G43gat), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n662_), .A2(new_n666_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n681_), .B1(new_n682_), .B2(new_n412_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT47), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n648_), .A2(G43gat), .A3(new_n251_), .ZN(new_n685_));
  OR3_X1    g484(.A1(new_n683_), .A2(new_n684_), .A3(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n684_), .B1(new_n683_), .B2(new_n685_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(G1330gat));
  INV_X1    g487(.A(G50gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n689_), .B1(new_n682_), .B2(new_n316_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT107), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n648_), .A2(G50gat), .A3(new_n413_), .ZN(new_n692_));
  OR3_X1    g491(.A1(new_n690_), .A2(new_n691_), .A3(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n691_), .B1(new_n690_), .B2(new_n692_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(G1331gat));
  NOR2_X1   g494(.A1(new_n611_), .A2(new_n571_), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n621_), .A2(new_n646_), .A3(new_n696_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n697_), .A2(G57gat), .A3(new_n614_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT108), .Z(new_n699_));
  NAND2_X1  g498(.A1(new_n547_), .A2(new_n696_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n498_), .B1(new_n700_), .B2(new_n399_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT109), .Z(G1332gat));
  AOI21_X1  g502(.A(new_n499_), .B1(new_n697_), .B2(new_n627_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(KEYINPUT110), .B(KEYINPUT48), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n704_), .B(new_n705_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n408_), .A2(G64gat), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT111), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n706_), .B1(new_n700_), .B2(new_n708_), .ZN(G1333gat));
  AOI21_X1  g508(.A(new_n507_), .B1(new_n697_), .B2(new_n412_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT49), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n700_), .A2(G71gat), .A3(new_n251_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT112), .ZN(G1334gat));
  AOI21_X1  g513(.A(new_n505_), .B1(new_n697_), .B2(new_n316_), .ZN(new_n715_));
  XOR2_X1   g514(.A(new_n715_), .B(KEYINPUT50), .Z(new_n716_));
  NAND2_X1  g515(.A1(new_n316_), .A2(new_n505_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n716_), .B1(new_n700_), .B2(new_n717_), .ZN(G1335gat));
  NOR3_X1   g517(.A1(new_n611_), .A2(new_n571_), .A3(new_n646_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n645_), .A2(new_n719_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n435_), .B1(new_n720_), .B2(new_n399_), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT113), .Z(new_n722_));
  NAND2_X1  g521(.A1(new_n665_), .A2(new_n719_), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n723_), .A2(new_n435_), .A3(new_n399_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n722_), .A2(new_n724_), .ZN(G1336gat));
  INV_X1    g524(.A(new_n720_), .ZN(new_n726_));
  AOI21_X1  g525(.A(G92gat), .B1(new_n726_), .B2(new_n627_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n723_), .A2(new_n344_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n727_), .B1(new_n728_), .B2(new_n627_), .ZN(G1337gat));
  OAI21_X1  g528(.A(G99gat), .B1(new_n723_), .B2(new_n251_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n726_), .A2(new_n412_), .A3(new_n427_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n730_), .A2(new_n731_), .A3(new_n732_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n733_), .B(new_n734_), .Z(G1338gat));
  OAI21_X1  g534(.A(G106gat), .B1(new_n723_), .B2(new_n413_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT52), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  OAI211_X1 g537(.A(KEYINPUT52), .B(G106gat), .C1(new_n723_), .C2(new_n413_), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n720_), .A2(G106gat), .A3(new_n413_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT115), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n738_), .A2(new_n739_), .A3(new_n741_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g542(.A1(new_n546_), .A2(new_n617_), .A3(new_n611_), .ZN(new_n744_));
  OR2_X1    g543(.A1(new_n744_), .A2(KEYINPUT54), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(KEYINPUT54), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT118), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT116), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT55), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n596_), .A2(new_n749_), .A3(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(new_n596_), .B2(new_n749_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n580_), .B1(new_n579_), .B2(new_n594_), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n751_), .A2(new_n752_), .A3(new_n753_), .ZN(new_n754_));
  OAI21_X1  g553(.A(KEYINPUT56), .B1(new_n754_), .B2(new_n605_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n555_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n756_));
  AOI211_X1 g555(.A(new_n562_), .B(new_n756_), .C1(new_n549_), .C2(new_n555_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n757_), .B1(new_n563_), .B2(new_n565_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n605_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n600_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n477_), .A2(KEYINPUT12), .A3(new_n522_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n762_), .B1(new_n598_), .B2(KEYINPUT12), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n594_), .A2(new_n580_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT70), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n763_), .B1(new_n766_), .B2(new_n581_), .ZN(new_n767_));
  OAI21_X1  g566(.A(KEYINPUT55), .B1(new_n767_), .B2(KEYINPUT116), .ZN(new_n768_));
  INV_X1    g567(.A(new_n753_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n596_), .A2(new_n749_), .A3(new_n750_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n768_), .A2(new_n769_), .A3(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT56), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n771_), .A2(new_n772_), .A3(new_n759_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n755_), .A2(new_n758_), .A3(new_n761_), .A4(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT58), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n748_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n771_), .A2(new_n772_), .A3(new_n759_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n772_), .B1(new_n771_), .B2(new_n759_), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n777_), .A2(new_n778_), .A3(new_n760_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n779_), .A2(KEYINPUT118), .A3(KEYINPUT58), .A4(new_n758_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n496_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n776_), .A2(new_n780_), .A3(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT117), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n755_), .A2(new_n571_), .A3(new_n761_), .A4(new_n773_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n607_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n758_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n783_), .B1(new_n787_), .B2(new_n644_), .ZN(new_n788_));
  AOI211_X1 g587(.A(KEYINPUT117), .B(new_n620_), .C1(new_n784_), .C2(new_n786_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT57), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n782_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n787_), .A2(new_n644_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n793_), .A2(new_n791_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n792_), .A2(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n747_), .B1(new_n796_), .B2(new_n545_), .ZN(new_n797_));
  NOR4_X1   g596(.A1(new_n251_), .A2(new_n399_), .A3(new_n316_), .A4(new_n627_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n797_), .A2(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(G113gat), .B1(new_n800_), .B2(new_n571_), .ZN(new_n801_));
  INV_X1    g600(.A(G113gat), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT121), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n802_), .B1(new_n571_), .B2(new_n803_), .ZN(new_n804_));
  NOR3_X1   g603(.A1(new_n788_), .A2(new_n789_), .A3(KEYINPUT57), .ZN(new_n805_));
  OAI21_X1  g604(.A(KEYINPUT119), .B1(new_n805_), .B2(new_n782_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n793_), .A2(KEYINPUT117), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n787_), .A2(new_n783_), .A3(new_n644_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n807_), .A2(new_n791_), .A3(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT119), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n776_), .A2(new_n780_), .A3(new_n781_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n809_), .A2(new_n810_), .A3(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n806_), .A2(new_n795_), .A3(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n747_), .B1(new_n813_), .B2(new_n545_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n799_), .A2(KEYINPUT59), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT59), .ZN(new_n817_));
  OAI221_X1 g616(.A(KEYINPUT120), .B1(new_n814_), .B2(new_n816_), .C1(new_n800_), .C2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT120), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n814_), .A2(new_n816_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n796_), .A2(new_n545_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n747_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n817_), .B1(new_n823_), .B2(new_n798_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n819_), .B1(new_n820_), .B2(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n804_), .B1(new_n818_), .B2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n803_), .A2(new_n802_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n801_), .B1(new_n826_), .B2(new_n827_), .ZN(G1340gat));
  INV_X1    g627(.A(G120gat), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n829_), .B1(new_n611_), .B2(KEYINPUT60), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n800_), .B(new_n830_), .C1(KEYINPUT60), .C2(new_n829_), .ZN(new_n831_));
  OR3_X1    g630(.A1(new_n820_), .A2(new_n824_), .A3(new_n611_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n831_), .B1(new_n833_), .B2(new_n829_), .ZN(G1341gat));
  AOI21_X1  g633(.A(G127gat), .B1(new_n800_), .B2(new_n646_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n545_), .B1(new_n818_), .B2(new_n825_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n835_), .B1(new_n836_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g636(.A(G134gat), .B1(new_n800_), .B2(new_n620_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n496_), .B1(new_n818_), .B2(new_n825_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n838_), .B1(new_n839_), .B2(G134gat), .ZN(G1343gat));
  NOR2_X1   g639(.A1(new_n412_), .A2(new_n413_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n627_), .A2(new_n399_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n823_), .A2(new_n841_), .A3(new_n842_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n843_), .A2(new_n617_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(new_n269_), .ZN(G1344gat));
  NOR2_X1   g644(.A1(new_n843_), .A2(new_n611_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(new_n270_), .ZN(G1345gat));
  NAND4_X1  g646(.A1(new_n823_), .A2(new_n646_), .A3(new_n841_), .A4(new_n842_), .ZN(new_n848_));
  OR2_X1    g647(.A1(new_n848_), .A2(KEYINPUT122), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(KEYINPUT122), .ZN(new_n850_));
  XNOR2_X1  g649(.A(KEYINPUT61), .B(G155gat), .ZN(new_n851_));
  AND3_X1   g650(.A1(new_n849_), .A2(new_n850_), .A3(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n851_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n852_), .A2(new_n853_), .ZN(G1346gat));
  NOR2_X1   g653(.A1(new_n843_), .A2(new_n644_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n855_), .A2(G162gat), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n843_), .A2(new_n496_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n856_), .B1(G162gat), .B2(new_n857_), .ZN(G1347gat));
  NOR2_X1   g657(.A1(new_n251_), .A2(new_n614_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n859_), .A2(new_n413_), .A3(new_n627_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n812_), .A2(new_n795_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n810_), .B1(new_n809_), .B2(new_n811_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n545_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n860_), .B1(new_n863_), .B2(new_n822_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n209_), .B1(new_n864_), .B2(new_n571_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT62), .ZN(new_n866_));
  OAI21_X1  g665(.A(KEYINPUT124), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n860_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n794_), .B1(new_n792_), .B2(new_n810_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n646_), .B1(new_n869_), .B2(new_n806_), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n571_), .B(new_n868_), .C1(new_n870_), .C2(new_n747_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n871_), .A2(new_n866_), .A3(G169gat), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT123), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n871_), .A2(KEYINPUT123), .A3(new_n866_), .A4(G169gat), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT124), .ZN(new_n876_));
  NOR3_X1   g675(.A1(new_n814_), .A2(new_n617_), .A3(new_n860_), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n876_), .B(KEYINPUT62), .C1(new_n877_), .C2(new_n209_), .ZN(new_n878_));
  NAND4_X1  g677(.A1(new_n867_), .A2(new_n874_), .A3(new_n875_), .A4(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n333_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(G1348gat));
  NOR2_X1   g680(.A1(new_n797_), .A2(new_n860_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n882_), .A2(G176gat), .A3(new_n610_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT125), .ZN(new_n884_));
  AND2_X1   g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n883_), .A2(new_n884_), .ZN(new_n886_));
  AOI21_X1  g685(.A(G176gat), .B1(new_n864_), .B2(new_n610_), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n885_), .A2(new_n886_), .A3(new_n887_), .ZN(G1349gat));
  AOI21_X1  g687(.A(G183gat), .B1(new_n882_), .B2(new_n646_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n545_), .A2(new_n218_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n889_), .B1(new_n864_), .B2(new_n890_), .ZN(G1350gat));
  INV_X1    g690(.A(new_n864_), .ZN(new_n892_));
  OAI21_X1  g691(.A(G190gat), .B1(new_n892_), .B2(new_n496_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n864_), .A2(new_n219_), .A3(new_n620_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(G1351gat));
  NOR2_X1   g694(.A1(new_n614_), .A2(new_n413_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n896_), .A2(new_n251_), .A3(new_n627_), .ZN(new_n897_));
  OAI21_X1  g696(.A(KEYINPUT126), .B1(new_n797_), .B2(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT126), .ZN(new_n899_));
  INV_X1    g698(.A(new_n897_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n823_), .A2(new_n899_), .A3(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n898_), .A2(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(new_n571_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g703(.A1(new_n902_), .A2(new_n610_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g705(.A(new_n545_), .B1(new_n898_), .B2(new_n901_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n907_), .A2(new_n908_), .ZN(new_n909_));
  XOR2_X1   g708(.A(KEYINPUT63), .B(G211gat), .Z(new_n910_));
  AOI211_X1 g709(.A(new_n545_), .B(new_n910_), .C1(new_n898_), .C2(new_n901_), .ZN(new_n911_));
  OAI21_X1  g710(.A(KEYINPUT127), .B1(new_n909_), .B2(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n910_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n907_), .A2(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT127), .ZN(new_n915_));
  OAI211_X1 g714(.A(new_n914_), .B(new_n915_), .C1(new_n907_), .C2(new_n908_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n912_), .A2(new_n916_), .ZN(G1354gat));
  AOI21_X1  g716(.A(G218gat), .B1(new_n902_), .B2(new_n620_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n496_), .B1(new_n898_), .B2(new_n901_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n918_), .B1(G218gat), .B2(new_n919_), .ZN(G1355gat));
endmodule


