//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 1 1 0 0 1 1 0 0 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 0 0 0 0 0 1 0 1 1 0 0 0 1 0 0 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n931_, new_n932_, new_n934_,
    new_n935_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n943_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n953_, new_n954_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n966_, new_n967_, new_n969_, new_n970_, new_n972_,
    new_n973_, new_n975_, new_n976_, new_n977_, new_n979_, new_n980_,
    new_n981_, new_n982_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n992_, new_n993_, new_n994_;
  INV_X1    g000(.A(KEYINPUT71), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT70), .ZN(new_n203_));
  XOR2_X1   g002(.A(KEYINPUT10), .B(G99gat), .Z(new_n204_));
  INV_X1    g003(.A(G106gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  XOR2_X1   g005(.A(G85gat), .B(G92gat), .Z(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT9), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G99gat), .A2(G106gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT6), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT6), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n211_), .A2(G99gat), .A3(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT9), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(G85gat), .A3(G92gat), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n206_), .A2(new_n208_), .A3(new_n213_), .A4(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT8), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n211_), .B1(G99gat), .B2(G106gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n209_), .A2(KEYINPUT6), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT65), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n210_), .A2(new_n212_), .A3(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(G99gat), .A2(G106gat), .ZN(new_n223_));
  AND2_X1   g022(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n224_));
  NOR2_X1   g023(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n223_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  OAI22_X1  g025(.A1(KEYINPUT64), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n220_), .A2(new_n222_), .A3(new_n226_), .A4(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n217_), .B1(new_n228_), .B2(new_n207_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n207_), .A2(new_n217_), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n226_), .A2(new_n227_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n230_), .B1(new_n231_), .B2(new_n213_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n216_), .B1(new_n229_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT66), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G29gat), .B(G36gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G43gat), .B(G50gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  OAI211_X1 g037(.A(KEYINPUT66), .B(new_n216_), .C1(new_n229_), .C2(new_n232_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n235_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G232gat), .A2(G233gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT34), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT35), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT69), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n244_), .B1(new_n242_), .B2(KEYINPUT35), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n238_), .B(KEYINPUT15), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n245_), .B1(new_n233_), .B2(new_n246_), .ZN(new_n247_));
  AND3_X1   g046(.A1(new_n240_), .A2(new_n243_), .A3(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n243_), .B1(new_n240_), .B2(new_n247_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n203_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n240_), .A2(new_n247_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n243_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n240_), .A2(new_n243_), .A3(new_n247_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n253_), .A2(KEYINPUT70), .A3(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n250_), .A2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G190gat), .B(G218gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G134gat), .B(G162gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  XOR2_X1   g058(.A(new_n259_), .B(KEYINPUT36), .Z(new_n260_));
  NAND2_X1  g059(.A1(new_n256_), .A2(new_n260_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n259_), .A2(KEYINPUT36), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n253_), .A2(new_n262_), .A3(new_n254_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT37), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n261_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n262_), .ZN(new_n268_));
  NOR3_X1   g067(.A1(new_n248_), .A2(new_n249_), .A3(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n260_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n270_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n271_));
  OAI21_X1  g070(.A(KEYINPUT37), .B1(new_n269_), .B2(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n202_), .B1(new_n267_), .B2(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n270_), .B1(new_n250_), .B2(new_n255_), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n272_), .B(new_n202_), .C1(new_n274_), .C2(new_n265_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n273_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(G230gat), .ZN(new_n278_));
  INV_X1    g077(.A(G233gat), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G57gat), .B(G64gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT11), .ZN(new_n282_));
  XOR2_X1   g081(.A(G71gat), .B(G78gat), .Z(new_n283_));
  OR2_X1    g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n281_), .A2(KEYINPUT11), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n282_), .A2(new_n283_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n284_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  AND3_X1   g086(.A1(new_n235_), .A2(new_n287_), .A3(new_n239_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n287_), .B1(new_n235_), .B2(new_n239_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n280_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  XOR2_X1   g089(.A(G120gat), .B(G148gat), .Z(new_n291_));
  XNOR2_X1  g090(.A(G176gat), .B(G204gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n287_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n233_), .A2(KEYINPUT12), .A3(new_n296_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n297_), .B1(new_n289_), .B2(KEYINPUT12), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n235_), .A2(new_n287_), .A3(new_n239_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n299_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n300_));
  OAI211_X1 g099(.A(new_n290_), .B(new_n295_), .C1(new_n298_), .C2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT68), .ZN(new_n302_));
  INV_X1    g101(.A(new_n297_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n232_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n207_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n226_), .A2(new_n227_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n221_), .B1(new_n210_), .B2(new_n212_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n305_), .B1(new_n308_), .B2(new_n222_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n304_), .B1(new_n309_), .B2(new_n217_), .ZN(new_n310_));
  AOI21_X1  g109(.A(KEYINPUT66), .B1(new_n310_), .B2(new_n216_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n239_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n296_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT12), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n303_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n288_), .A2(new_n280_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT68), .ZN(new_n318_));
  NAND4_X1  g117(.A1(new_n317_), .A2(new_n318_), .A3(new_n290_), .A4(new_n295_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n302_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n317_), .A2(new_n290_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n295_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n320_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT13), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n320_), .A2(KEYINPUT13), .A3(new_n323_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G127gat), .B(G155gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT16), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G183gat), .B(G211gat), .ZN(new_n331_));
  XOR2_X1   g130(.A(new_n330_), .B(new_n331_), .Z(new_n332_));
  AND2_X1   g131(.A1(G231gat), .A2(G233gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n287_), .B(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT72), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G15gat), .B(G22gat), .ZN(new_n337_));
  INV_X1    g136(.A(G1gat), .ZN(new_n338_));
  INV_X1    g137(.A(G8gat), .ZN(new_n339_));
  OAI21_X1  g138(.A(KEYINPUT14), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n337_), .A2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G1gat), .B(G8gat), .ZN(new_n342_));
  XOR2_X1   g141(.A(new_n341_), .B(new_n342_), .Z(new_n343_));
  NAND2_X1  g142(.A1(new_n334_), .A2(new_n335_), .ZN(new_n344_));
  AND3_X1   g143(.A1(new_n336_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n343_), .B1(new_n336_), .B2(new_n344_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n332_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT73), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n348_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n332_), .ZN(new_n350_));
  AOI22_X1  g149(.A1(KEYINPUT17), .A2(new_n347_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n334_), .B(new_n335_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n343_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n336_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n355_));
  AOI21_X1  g154(.A(KEYINPUT73), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT17), .ZN(new_n357_));
  NOR3_X1   g156(.A1(new_n356_), .A2(new_n357_), .A3(new_n332_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n351_), .A2(new_n358_), .ZN(new_n359_));
  NOR3_X1   g158(.A1(new_n277_), .A2(new_n328_), .A3(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT74), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G1gat), .B(G29gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(G85gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT0), .B(G57gat), .ZN(new_n365_));
  XOR2_X1   g164(.A(new_n364_), .B(new_n365_), .Z(new_n366_));
  NAND2_X1  g165(.A1(G225gat), .A2(G233gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(KEYINPUT92), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  XOR2_X1   g168(.A(G127gat), .B(G134gat), .Z(new_n370_));
  XOR2_X1   g169(.A(G113gat), .B(G120gat), .Z(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G127gat), .B(G134gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G113gat), .B(G120gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n372_), .A2(KEYINPUT83), .A3(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(KEYINPUT83), .B1(new_n372_), .B2(new_n375_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(G155gat), .ZN(new_n379_));
  INV_X1    g178(.A(G162gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G155gat), .A2(G162gat), .ZN(new_n382_));
  AND2_X1   g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT86), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G141gat), .A2(G148gat), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT2), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n390_));
  INV_X1    g189(.A(G141gat), .ZN(new_n391_));
  INV_X1    g190(.A(G148gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n389_), .B(new_n390_), .C1(new_n393_), .C2(KEYINPUT3), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n383_), .B1(new_n386_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT85), .ZN(new_n396_));
  NAND3_X1  g195(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(new_n387_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT84), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n399_), .B1(G141gat), .B2(G148gat), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n391_), .A2(new_n392_), .A3(KEYINPUT84), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n398_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT1), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n381_), .A2(new_n403_), .A3(new_n382_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n396_), .B1(new_n402_), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n401_), .A2(new_n400_), .ZN(new_n406_));
  AND2_X1   g205(.A1(new_n397_), .A2(new_n387_), .ZN(new_n407_));
  AND4_X1   g206(.A1(new_n396_), .A2(new_n406_), .A3(new_n404_), .A4(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n395_), .B1(new_n405_), .B2(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(KEYINPUT4), .B1(new_n378_), .B2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n378_), .A2(new_n409_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n372_), .A2(new_n375_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n411_), .B1(new_n409_), .B2(new_n413_), .ZN(new_n414_));
  AOI211_X1 g213(.A(new_n369_), .B(new_n410_), .C1(new_n414_), .C2(KEYINPUT4), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n369_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n366_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT97), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n414_), .A2(KEYINPUT4), .ZN(new_n420_));
  INV_X1    g219(.A(new_n410_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n420_), .A2(new_n368_), .A3(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n366_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n422_), .A2(new_n423_), .A3(new_n416_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n418_), .A2(new_n419_), .A3(new_n424_), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n422_), .A2(KEYINPUT97), .A3(new_n423_), .A4(new_n416_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G22gat), .B(G50gat), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n406_), .A2(new_n404_), .A3(new_n407_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT85), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n406_), .A2(new_n404_), .A3(new_n407_), .A4(new_n396_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT29), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n434_), .A2(new_n435_), .A3(new_n395_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(KEYINPUT28), .ZN(new_n437_));
  INV_X1    g236(.A(G228gat), .ZN(new_n438_));
  OR2_X1    g237(.A1(new_n438_), .A2(KEYINPUT88), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(KEYINPUT88), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n279_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n409_), .A2(KEYINPUT29), .ZN(new_n443_));
  XOR2_X1   g242(.A(G211gat), .B(G218gat), .Z(new_n444_));
  NOR2_X1   g243(.A1(G197gat), .A2(G204gat), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G197gat), .A2(G204gat), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n444_), .A2(KEYINPUT21), .A3(new_n446_), .A4(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n446_), .A2(KEYINPUT21), .A3(new_n447_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT21), .ZN(new_n450_));
  AND2_X1   g249(.A1(G197gat), .A2(G204gat), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n450_), .B1(new_n451_), .B2(new_n445_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G211gat), .B(G218gat), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n449_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n448_), .A2(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n442_), .B1(new_n443_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT89), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n448_), .A2(new_n454_), .A3(KEYINPUT89), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n458_), .A2(new_n459_), .A3(new_n442_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n435_), .B1(new_n434_), .B2(new_n395_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(G78gat), .B1(new_n456_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n455_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n441_), .B1(new_n461_), .B2(new_n464_), .ZN(new_n465_));
  AND3_X1   g264(.A1(new_n448_), .A2(new_n454_), .A3(KEYINPUT89), .ZN(new_n466_));
  AOI21_X1  g265(.A(KEYINPUT89), .B1(new_n448_), .B2(new_n454_), .ZN(new_n467_));
  NOR3_X1   g266(.A1(new_n466_), .A2(new_n467_), .A3(new_n441_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(new_n443_), .ZN(new_n469_));
  INV_X1    g268(.A(G78gat), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n465_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n463_), .A2(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(KEYINPUT87), .B1(new_n472_), .B2(new_n205_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n463_), .A2(G106gat), .A3(new_n471_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n437_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT87), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n465_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n470_), .B1(new_n465_), .B2(new_n469_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n205_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  AND4_X1   g278(.A1(new_n476_), .A2(new_n479_), .A3(new_n437_), .A4(new_n474_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n430_), .B1(new_n475_), .B2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n479_), .A2(new_n476_), .A3(new_n474_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n437_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n473_), .A2(new_n437_), .A3(new_n474_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n484_), .A2(new_n485_), .A3(new_n429_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n428_), .B1(new_n481_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G226gat), .A2(G233gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(KEYINPUT19), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n466_), .A2(new_n467_), .ZN(new_n491_));
  INV_X1    g290(.A(G169gat), .ZN(new_n492_));
  INV_X1    g291(.A(G176gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G169gat), .A2(G176gat), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n494_), .A2(KEYINPUT24), .A3(new_n495_), .ZN(new_n496_));
  OR3_X1    g295(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n497_));
  AND2_X1   g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(KEYINPUT25), .B(G183gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(KEYINPUT26), .B(G190gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  AND2_X1   g300(.A1(G183gat), .A2(G190gat), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT23), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT78), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT78), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT23), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n502_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G183gat), .A2(G190gat), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n508_), .A2(KEYINPUT23), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n498_), .B(new_n501_), .C1(new_n507_), .C2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT80), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT22), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(G169gat), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n492_), .A2(KEYINPUT22), .ZN(new_n514_));
  AOI21_X1  g313(.A(KEYINPUT79), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(KEYINPUT79), .B1(new_n492_), .B2(KEYINPUT22), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(new_n493_), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n511_), .B(new_n495_), .C1(new_n515_), .C2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n504_), .A2(new_n506_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(new_n502_), .ZN(new_n520_));
  INV_X1    g319(.A(G183gat), .ZN(new_n521_));
  INV_X1    g320(.A(G190gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n508_), .A2(new_n503_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n520_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n518_), .A2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT22), .B(G169gat), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n493_), .B(new_n516_), .C1(new_n527_), .C2(KEYINPUT79), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n511_), .B1(new_n528_), .B2(new_n495_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n510_), .B1(new_n526_), .B2(new_n529_), .ZN(new_n530_));
  OR2_X1    g329(.A1(new_n491_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT20), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n523_), .B1(new_n507_), .B2(new_n509_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n495_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n534_), .B1(new_n527_), .B2(new_n493_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT90), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n500_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT26), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n539_), .A2(G190gat), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n522_), .A2(KEYINPUT26), .ZN(new_n541_));
  OAI21_X1  g340(.A(KEYINPUT90), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  AND3_X1   g341(.A1(new_n538_), .A2(new_n542_), .A3(new_n499_), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n520_), .A2(new_n524_), .A3(new_n496_), .A4(new_n497_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n536_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n532_), .B1(new_n545_), .B2(new_n455_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n490_), .B1(new_n531_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(G8gat), .B(G36gat), .Z(new_n549_));
  XNOR2_X1  g348(.A(G64gat), .B(G92gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(KEYINPUT78), .B(KEYINPUT23), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n524_), .B1(new_n555_), .B2(new_n508_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n496_), .A2(new_n497_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n538_), .A2(new_n542_), .A3(new_n499_), .ZN(new_n559_));
  AOI22_X1  g358(.A1(new_n558_), .A2(new_n559_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n560_));
  AOI211_X1 g359(.A(new_n532_), .B(new_n489_), .C1(new_n560_), .C2(new_n464_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n491_), .A2(new_n530_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n548_), .A2(new_n554_), .A3(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n563_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n553_), .B1(new_n565_), .B2(new_n547_), .ZN(new_n566_));
  AOI21_X1  g365(.A(KEYINPUT27), .B1(new_n564_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT94), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n455_), .B1(new_n545_), .B2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n560_), .A2(KEYINPUT94), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n532_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  AOI22_X1  g370(.A1(new_n571_), .A2(KEYINPUT95), .B1(new_n491_), .B2(new_n530_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n464_), .B1(new_n560_), .B2(KEYINPUT94), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n545_), .A2(new_n568_), .ZN(new_n574_));
  OAI21_X1  g373(.A(KEYINPUT20), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT95), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n490_), .B1(new_n572_), .B2(new_n577_), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n531_), .A2(new_n490_), .A3(new_n546_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n553_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n564_), .A2(KEYINPUT27), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n567_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  AND3_X1   g381(.A1(new_n484_), .A2(new_n485_), .A3(new_n429_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n429_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT33), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n418_), .A2(KEYINPUT93), .A3(new_n586_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n564_), .A2(new_n566_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n410_), .B1(new_n414_), .B2(KEYINPUT4), .ZN(new_n589_));
  OR2_X1    g388(.A1(new_n589_), .A2(new_n368_), .ZN(new_n590_));
  OAI211_X1 g389(.A(new_n590_), .B(new_n423_), .C1(new_n414_), .C2(new_n369_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n586_), .A2(KEYINPUT93), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n366_), .B(new_n592_), .C1(new_n415_), .C2(new_n417_), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n587_), .A2(new_n588_), .A3(new_n591_), .A4(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT96), .ZN(new_n595_));
  OAI211_X1 g394(.A(KEYINPUT95), .B(KEYINPUT20), .C1(new_n573_), .C2(new_n574_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n577_), .A2(new_n562_), .A3(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n579_), .B1(new_n597_), .B2(new_n489_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n554_), .A2(KEYINPUT32), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n595_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n599_), .ZN(new_n601_));
  OAI211_X1 g400(.A(KEYINPUT96), .B(new_n601_), .C1(new_n578_), .C2(new_n579_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n548_), .A2(new_n563_), .A3(new_n599_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n425_), .A2(new_n426_), .A3(new_n604_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n594_), .B1(new_n603_), .B2(new_n605_), .ZN(new_n606_));
  AOI22_X1  g405(.A1(new_n487_), .A2(new_n582_), .B1(new_n585_), .B2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(G227gat), .A2(G233gat), .ZN(new_n608_));
  INV_X1    g407(.A(G15gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(G71gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(G99gat), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT30), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n530_), .A2(new_n614_), .ZN(new_n615_));
  OAI211_X1 g414(.A(new_n510_), .B(KEYINPUT30), .C1(new_n526_), .C2(new_n529_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(KEYINPUT81), .B(G43gat), .ZN(new_n617_));
  AND3_X1   g416(.A1(new_n615_), .A2(new_n616_), .A3(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n617_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT31), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n620_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT83), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n412_), .A2(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n372_), .A2(KEYINPUT83), .A3(new_n375_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n623_), .A2(KEYINPUT31), .A3(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n621_), .A2(new_n625_), .A3(KEYINPUT82), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NOR3_X1   g426(.A1(new_n618_), .A2(new_n619_), .A3(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n617_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n616_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n495_), .B1(new_n515_), .B2(new_n517_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(KEYINPUT80), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n632_), .A2(new_n525_), .A3(new_n518_), .ZN(new_n633_));
  AOI21_X1  g432(.A(KEYINPUT30), .B1(new_n633_), .B2(new_n510_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n629_), .B1(new_n630_), .B2(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n615_), .A2(new_n616_), .A3(new_n617_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n626_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n613_), .B1(new_n628_), .B2(new_n637_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n627_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n635_), .A2(new_n636_), .A3(new_n626_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n639_), .A2(new_n612_), .A3(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n638_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n642_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n481_), .A2(new_n644_), .A3(new_n486_), .A4(new_n582_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT98), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n645_), .A2(new_n646_), .ZN(new_n648_));
  OAI22_X1  g447(.A1(new_n607_), .A2(new_n643_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n246_), .A2(new_n353_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT76), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n650_), .B(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(G229gat), .A2(G233gat), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n238_), .B(KEYINPUT75), .Z(new_n655_));
  AOI21_X1  g454(.A(new_n654_), .B1(new_n655_), .B2(new_n343_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n655_), .B(new_n343_), .ZN(new_n657_));
  AOI22_X1  g456(.A1(new_n652_), .A2(new_n656_), .B1(new_n657_), .B2(new_n654_), .ZN(new_n658_));
  XOR2_X1   g457(.A(G113gat), .B(G141gat), .Z(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT77), .ZN(new_n660_));
  XNOR2_X1  g459(.A(G169gat), .B(G197gat), .ZN(new_n661_));
  XOR2_X1   g460(.A(new_n660_), .B(new_n661_), .Z(new_n662_));
  XNOR2_X1  g461(.A(new_n658_), .B(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n649_), .A2(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(KEYINPUT99), .B1(new_n362_), .B2(new_n664_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n360_), .B(KEYINPUT74), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT99), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n666_), .A2(new_n667_), .A3(new_n649_), .A4(new_n663_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n665_), .A2(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n669_), .A2(new_n338_), .A3(new_n428_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT38), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n585_), .A2(new_n606_), .ZN(new_n673_));
  OAI211_X1 g472(.A(new_n427_), .B(new_n582_), .C1(new_n583_), .C2(new_n584_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n585_), .A2(KEYINPUT98), .A3(new_n582_), .A4(new_n644_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n645_), .A2(new_n646_), .ZN(new_n677_));
  AOI22_X1  g476(.A1(new_n675_), .A2(new_n642_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT100), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n261_), .A2(new_n679_), .A3(new_n263_), .ZN(new_n680_));
  OAI21_X1  g479(.A(KEYINPUT100), .B1(new_n274_), .B2(new_n269_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n678_), .A2(new_n683_), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n320_), .A2(KEYINPUT13), .A3(new_n323_), .ZN(new_n685_));
  AOI21_X1  g484(.A(KEYINPUT13), .B1(new_n320_), .B2(new_n323_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n359_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n684_), .A2(new_n663_), .A3(new_n687_), .A4(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(G1gat), .B1(new_n689_), .B2(new_n427_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n670_), .A2(new_n671_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n672_), .A2(new_n690_), .A3(new_n691_), .ZN(G1324gat));
  NOR2_X1   g491(.A1(new_n582_), .A2(G8gat), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n665_), .A2(new_n668_), .A3(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(KEYINPUT101), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT101), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n665_), .A2(new_n668_), .A3(new_n696_), .A4(new_n693_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(new_n698_));
  OAI21_X1  g497(.A(G8gat), .B1(new_n689_), .B2(new_n582_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT39), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n698_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT40), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n698_), .A2(KEYINPUT40), .A3(new_n700_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(G1325gat));
  OAI21_X1  g504(.A(G15gat), .B1(new_n689_), .B2(new_n642_), .ZN(new_n706_));
  XOR2_X1   g505(.A(new_n706_), .B(KEYINPUT41), .Z(new_n707_));
  NAND3_X1  g506(.A1(new_n669_), .A2(new_n609_), .A3(new_n643_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(KEYINPUT102), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT102), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n707_), .A2(new_n711_), .A3(new_n708_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(G1326gat));
  OAI21_X1  g512(.A(G22gat), .B1(new_n689_), .B2(new_n585_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT42), .ZN(new_n715_));
  INV_X1    g514(.A(G22gat), .ZN(new_n716_));
  INV_X1    g515(.A(new_n585_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n669_), .A2(new_n716_), .A3(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n715_), .A2(new_n718_), .ZN(G1327gat));
  NAND3_X1  g518(.A1(new_n359_), .A2(new_n681_), .A3(new_n680_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n328_), .A2(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n645_), .B(KEYINPUT98), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n643_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n723_));
  OAI211_X1 g522(.A(new_n663_), .B(new_n721_), .C1(new_n722_), .C2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT106), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n649_), .A2(KEYINPUT106), .A3(new_n663_), .A4(new_n721_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  OR3_X1    g527(.A1(new_n728_), .A2(G29gat), .A3(new_n427_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n662_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n658_), .B(new_n730_), .ZN(new_n731_));
  NOR3_X1   g530(.A1(new_n328_), .A2(new_n731_), .A3(new_n688_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n265_), .B1(new_n256_), .B2(new_n260_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n271_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n264_), .B1(new_n735_), .B2(new_n263_), .ZN(new_n736_));
  OAI21_X1  g535(.A(KEYINPUT71), .B1(new_n734_), .B2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(new_n275_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT103), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n649_), .B2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n678_), .A2(KEYINPUT103), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n733_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n649_), .A2(KEYINPUT104), .A3(new_n733_), .A4(new_n277_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT104), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n277_), .A2(new_n733_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n744_), .B1(new_n678_), .B2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n743_), .A2(new_n746_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n732_), .B1(new_n742_), .B2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT44), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  OAI211_X1 g549(.A(KEYINPUT44), .B(new_n732_), .C1(new_n742_), .C2(new_n747_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n750_), .A2(new_n428_), .A3(new_n751_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n752_), .A2(KEYINPUT105), .ZN(new_n753_));
  OAI21_X1  g552(.A(G29gat), .B1(new_n752_), .B2(KEYINPUT105), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n729_), .B1(new_n753_), .B2(new_n754_), .ZN(G1328gat));
  INV_X1    g554(.A(KEYINPUT46), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n756_), .A2(KEYINPUT107), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n582_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n750_), .A2(new_n759_), .A3(new_n751_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(G36gat), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n582_), .A2(G36gat), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n726_), .A2(new_n727_), .A3(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT45), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT45), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n726_), .A2(new_n765_), .A3(new_n727_), .A4(new_n762_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n756_), .A2(KEYINPUT107), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n758_), .B1(new_n761_), .B2(new_n770_), .ZN(new_n771_));
  AOI211_X1 g570(.A(new_n757_), .B(new_n769_), .C1(new_n760_), .C2(G36gat), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n771_), .A2(new_n772_), .ZN(G1329gat));
  NAND4_X1  g572(.A1(new_n750_), .A2(G43gat), .A3(new_n643_), .A4(new_n751_), .ZN(new_n774_));
  INV_X1    g573(.A(G43gat), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n775_), .B1(new_n728_), .B2(new_n642_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g577(.A(new_n728_), .ZN(new_n779_));
  AOI21_X1  g578(.A(G50gat), .B1(new_n779_), .B2(new_n717_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n750_), .A2(new_n751_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n717_), .A2(G50gat), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n780_), .B1(new_n781_), .B2(new_n782_), .ZN(G1331gat));
  OAI21_X1  g582(.A(new_n731_), .B1(new_n351_), .B2(new_n358_), .ZN(new_n784_));
  NOR4_X1   g583(.A1(new_n678_), .A2(new_n687_), .A3(new_n683_), .A4(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n428_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n328_), .A2(new_n738_), .A3(new_n688_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT108), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n787_), .A2(new_n788_), .ZN(new_n790_));
  NOR4_X1   g589(.A1(new_n789_), .A2(new_n790_), .A3(new_n678_), .A4(new_n663_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n427_), .A2(G57gat), .ZN(new_n792_));
  AOI22_X1  g591(.A1(G57gat), .A2(new_n786_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT109), .ZN(G1332gat));
  INV_X1    g593(.A(G64gat), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n795_), .B1(new_n785_), .B2(new_n759_), .ZN(new_n796_));
  XOR2_X1   g595(.A(new_n796_), .B(KEYINPUT48), .Z(new_n797_));
  NAND3_X1  g596(.A1(new_n791_), .A2(new_n795_), .A3(new_n759_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(G1333gat));
  INV_X1    g598(.A(G71gat), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n800_), .B1(new_n785_), .B2(new_n643_), .ZN(new_n801_));
  XOR2_X1   g600(.A(new_n801_), .B(KEYINPUT49), .Z(new_n802_));
  NAND3_X1  g601(.A1(new_n791_), .A2(new_n800_), .A3(new_n643_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(G1334gat));
  AOI21_X1  g603(.A(new_n470_), .B1(new_n785_), .B2(new_n717_), .ZN(new_n805_));
  XOR2_X1   g604(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n806_));
  XNOR2_X1  g605(.A(new_n805_), .B(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n791_), .A2(new_n470_), .A3(new_n717_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(G1335gat));
  NOR4_X1   g608(.A1(new_n678_), .A2(new_n663_), .A3(new_n687_), .A4(new_n720_), .ZN(new_n810_));
  INV_X1    g609(.A(G85gat), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n810_), .A2(new_n811_), .A3(new_n428_), .ZN(new_n812_));
  NOR3_X1   g611(.A1(new_n687_), .A2(new_n663_), .A3(new_n688_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n813_), .B1(new_n742_), .B2(new_n747_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT111), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT111), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n816_), .B(new_n813_), .C1(new_n742_), .C2(new_n747_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n427_), .B1(new_n815_), .B2(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n812_), .B1(new_n818_), .B2(new_n811_), .ZN(G1336gat));
  AOI21_X1  g618(.A(G92gat), .B1(new_n810_), .B2(new_n759_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n815_), .A2(new_n817_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n759_), .A2(G92gat), .ZN(new_n822_));
  XOR2_X1   g621(.A(new_n822_), .B(KEYINPUT112), .Z(new_n823_));
  AOI21_X1  g622(.A(new_n820_), .B1(new_n821_), .B2(new_n823_), .ZN(G1337gat));
  NAND3_X1  g623(.A1(new_n810_), .A2(new_n643_), .A3(new_n204_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n642_), .B1(new_n815_), .B2(new_n817_), .ZN(new_n826_));
  INV_X1    g625(.A(G99gat), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n825_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT113), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT51), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n828_), .A2(new_n831_), .ZN(new_n832_));
  OAI221_X1 g631(.A(new_n825_), .B1(new_n829_), .B2(new_n830_), .C1(new_n826_), .C2(new_n827_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(G1338gat));
  NAND3_X1  g633(.A1(new_n810_), .A2(new_n205_), .A3(new_n717_), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n717_), .B(new_n813_), .C1(new_n742_), .C2(new_n747_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(KEYINPUT114), .B(KEYINPUT52), .ZN(new_n837_));
  AND3_X1   g636(.A1(new_n836_), .A2(G106gat), .A3(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n837_), .B1(new_n836_), .B2(G106gat), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n835_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(KEYINPUT53), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n842_), .B(new_n835_), .C1(new_n838_), .C2(new_n839_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n843_), .ZN(G1339gat));
  NAND2_X1  g643(.A1(new_n658_), .A2(new_n662_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n662_), .B1(new_n657_), .B2(new_n653_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n653_), .B1(new_n655_), .B2(new_n343_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n652_), .A2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n324_), .A2(new_n845_), .A3(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n315_), .A2(KEYINPUT55), .A3(new_n316_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n280_), .B1(new_n298_), .B2(new_n288_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT55), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n853_), .B1(new_n298_), .B2(new_n300_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n851_), .A2(new_n852_), .A3(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n322_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT118), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n856_), .A2(new_n857_), .A3(KEYINPUT56), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n731_), .B1(new_n302_), .B2(new_n319_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(KEYINPUT56), .B1(new_n856_), .B2(new_n857_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n850_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n682_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT58), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n856_), .A2(KEYINPUT56), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n845_), .A2(new_n849_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT56), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n855_), .A2(new_n868_), .A3(new_n322_), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n866_), .A2(new_n320_), .A3(new_n867_), .A4(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n738_), .B1(new_n865_), .B2(new_n870_), .ZN(new_n871_));
  OR2_X1    g670(.A1(new_n870_), .A2(new_n865_), .ZN(new_n872_));
  AOI22_X1  g671(.A1(new_n863_), .A2(new_n864_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n862_), .A2(KEYINPUT57), .A3(new_n682_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n688_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT117), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT54), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n685_), .A2(new_n784_), .A3(new_n686_), .ZN(new_n879_));
  AOI211_X1 g678(.A(KEYINPUT116), .B(new_n878_), .C1(new_n879_), .C2(new_n738_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT116), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n350_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n882_));
  OAI22_X1  g681(.A1(new_n357_), .A2(new_n882_), .B1(new_n356_), .B2(new_n332_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n349_), .A2(KEYINPUT17), .A3(new_n350_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n663_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n687_), .A2(new_n738_), .A3(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n881_), .B1(new_n886_), .B2(KEYINPUT54), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n880_), .A2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT115), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n878_), .B1(new_n273_), .B2(new_n276_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n326_), .A2(new_n327_), .A3(new_n885_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n889_), .B1(new_n890_), .B2(new_n891_), .ZN(new_n892_));
  AOI21_X1  g691(.A(KEYINPUT54), .B1(new_n737_), .B2(new_n275_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n879_), .A2(KEYINPUT115), .A3(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n894_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n877_), .B1(new_n888_), .B2(new_n895_), .ZN(new_n896_));
  OAI21_X1  g695(.A(KEYINPUT54), .B1(new_n277_), .B2(new_n891_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(KEYINPUT116), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n886_), .A2(new_n881_), .A3(KEYINPUT54), .ZN(new_n899_));
  NAND4_X1  g698(.A1(new_n895_), .A2(new_n898_), .A3(new_n877_), .A4(new_n899_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n876_), .B1(new_n896_), .B2(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n717_), .A2(new_n759_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n903_), .A2(new_n428_), .A3(new_n643_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n902_), .A2(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n906_), .ZN(new_n907_));
  AOI21_X1  g706(.A(G113gat), .B1(new_n907_), .B2(new_n663_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n909_), .B1(new_n902_), .B2(new_n905_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n895_), .A2(new_n898_), .A3(new_n899_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(KEYINPUT117), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n875_), .B1(new_n912_), .B2(new_n900_), .ZN(new_n913_));
  XOR2_X1   g712(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n914_));
  NOR3_X1   g713(.A1(new_n913_), .A2(new_n904_), .A3(new_n914_), .ZN(new_n915_));
  OAI21_X1  g714(.A(KEYINPUT120), .B1(new_n910_), .B2(new_n915_), .ZN(new_n916_));
  OAI22_X1  g715(.A1(new_n913_), .A2(new_n904_), .B1(KEYINPUT119), .B2(KEYINPUT59), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT120), .ZN(new_n918_));
  OAI211_X1 g717(.A(new_n917_), .B(new_n918_), .C1(new_n906_), .C2(new_n914_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n916_), .A2(new_n919_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT121), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n921_), .A2(G113gat), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n663_), .A2(KEYINPUT121), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n922_), .B1(new_n923_), .B2(G113gat), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n908_), .B1(new_n920_), .B2(new_n924_), .ZN(G1340gat));
  INV_X1    g724(.A(G120gat), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n926_), .B1(new_n687_), .B2(KEYINPUT60), .ZN(new_n927_));
  OAI211_X1 g726(.A(new_n907_), .B(new_n927_), .C1(KEYINPUT60), .C2(new_n926_), .ZN(new_n928_));
  NOR3_X1   g727(.A1(new_n910_), .A2(new_n915_), .A3(new_n687_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n929_), .B2(new_n926_), .ZN(G1341gat));
  AOI21_X1  g729(.A(G127gat), .B1(new_n907_), .B2(new_n688_), .ZN(new_n931_));
  AND2_X1   g730(.A1(new_n688_), .A2(G127gat), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n931_), .B1(new_n920_), .B2(new_n932_), .ZN(G1342gat));
  AOI21_X1  g732(.A(G134gat), .B1(new_n907_), .B2(new_n683_), .ZN(new_n934_));
  AND2_X1   g733(.A1(new_n277_), .A2(G134gat), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n934_), .B1(new_n920_), .B2(new_n935_), .ZN(G1343gat));
  NOR3_X1   g735(.A1(new_n759_), .A2(new_n427_), .A3(new_n643_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n717_), .A2(new_n937_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n913_), .A2(new_n938_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n939_), .A2(new_n663_), .ZN(new_n940_));
  XNOR2_X1  g739(.A(KEYINPUT122), .B(G141gat), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n940_), .B(new_n941_), .ZN(G1344gat));
  NAND2_X1  g741(.A1(new_n939_), .A2(new_n328_), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n943_), .B(G148gat), .ZN(G1345gat));
  NAND4_X1  g743(.A1(new_n902_), .A2(new_n717_), .A3(new_n688_), .A4(new_n937_), .ZN(new_n945_));
  INV_X1    g744(.A(KEYINPUT123), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n945_), .A2(new_n946_), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n939_), .A2(KEYINPUT123), .A3(new_n688_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(KEYINPUT61), .B(G155gat), .ZN(new_n949_));
  AND3_X1   g748(.A1(new_n947_), .A2(new_n948_), .A3(new_n949_), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n949_), .B1(new_n947_), .B2(new_n948_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n950_), .A2(new_n951_), .ZN(G1346gat));
  NAND3_X1  g751(.A1(new_n939_), .A2(new_n380_), .A3(new_n683_), .ZN(new_n953_));
  NOR3_X1   g752(.A1(new_n913_), .A2(new_n738_), .A3(new_n938_), .ZN(new_n954_));
  OAI21_X1  g753(.A(new_n953_), .B1(new_n954_), .B2(new_n380_), .ZN(G1347gat));
  NAND3_X1  g754(.A1(new_n585_), .A2(new_n759_), .A3(new_n644_), .ZN(new_n956_));
  NOR3_X1   g755(.A1(new_n913_), .A2(new_n731_), .A3(new_n956_), .ZN(new_n957_));
  NOR2_X1   g756(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n958_));
  INV_X1    g757(.A(KEYINPUT124), .ZN(new_n959_));
  INV_X1    g758(.A(KEYINPUT62), .ZN(new_n960_));
  OAI21_X1  g759(.A(G169gat), .B1(new_n959_), .B2(new_n960_), .ZN(new_n961_));
  OR3_X1    g760(.A1(new_n957_), .A2(new_n958_), .A3(new_n961_), .ZN(new_n962_));
  OAI21_X1  g761(.A(new_n958_), .B1(new_n957_), .B2(new_n961_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n957_), .A2(new_n527_), .ZN(new_n964_));
  NAND3_X1  g763(.A1(new_n962_), .A2(new_n963_), .A3(new_n964_), .ZN(G1348gat));
  NOR2_X1   g764(.A1(new_n913_), .A2(new_n956_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n966_), .A2(new_n328_), .ZN(new_n967_));
  XNOR2_X1  g766(.A(new_n967_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g767(.A1(new_n966_), .A2(new_n688_), .ZN(new_n969_));
  NOR2_X1   g768(.A1(new_n969_), .A2(new_n499_), .ZN(new_n970_));
  AOI21_X1  g769(.A(new_n970_), .B1(new_n521_), .B2(new_n969_), .ZN(G1350gat));
  NAND4_X1  g770(.A1(new_n966_), .A2(new_n542_), .A3(new_n538_), .A4(new_n683_), .ZN(new_n972_));
  NOR3_X1   g771(.A1(new_n913_), .A2(new_n738_), .A3(new_n956_), .ZN(new_n973_));
  OAI21_X1  g772(.A(new_n972_), .B1(new_n973_), .B2(new_n522_), .ZN(G1351gat));
  NAND3_X1  g773(.A1(new_n487_), .A2(new_n759_), .A3(new_n642_), .ZN(new_n975_));
  NOR2_X1   g774(.A1(new_n913_), .A2(new_n975_), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n976_), .A2(new_n663_), .ZN(new_n977_));
  XNOR2_X1  g776(.A(new_n977_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g777(.A1(new_n976_), .A2(new_n328_), .ZN(new_n979_));
  INV_X1    g778(.A(KEYINPUT125), .ZN(new_n980_));
  OAI21_X1  g779(.A(new_n979_), .B1(new_n980_), .B2(G204gat), .ZN(new_n981_));
  XNOR2_X1  g780(.A(KEYINPUT125), .B(G204gat), .ZN(new_n982_));
  OAI21_X1  g781(.A(new_n981_), .B1(new_n979_), .B2(new_n982_), .ZN(G1353gat));
  AOI21_X1  g782(.A(new_n359_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n984_));
  NAND2_X1  g783(.A1(new_n976_), .A2(new_n984_), .ZN(new_n985_));
  INV_X1    g784(.A(KEYINPUT127), .ZN(new_n986_));
  NOR2_X1   g785(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n987_));
  XNOR2_X1  g786(.A(new_n987_), .B(KEYINPUT126), .ZN(new_n988_));
  AOI21_X1  g787(.A(new_n985_), .B1(new_n986_), .B2(new_n988_), .ZN(new_n989_));
  XNOR2_X1  g788(.A(new_n988_), .B(new_n986_), .ZN(new_n990_));
  AOI21_X1  g789(.A(new_n989_), .B1(new_n985_), .B2(new_n990_), .ZN(G1354gat));
  INV_X1    g790(.A(G218gat), .ZN(new_n992_));
  NAND3_X1  g791(.A1(new_n976_), .A2(new_n992_), .A3(new_n683_), .ZN(new_n993_));
  NOR3_X1   g792(.A1(new_n913_), .A2(new_n738_), .A3(new_n975_), .ZN(new_n994_));
  OAI21_X1  g793(.A(new_n993_), .B1(new_n994_), .B2(new_n992_), .ZN(G1355gat));
endmodule


