//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 0 0 1 1 0 1 1 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 1 0 1 1 1 0 1 0 1 1 0 1 1 1 0 0 0 1 0 0 1 0 0 0 1 0 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n764_, new_n765_, new_n766_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n882_, new_n883_,
    new_n885_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n908_, new_n909_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n923_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_;
  INV_X1    g000(.A(KEYINPUT105), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT27), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G226gat), .A2(G233gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT19), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT96), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT23), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT23), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n209_), .A2(G183gat), .A3(G190gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  OR3_X1    g010(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT79), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT78), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT78), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(G169gat), .A3(G176gat), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(G169gat), .ZN(new_n221_));
  INV_X1    g020(.A(G176gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT24), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n220_), .A2(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n211_), .A2(KEYINPUT79), .A3(new_n212_), .ZN(new_n227_));
  INV_X1    g026(.A(G190gat), .ZN(new_n228_));
  OR2_X1    g027(.A1(new_n228_), .A2(KEYINPUT26), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT25), .B(G183gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n228_), .A2(KEYINPUT77), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT77), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(G190gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n231_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT26), .ZN(new_n235_));
  OAI211_X1 g034(.A(new_n229_), .B(new_n230_), .C1(new_n234_), .C2(new_n235_), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n215_), .A2(new_n226_), .A3(new_n227_), .A4(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT80), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n208_), .A2(new_n210_), .A3(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n207_), .A2(KEYINPUT80), .A3(KEYINPUT23), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n239_), .B(new_n240_), .C1(new_n234_), .C2(G183gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT22), .B(G169gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(new_n222_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n241_), .A2(new_n243_), .A3(new_n220_), .ZN(new_n244_));
  AND3_X1   g043(.A1(new_n237_), .A2(KEYINPUT81), .A3(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(G204gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT91), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT91), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(G204gat), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n247_), .A2(new_n249_), .A3(G197gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT93), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT93), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n247_), .A2(new_n249_), .A3(new_n252_), .A4(G197gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT90), .B(G197gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(G204gat), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n251_), .A2(new_n253_), .A3(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G211gat), .B(G218gat), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n256_), .A2(KEYINPUT21), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT21), .ZN(new_n260_));
  INV_X1    g059(.A(G197gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT90), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT90), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(G197gat), .ZN(new_n264_));
  AOI21_X1  g063(.A(G204gat), .B1(new_n262_), .B2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n247_), .A2(new_n249_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(new_n261_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n265_), .B1(new_n267_), .B2(KEYINPUT92), .ZN(new_n268_));
  AOI21_X1  g067(.A(G197gat), .B1(new_n247_), .B2(new_n249_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT92), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n260_), .B1(new_n268_), .B2(new_n271_), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n251_), .A2(new_n260_), .A3(new_n253_), .A4(new_n255_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(new_n257_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n259_), .B1(new_n272_), .B2(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(KEYINPUT81), .B1(new_n237_), .B2(new_n244_), .ZN(new_n276_));
  NOR3_X1   g075(.A1(new_n245_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n258_), .A2(KEYINPUT21), .ZN(new_n278_));
  AOI22_X1  g077(.A1(new_n250_), .A2(KEYINPUT93), .B1(new_n254_), .B2(G204gat), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n278_), .B1(new_n279_), .B2(new_n253_), .ZN(new_n280_));
  AND2_X1   g079(.A1(new_n273_), .A2(new_n257_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n271_), .ZN(new_n282_));
  OAI22_X1  g081(.A1(new_n269_), .A2(new_n270_), .B1(G204gat), .B2(new_n254_), .ZN(new_n283_));
  OAI21_X1  g082(.A(KEYINPUT21), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n280_), .B1(new_n281_), .B2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n239_), .A2(new_n240_), .A3(new_n212_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT97), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n239_), .A2(KEYINPUT97), .A3(new_n240_), .A4(new_n212_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n230_), .A2(new_n229_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n228_), .A2(KEYINPUT26), .ZN(new_n292_));
  AOI22_X1  g091(.A1(new_n291_), .A2(new_n292_), .B1(new_n216_), .B2(new_n225_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(G183gat), .A2(G190gat), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n294_), .B1(new_n208_), .B2(new_n210_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT99), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT98), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n221_), .A2(KEYINPUT22), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT22), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(G169gat), .ZN(new_n300_));
  AND3_X1   g099(.A1(new_n298_), .A2(new_n300_), .A3(new_n222_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n217_), .A2(new_n219_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n297_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n243_), .A2(new_n220_), .A3(KEYINPUT98), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  AOI22_X1  g104(.A1(new_n290_), .A2(new_n293_), .B1(new_n296_), .B2(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(KEYINPUT20), .B1(new_n285_), .B2(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n206_), .B1(new_n277_), .B2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT20), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n309_), .B1(new_n285_), .B2(new_n306_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n205_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n275_), .B1(new_n245_), .B2(new_n276_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n310_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n313_));
  XOR2_X1   g112(.A(G8gat), .B(G36gat), .Z(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT18), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G64gat), .B(G92gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n308_), .A2(new_n313_), .A3(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT100), .ZN(new_n319_));
  AND2_X1   g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n317_), .ZN(new_n321_));
  AND3_X1   g120(.A1(new_n310_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n206_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n290_), .A2(new_n293_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n296_), .A2(new_n305_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n309_), .B1(new_n326_), .B2(new_n275_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n237_), .A2(new_n244_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT81), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n237_), .A2(KEYINPUT81), .A3(new_n244_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n285_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n323_), .B1(new_n327_), .B2(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n321_), .B1(new_n322_), .B2(new_n333_), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n308_), .A2(KEYINPUT100), .A3(new_n313_), .A4(new_n317_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n203_), .B1(new_n320_), .B2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT104), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n318_), .A2(new_n319_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n340_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n341_), .A2(KEYINPUT104), .A3(new_n203_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n339_), .A2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G1gat), .B(G29gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(G85gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT0), .B(G57gat), .ZN(new_n346_));
  XOR2_X1   g145(.A(new_n345_), .B(new_n346_), .Z(new_n347_));
  INV_X1    g146(.A(G155gat), .ZN(new_n348_));
  INV_X1    g147(.A(G162gat), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(G155gat), .A2(G162gat), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT2), .ZN(new_n353_));
  AND3_X1   g152(.A1(KEYINPUT84), .A2(G141gat), .A3(G148gat), .ZN(new_n354_));
  AOI21_X1  g153(.A(KEYINPUT84), .B1(G141gat), .B2(G148gat), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n353_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT87), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n357_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n358_));
  NAND3_X1  g157(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(KEYINPUT87), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n356_), .A2(new_n358_), .A3(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT86), .ZN(new_n362_));
  NOR2_X1   g161(.A1(G141gat), .A2(G148gat), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n362_), .B1(new_n363_), .B2(KEYINPUT85), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT3), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT85), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n366_), .B1(new_n365_), .B2(KEYINPUT86), .ZN(new_n367_));
  AOI22_X1  g166(.A1(new_n364_), .A2(new_n365_), .B1(new_n363_), .B2(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n352_), .B1(new_n361_), .B2(new_n368_), .ZN(new_n369_));
  XOR2_X1   g168(.A(G127gat), .B(G134gat), .Z(new_n370_));
  XOR2_X1   g169(.A(G113gat), .B(G120gat), .Z(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT1), .B1(new_n348_), .B2(new_n349_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n351_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT1), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n375_), .A2(G155gat), .A3(G162gat), .ZN(new_n376_));
  AND3_X1   g175(.A1(new_n373_), .A2(new_n374_), .A3(new_n376_), .ZN(new_n377_));
  OR2_X1    g176(.A1(G141gat), .A2(G148gat), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n378_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n379_));
  OR2_X1    g178(.A1(new_n377_), .A2(new_n379_), .ZN(new_n380_));
  AND3_X1   g179(.A1(new_n369_), .A2(new_n372_), .A3(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n372_), .B1(new_n369_), .B2(new_n380_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT4), .ZN(new_n383_));
  NOR3_X1   g182(.A1(new_n381_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n369_), .A2(new_n380_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n372_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(new_n383_), .A3(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G225gat), .A2(G233gat), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n387_), .A2(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT101), .B1(new_n384_), .B2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n352_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n360_), .A2(new_n358_), .ZN(new_n393_));
  OR2_X1    g192(.A1(new_n354_), .A2(new_n355_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n393_), .B1(new_n394_), .B2(new_n353_), .ZN(new_n395_));
  AOI21_X1  g194(.A(KEYINPUT86), .B1(new_n378_), .B2(new_n366_), .ZN(new_n396_));
  AOI21_X1  g195(.A(KEYINPUT85), .B1(new_n362_), .B2(KEYINPUT3), .ZN(new_n397_));
  OAI22_X1  g196(.A1(new_n396_), .A2(KEYINPUT3), .B1(new_n378_), .B2(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n392_), .B1(new_n395_), .B2(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n377_), .A2(new_n379_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n386_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n369_), .A2(new_n372_), .A3(new_n380_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n401_), .A2(KEYINPUT4), .A3(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n388_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT101), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n403_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n406_));
  NOR3_X1   g205(.A1(new_n381_), .A2(new_n382_), .A3(new_n389_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  AND4_X1   g207(.A1(new_n347_), .A2(new_n391_), .A3(new_n406_), .A4(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n403_), .A2(new_n404_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n407_), .B1(new_n410_), .B2(KEYINPUT101), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n347_), .B1(new_n411_), .B2(new_n406_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n409_), .A2(new_n412_), .ZN(new_n413_));
  AND3_X1   g212(.A1(new_n327_), .A2(new_n332_), .A3(new_n323_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n311_), .B1(new_n310_), .B2(new_n312_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n321_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n416_), .A2(KEYINPUT27), .A3(new_n318_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n413_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT95), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G228gat), .A2(G233gat), .ZN(new_n420_));
  XOR2_X1   g219(.A(new_n420_), .B(KEYINPUT89), .Z(new_n421_));
  NAND2_X1  g220(.A1(new_n385_), .A2(KEYINPUT29), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n421_), .B1(new_n275_), .B2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n393_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n397_), .A2(new_n378_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n366_), .B1(G141gat), .B2(G148gat), .ZN(new_n426_));
  AOI21_X1  g225(.A(KEYINPUT3), .B1(new_n426_), .B2(new_n362_), .ZN(new_n427_));
  OAI211_X1 g226(.A(new_n424_), .B(new_n356_), .C1(new_n425_), .C2(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n400_), .B1(new_n428_), .B2(new_n352_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT29), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT88), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT88), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n385_), .A2(new_n432_), .A3(KEYINPUT29), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n431_), .A2(new_n433_), .A3(new_n275_), .A4(new_n421_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT94), .ZN(new_n435_));
  INV_X1    g234(.A(new_n421_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n281_), .A2(new_n284_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n436_), .B1(new_n437_), .B2(new_n259_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT94), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n438_), .A2(new_n439_), .A3(new_n431_), .A4(new_n433_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n423_), .B1(new_n435_), .B2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G78gat), .B(G106gat), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n419_), .B1(new_n441_), .B2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n429_), .A2(new_n430_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G22gat), .B(G50gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(KEYINPUT28), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n445_), .B(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n441_), .A2(new_n443_), .ZN(new_n450_));
  AOI211_X1 g249(.A(new_n423_), .B(new_n442_), .C1(new_n435_), .C2(new_n440_), .ZN(new_n451_));
  OAI22_X1  g250(.A1(new_n444_), .A2(new_n449_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  AND2_X1   g251(.A1(new_n435_), .A2(new_n440_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n442_), .B1(new_n453_), .B2(new_n423_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n441_), .A2(new_n443_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n454_), .A2(new_n419_), .A3(new_n455_), .A4(new_n448_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n418_), .B1(new_n452_), .B2(new_n456_), .ZN(new_n457_));
  AND2_X1   g256(.A1(new_n452_), .A2(new_n456_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n317_), .A2(KEYINPUT32), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(KEYINPUT102), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n460_), .A2(new_n308_), .A3(new_n313_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT103), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n414_), .A2(new_n415_), .ZN(new_n464_));
  OAI22_X1  g263(.A1(new_n409_), .A2(new_n412_), .B1(new_n464_), .B2(new_n459_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n411_), .A2(new_n347_), .A3(new_n406_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT33), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n411_), .A2(KEYINPUT33), .A3(new_n347_), .A4(new_n406_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n403_), .A2(new_n388_), .A3(new_n387_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n347_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n401_), .A2(new_n402_), .A3(new_n389_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n470_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n468_), .A2(new_n469_), .A3(new_n473_), .ZN(new_n474_));
  OAI22_X1  g273(.A1(new_n463_), .A2(new_n465_), .B1(new_n474_), .B2(new_n341_), .ZN(new_n475_));
  AOI22_X1  g274(.A1(new_n343_), .A2(new_n457_), .B1(new_n458_), .B2(new_n475_), .ZN(new_n476_));
  XOR2_X1   g275(.A(KEYINPUT83), .B(G15gat), .Z(new_n477_));
  NAND2_X1  g276(.A1(G227gat), .A2(G233gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(KEYINPUT82), .B(G43gat), .ZN(new_n480_));
  XOR2_X1   g279(.A(new_n479_), .B(new_n480_), .Z(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(new_n386_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n245_), .A2(new_n276_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(KEYINPUT30), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G71gat), .B(G99gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n485_), .A2(new_n486_), .ZN(new_n489_));
  NOR3_X1   g288(.A1(new_n488_), .A2(new_n489_), .A3(KEYINPUT31), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT31), .ZN(new_n491_));
  OR2_X1    g290(.A1(new_n485_), .A2(new_n486_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n491_), .B1(new_n492_), .B2(new_n487_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n483_), .B1(new_n490_), .B2(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(KEYINPUT31), .B1(new_n488_), .B2(new_n489_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n492_), .A2(new_n491_), .A3(new_n487_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n495_), .A2(new_n496_), .A3(new_n482_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n494_), .A2(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n202_), .B1(new_n476_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n342_), .ZN(new_n500_));
  AOI21_X1  g299(.A(KEYINPUT104), .B1(new_n341_), .B2(new_n203_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n457_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n475_), .A2(new_n458_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n498_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n504_), .A2(KEYINPUT105), .A3(new_n505_), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n343_), .A2(new_n417_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n413_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n508_), .B1(new_n494_), .B2(new_n497_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n507_), .A2(new_n458_), .A3(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n499_), .A2(new_n506_), .A3(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G15gat), .B(G22gat), .ZN(new_n513_));
  INV_X1    g312(.A(G1gat), .ZN(new_n514_));
  INV_X1    g313(.A(G8gat), .ZN(new_n515_));
  OAI21_X1  g314(.A(KEYINPUT14), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n513_), .A2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G1gat), .B(G8gat), .ZN(new_n518_));
  XOR2_X1   g317(.A(new_n517_), .B(new_n518_), .Z(new_n519_));
  XNOR2_X1  g318(.A(G29gat), .B(G36gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G43gat), .B(G50gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n519_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT75), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n519_), .A2(new_n522_), .ZN(new_n525_));
  XOR2_X1   g324(.A(new_n524_), .B(new_n525_), .Z(new_n526_));
  NAND2_X1  g325(.A1(G229gat), .A2(G233gat), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n522_), .B(KEYINPUT15), .ZN(new_n529_));
  INV_X1    g328(.A(new_n519_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT76), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n528_), .B1(new_n519_), .B2(new_n522_), .ZN(new_n533_));
  AOI22_X1  g332(.A1(new_n526_), .A2(new_n528_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G113gat), .B(G141gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G169gat), .B(G197gat), .ZN(new_n536_));
  XOR2_X1   g335(.A(new_n535_), .B(new_n536_), .Z(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n534_), .B(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n512_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G127gat), .B(G155gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT16), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G183gat), .B(G211gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(KEYINPUT74), .B1(new_n544_), .B2(KEYINPUT17), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(new_n530_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G231gat), .A2(G233gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(G57gat), .B(G64gat), .Z(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT66), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(KEYINPUT11), .ZN(new_n551_));
  XOR2_X1   g350(.A(G71gat), .B(G78gat), .Z(new_n552_));
  NOR2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n551_), .A2(new_n552_), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n550_), .A2(KEYINPUT11), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n553_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  OR2_X1    g355(.A1(new_n548_), .A2(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n544_), .A2(KEYINPUT17), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n558_), .B1(new_n548_), .B2(new_n556_), .ZN(new_n559_));
  AND2_X1   g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  XOR2_X1   g360(.A(G120gat), .B(G148gat), .Z(new_n562_));
  XNOR2_X1  g361(.A(G176gat), .B(G204gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  XOR2_X1   g365(.A(G85gat), .B(G92gat), .Z(new_n567_));
  NAND2_X1  g366(.A1(G99gat), .A2(G106gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT6), .ZN(new_n569_));
  OR2_X1    g368(.A1(G99gat), .A2(G106gat), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n569_), .B1(KEYINPUT7), .B2(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT65), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n567_), .B1(new_n571_), .B2(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT8), .ZN(new_n575_));
  XOR2_X1   g374(.A(KEYINPUT10), .B(G99gat), .Z(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT64), .B(G106gat), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n567_), .A2(KEYINPUT9), .ZN(new_n579_));
  INV_X1    g378(.A(G85gat), .ZN(new_n580_));
  INV_X1    g379(.A(G92gat), .ZN(new_n581_));
  OR3_X1    g380(.A1(new_n580_), .A2(new_n581_), .A3(KEYINPUT9), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n578_), .A2(new_n579_), .A3(new_n582_), .A4(new_n569_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n575_), .A2(new_n583_), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n584_), .A2(new_n556_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(KEYINPUT12), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(new_n556_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G230gat), .A2(G233gat), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n589_), .B1(new_n585_), .B2(new_n587_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n566_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT68), .ZN(new_n595_));
  NOR3_X1   g394(.A1(new_n591_), .A2(new_n592_), .A3(new_n566_), .ZN(new_n596_));
  NOR3_X1   g395(.A1(new_n594_), .A2(new_n595_), .A3(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n596_), .ZN(new_n598_));
  AOI21_X1  g397(.A(KEYINPUT68), .B1(new_n598_), .B2(new_n593_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT13), .ZN(new_n600_));
  OAI22_X1  g399(.A1(new_n597_), .A2(new_n599_), .B1(KEYINPUT69), .B2(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n595_), .B1(new_n594_), .B2(new_n596_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n598_), .A2(KEYINPUT68), .A3(new_n593_), .ZN(new_n603_));
  XOR2_X1   g402(.A(KEYINPUT69), .B(KEYINPUT13), .Z(new_n604_));
  NAND3_X1  g403(.A1(new_n602_), .A2(new_n603_), .A3(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n601_), .A2(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n575_), .A2(new_n522_), .A3(new_n583_), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n607_), .B(KEYINPUT71), .Z(new_n608_));
  XOR2_X1   g407(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n609_));
  NAND2_X1  g408(.A1(G232gat), .A2(G233gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(KEYINPUT35), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n612_), .A2(KEYINPUT72), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n611_), .A2(KEYINPUT35), .ZN(new_n614_));
  AOI211_X1 g413(.A(new_n613_), .B(new_n614_), .C1(new_n584_), .C2(new_n529_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n608_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n612_), .A2(KEYINPUT72), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n608_), .A2(new_n617_), .A3(new_n615_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G190gat), .B(G218gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G134gat), .B(G162gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n624_), .A2(KEYINPUT36), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n621_), .A2(new_n625_), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n624_), .B(KEYINPUT36), .Z(new_n627_));
  NAND3_X1  g426(.A1(new_n619_), .A2(new_n620_), .A3(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n626_), .A2(KEYINPUT37), .A3(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n627_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n631_), .B1(new_n621_), .B2(KEYINPUT73), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n632_), .B1(KEYINPUT73), .B2(new_n621_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(new_n626_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT37), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n630_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n540_), .A2(new_n561_), .A3(new_n606_), .A4(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n638_), .A2(new_n514_), .A3(new_n508_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT38), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n511_), .A2(new_n634_), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n641_), .B(KEYINPUT106), .Z(new_n642_));
  INV_X1    g441(.A(new_n606_), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n643_), .A2(new_n560_), .A3(new_n539_), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n642_), .A2(new_n644_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n645_), .A2(new_n508_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n640_), .B1(new_n514_), .B2(new_n646_), .ZN(G1324gat));
  INV_X1    g446(.A(new_n507_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n638_), .A2(new_n515_), .A3(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT39), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n645_), .A2(new_n648_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n650_), .B1(new_n651_), .B2(G8gat), .ZN(new_n652_));
  AOI211_X1 g451(.A(KEYINPUT39), .B(new_n515_), .C1(new_n645_), .C2(new_n648_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n649_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n654_), .B(new_n656_), .ZN(G1325gat));
  OR3_X1    g456(.A1(new_n637_), .A2(G15gat), .A3(new_n505_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n645_), .A2(new_n498_), .ZN(new_n659_));
  AND3_X1   g458(.A1(new_n659_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n660_));
  AOI21_X1  g459(.A(KEYINPUT41), .B1(new_n659_), .B2(G15gat), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n658_), .B1(new_n660_), .B2(new_n661_), .ZN(G1326gat));
  OR3_X1    g461(.A1(new_n637_), .A2(G22gat), .A3(new_n458_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n458_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n645_), .A2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(G22gat), .ZN(new_n666_));
  XOR2_X1   g465(.A(KEYINPUT108), .B(KEYINPUT42), .Z(new_n667_));
  AND2_X1   g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n666_), .A2(new_n667_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n663_), .B1(new_n668_), .B2(new_n669_), .ZN(G1327gat));
  NOR2_X1   g469(.A1(new_n634_), .A2(new_n561_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n606_), .A2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(new_n540_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(G29gat), .B1(new_n674_), .B2(new_n508_), .ZN(new_n675_));
  AOI211_X1 g474(.A(new_n561_), .B(new_n539_), .C1(new_n601_), .C2(new_n605_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n633_), .A2(new_n626_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n629_), .B1(new_n677_), .B2(KEYINPUT37), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT43), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n511_), .A2(new_n678_), .A3(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(KEYINPUT109), .B(KEYINPUT43), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n681_), .B1(new_n511_), .B2(new_n678_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT110), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n680_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  AOI211_X1 g483(.A(KEYINPUT110), .B(new_n681_), .C1(new_n511_), .C2(new_n678_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n676_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n688_), .A2(G29gat), .A3(new_n508_), .ZN(new_n689_));
  OAI211_X1 g488(.A(KEYINPUT44), .B(new_n676_), .C1(new_n684_), .C2(new_n685_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(KEYINPUT111), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n343_), .A2(new_n458_), .A3(new_n417_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n498_), .A2(new_n413_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n504_), .A2(new_n505_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n695_), .B2(new_n202_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n636_), .B1(new_n696_), .B2(new_n506_), .ZN(new_n697_));
  OAI21_X1  g496(.A(KEYINPUT110), .B1(new_n697_), .B2(new_n681_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n682_), .A2(new_n683_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n698_), .A2(new_n699_), .A3(new_n680_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT111), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n700_), .A2(new_n701_), .A3(KEYINPUT44), .A4(new_n676_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n691_), .A2(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n675_), .B1(new_n689_), .B2(new_n703_), .ZN(G1328gat));
  INV_X1    g503(.A(G36gat), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n674_), .A2(new_n705_), .A3(new_n648_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT45), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n507_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n703_), .A2(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(KEYINPUT112), .B1(new_n709_), .B2(G36gat), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT112), .ZN(new_n711_));
  AOI211_X1 g510(.A(new_n711_), .B(new_n705_), .C1(new_n703_), .C2(new_n708_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n707_), .B1(new_n710_), .B2(new_n712_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(KEYINPUT113), .A2(KEYINPUT46), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  OAI221_X1 g514(.A(new_n707_), .B1(KEYINPUT113), .B2(KEYINPUT46), .C1(new_n710_), .C2(new_n712_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1329gat));
  NAND4_X1  g516(.A1(new_n703_), .A2(G43gat), .A3(new_n498_), .A4(new_n688_), .ZN(new_n718_));
  INV_X1    g517(.A(G43gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n719_), .B1(new_n673_), .B2(new_n505_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT114), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n718_), .A2(new_n721_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(KEYINPUT115), .B(KEYINPUT47), .ZN(new_n723_));
  XOR2_X1   g522(.A(new_n722_), .B(new_n723_), .Z(G1330gat));
  AOI21_X1  g523(.A(G50gat), .B1(new_n674_), .B2(new_n664_), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n688_), .A2(G50gat), .A3(new_n664_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n726_), .B2(new_n703_), .ZN(G1331gat));
  INV_X1    g526(.A(G57gat), .ZN(new_n728_));
  INV_X1    g527(.A(new_n539_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n560_), .A2(new_n729_), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n642_), .A2(new_n643_), .A3(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n728_), .B1(new_n731_), .B2(new_n508_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n512_), .A2(new_n729_), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n733_), .A2(new_n561_), .A3(new_n643_), .A4(new_n636_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n734_), .A2(G57gat), .A3(new_n413_), .ZN(new_n735_));
  OR2_X1    g534(.A1(new_n732_), .A2(new_n735_), .ZN(G1332gat));
  OR3_X1    g535(.A1(new_n734_), .A2(G64gat), .A3(new_n507_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n731_), .A2(new_n648_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(G64gat), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n739_), .A2(KEYINPUT48), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n739_), .A2(KEYINPUT48), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n737_), .B1(new_n740_), .B2(new_n741_), .ZN(G1333gat));
  OR3_X1    g541(.A1(new_n734_), .A2(G71gat), .A3(new_n505_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n731_), .A2(new_n498_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(G71gat), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n745_), .A2(KEYINPUT49), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n745_), .A2(KEYINPUT49), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n743_), .B1(new_n746_), .B2(new_n747_), .ZN(G1334gat));
  OR3_X1    g547(.A1(new_n734_), .A2(G78gat), .A3(new_n458_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n731_), .A2(new_n664_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(G78gat), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n751_), .A2(KEYINPUT50), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n751_), .A2(KEYINPUT50), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n749_), .B1(new_n752_), .B2(new_n753_), .ZN(G1335gat));
  NAND3_X1  g553(.A1(new_n733_), .A2(new_n643_), .A3(new_n671_), .ZN(new_n755_));
  OR2_X1    g554(.A1(new_n755_), .A2(KEYINPUT116), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(KEYINPUT116), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n758_), .A2(new_n580_), .A3(new_n508_), .ZN(new_n759_));
  AND4_X1   g558(.A1(new_n560_), .A2(new_n700_), .A3(new_n539_), .A4(new_n643_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(new_n508_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n759_), .B1(new_n762_), .B2(new_n580_), .ZN(G1336gat));
  NAND3_X1  g562(.A1(new_n758_), .A2(new_n581_), .A3(new_n648_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n760_), .A2(new_n648_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n764_), .B1(new_n766_), .B2(new_n581_), .ZN(G1337gat));
  NAND2_X1  g566(.A1(new_n498_), .A2(new_n576_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n768_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT117), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n769_), .B(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(G99gat), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n772_), .B1(new_n760_), .B2(new_n498_), .ZN(new_n773_));
  OR3_X1    g572(.A1(new_n771_), .A2(KEYINPUT51), .A3(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(KEYINPUT51), .B1(new_n771_), .B2(new_n773_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(G1338gat));
  NAND3_X1  g575(.A1(new_n758_), .A2(new_n664_), .A3(new_n577_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n760_), .A2(new_n664_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n778_), .A2(new_n779_), .A3(G106gat), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n779_), .B1(new_n778_), .B2(G106gat), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n777_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT53), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT53), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n777_), .B(new_n784_), .C1(new_n780_), .C2(new_n781_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n785_), .ZN(G1339gat));
  NAND2_X1  g585(.A1(new_n526_), .A2(new_n527_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n532_), .A2(new_n528_), .A3(new_n523_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n787_), .A2(new_n788_), .A3(new_n538_), .ZN(new_n789_));
  OR2_X1    g588(.A1(new_n789_), .A2(KEYINPUT119), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n534_), .A2(new_n537_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(KEYINPUT119), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n790_), .A2(new_n791_), .A3(new_n792_), .ZN(new_n793_));
  OR3_X1    g592(.A1(new_n596_), .A2(KEYINPUT121), .A3(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(KEYINPUT121), .B1(new_n596_), .B2(new_n793_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT55), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n591_), .A2(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(KEYINPUT55), .B1(new_n588_), .B2(new_n590_), .ZN(new_n799_));
  AOI22_X1  g598(.A1(new_n798_), .A2(new_n799_), .B1(new_n590_), .B2(new_n588_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT56), .ZN(new_n801_));
  INV_X1    g600(.A(new_n566_), .ZN(new_n802_));
  NOR3_X1   g601(.A1(new_n800_), .A2(new_n801_), .A3(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n588_), .A2(new_n590_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n799_), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n588_), .A2(KEYINPUT55), .A3(new_n590_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n804_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT56), .B1(new_n807_), .B2(new_n566_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n796_), .B1(new_n803_), .B2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT58), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n796_), .B(KEYINPUT58), .C1(new_n808_), .C2(new_n803_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n811_), .A2(new_n678_), .A3(new_n812_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n596_), .A2(new_n539_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n814_), .B1(new_n803_), .B2(new_n808_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n793_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n602_), .A2(new_n603_), .A3(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n677_), .B1(new_n815_), .B2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT57), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n813_), .A2(new_n819_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n818_), .A2(KEYINPUT57), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n560_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n730_), .B(KEYINPUT118), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n606_), .A2(new_n636_), .A3(new_n823_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n824_), .B(KEYINPUT54), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n822_), .A2(new_n825_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n507_), .A2(new_n508_), .A3(new_n498_), .A4(new_n458_), .ZN(new_n827_));
  XOR2_X1   g626(.A(new_n827_), .B(KEYINPUT122), .Z(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n829_), .A2(KEYINPUT59), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n826_), .A2(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(KEYINPUT120), .B1(new_n818_), .B2(KEYINPUT57), .ZN(new_n832_));
  INV_X1    g631(.A(new_n817_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n814_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n801_), .B1(new_n800_), .B2(new_n802_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n807_), .A2(KEYINPUT56), .A3(new_n566_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n834_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n634_), .B1(new_n833_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT120), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT57), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n838_), .A2(new_n839_), .A3(new_n840_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n832_), .A2(new_n841_), .A3(new_n813_), .A4(new_n819_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n560_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n829_), .B1(new_n843_), .B2(new_n825_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT59), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n831_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(G113gat), .B1(new_n846_), .B2(new_n539_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n843_), .A2(new_n825_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n828_), .ZN(new_n849_));
  OR2_X1    g648(.A1(new_n539_), .A2(G113gat), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n847_), .B1(new_n849_), .B2(new_n850_), .ZN(G1340gat));
  OAI21_X1  g650(.A(G120gat), .B1(new_n846_), .B2(new_n606_), .ZN(new_n852_));
  INV_X1    g651(.A(G120gat), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n853_), .B1(new_n606_), .B2(KEYINPUT60), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n854_), .B1(KEYINPUT60), .B2(new_n853_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n852_), .B1(new_n849_), .B2(new_n855_), .ZN(G1341gat));
  OAI21_X1  g655(.A(G127gat), .B1(new_n846_), .B2(new_n560_), .ZN(new_n857_));
  OR2_X1    g656(.A1(new_n560_), .A2(G127gat), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n849_), .B2(new_n858_), .ZN(G1342gat));
  OAI21_X1  g658(.A(G134gat), .B1(new_n846_), .B2(new_n636_), .ZN(new_n860_));
  OR3_X1    g659(.A1(new_n849_), .A2(G134gat), .A3(new_n634_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT123), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT123), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n860_), .A2(new_n861_), .A3(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n863_), .A2(new_n865_), .ZN(G1343gat));
  XNOR2_X1  g665(.A(KEYINPUT124), .B(G141gat), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n498_), .A2(new_n458_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n648_), .A2(new_n413_), .ZN(new_n870_));
  AND3_X1   g669(.A1(new_n848_), .A2(new_n869_), .A3(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT125), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n871_), .A2(new_n872_), .A3(new_n729_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n872_), .B1(new_n871_), .B2(new_n729_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n868_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n875_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n877_), .A2(new_n873_), .A3(new_n867_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n878_), .ZN(G1344gat));
  NAND2_X1  g678(.A1(new_n871_), .A2(new_n643_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g680(.A1(new_n871_), .A2(new_n561_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(KEYINPUT61), .B(G155gat), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n882_), .B(new_n883_), .ZN(G1346gat));
  INV_X1    g683(.A(new_n871_), .ZN(new_n885_));
  OAI21_X1  g684(.A(G162gat), .B1(new_n885_), .B2(new_n636_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n871_), .A2(new_n349_), .A3(new_n677_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(G1347gat));
  AOI21_X1  g687(.A(new_n664_), .B1(new_n822_), .B2(new_n825_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n507_), .A2(new_n693_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  OAI21_X1  g690(.A(G169gat), .B1(new_n891_), .B2(new_n539_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT62), .ZN(new_n893_));
  OR2_X1    g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n891_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n895_), .A2(new_n242_), .A3(new_n729_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n892_), .A2(new_n893_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n894_), .A2(new_n896_), .A3(new_n897_), .ZN(G1348gat));
  AOI21_X1  g697(.A(G176gat), .B1(new_n895_), .B2(new_n643_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n664_), .B1(new_n843_), .B2(new_n825_), .ZN(new_n900_));
  NOR4_X1   g699(.A1(new_n606_), .A2(new_n222_), .A3(new_n507_), .A4(new_n693_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n899_), .B1(new_n900_), .B2(new_n901_), .ZN(G1349gat));
  NAND2_X1  g701(.A1(new_n890_), .A2(new_n561_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n903_), .ZN(new_n904_));
  AOI21_X1  g703(.A(G183gat), .B1(new_n900_), .B2(new_n904_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n903_), .A2(new_n230_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n905_), .B1(new_n889_), .B2(new_n906_), .ZN(G1350gat));
  OAI21_X1  g706(.A(G190gat), .B1(new_n891_), .B2(new_n636_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n677_), .A2(new_n229_), .A3(new_n292_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n891_), .B2(new_n909_), .ZN(G1351gat));
  AND2_X1   g709(.A1(new_n848_), .A2(new_n869_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n507_), .A2(new_n508_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n913_), .A2(new_n539_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(new_n261_), .ZN(G1352gat));
  NAND4_X1  g714(.A1(new_n911_), .A2(new_n266_), .A3(new_n643_), .A4(new_n912_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT126), .ZN(new_n917_));
  NAND4_X1  g716(.A1(new_n848_), .A2(new_n643_), .A3(new_n869_), .A4(new_n912_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(new_n246_), .ZN(new_n919_));
  AND3_X1   g718(.A1(new_n916_), .A2(new_n917_), .A3(new_n919_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n917_), .B1(new_n916_), .B2(new_n919_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n920_), .A2(new_n921_), .ZN(G1353gat));
  NAND3_X1  g721(.A1(new_n911_), .A2(new_n561_), .A3(new_n912_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n924_));
  AND2_X1   g723(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n925_));
  NOR3_X1   g724(.A1(new_n923_), .A2(new_n924_), .A3(new_n925_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n926_), .B1(new_n923_), .B2(new_n924_), .ZN(G1354gat));
  INV_X1    g726(.A(G218gat), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n677_), .A2(new_n928_), .ZN(new_n929_));
  AND4_X1   g728(.A1(new_n678_), .A2(new_n848_), .A3(new_n869_), .A4(new_n912_), .ZN(new_n930_));
  OAI22_X1  g729(.A1(new_n913_), .A2(new_n929_), .B1(new_n930_), .B2(new_n928_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n931_), .A2(KEYINPUT127), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT127), .ZN(new_n933_));
  OAI221_X1 g732(.A(new_n933_), .B1(new_n930_), .B2(new_n928_), .C1(new_n913_), .C2(new_n929_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n932_), .A2(new_n934_), .ZN(G1355gat));
endmodule


