//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 1 1 0 1 0 0 1 1 1 0 1 0 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 1 0 0 1 1 0 0 1 0 1 1 0 0 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n699_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n754_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n839_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n857_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_;
  XNOR2_X1  g000(.A(KEYINPUT88), .B(G176gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT22), .B(G169gat), .ZN(new_n203_));
  AOI22_X1  g002(.A1(new_n202_), .A2(new_n203_), .B1(G169gat), .B2(G176gat), .ZN(new_n204_));
  OR2_X1    g003(.A1(new_n204_), .A2(KEYINPUT89), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(KEYINPUT89), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT23), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT87), .B(G183gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n208_), .B1(G190gat), .B2(new_n209_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n205_), .A2(new_n206_), .A3(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT26), .B(G190gat), .ZN(new_n212_));
  AND2_X1   g011(.A1(new_n209_), .A2(KEYINPUT25), .ZN(new_n213_));
  NOR2_X1   g012(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n212_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n207_), .B(KEYINPUT23), .ZN(new_n216_));
  INV_X1    g015(.A(G169gat), .ZN(new_n217_));
  INV_X1    g016(.A(G176gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220_));
  AND3_X1   g019(.A1(new_n219_), .A2(KEYINPUT24), .A3(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n219_), .A2(KEYINPUT24), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n215_), .A2(new_n216_), .A3(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n211_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  XOR2_X1   g025(.A(G211gat), .B(G218gat), .Z(new_n227_));
  INV_X1    g026(.A(G197gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(G204gat), .ZN(new_n229_));
  INV_X1    g028(.A(G204gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(G197gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n227_), .B1(KEYINPUT21), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT97), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n229_), .B(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT96), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n231_), .A2(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n230_), .A2(KEYINPUT96), .A3(G197gat), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n235_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n233_), .B1(new_n239_), .B2(KEYINPUT21), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(KEYINPUT21), .A3(new_n227_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n226_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT20), .ZN(new_n245_));
  INV_X1    g044(.A(new_n212_), .ZN(new_n246_));
  XOR2_X1   g045(.A(KEYINPUT25), .B(G183gat), .Z(new_n247_));
  OAI211_X1 g046(.A(new_n223_), .B(new_n216_), .C1(new_n246_), .C2(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n208_), .B1(G183gat), .B2(G190gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(new_n204_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n245_), .B1(new_n242_), .B2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n244_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G226gat), .A2(G233gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(KEYINPUT19), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n225_), .A2(new_n242_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n240_), .A2(new_n241_), .A3(new_n250_), .A4(new_n248_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n255_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n259_), .A2(KEYINPUT20), .A3(new_n260_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n258_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G8gat), .B(G36gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT18), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G64gat), .B(G92gat), .ZN(new_n266_));
  XOR2_X1   g065(.A(new_n265_), .B(new_n266_), .Z(new_n267_));
  NAND3_X1  g066(.A1(new_n256_), .A2(new_n263_), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n267_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n260_), .B1(new_n244_), .B2(new_n252_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n269_), .B1(new_n270_), .B2(new_n262_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n268_), .A2(new_n271_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n272_), .A2(KEYINPUT27), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT103), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n268_), .A2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT102), .B(KEYINPUT20), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n259_), .A2(new_n276_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n255_), .B1(new_n258_), .B2(new_n277_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n278_), .B1(new_n255_), .B2(new_n253_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(new_n269_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n268_), .A2(new_n274_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n275_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n273_), .B1(new_n282_), .B2(KEYINPUT27), .ZN(new_n283_));
  XOR2_X1   g082(.A(G155gat), .B(G162gat), .Z(new_n284_));
  NAND3_X1  g083(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n285_));
  XOR2_X1   g084(.A(new_n285_), .B(KEYINPUT94), .Z(new_n286_));
  OR2_X1    g085(.A1(G141gat), .A2(G148gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT3), .ZN(new_n288_));
  OR3_X1    g087(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G141gat), .A2(G148gat), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT93), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n290_), .B1(new_n291_), .B2(KEYINPUT2), .ZN(new_n292_));
  AND2_X1   g091(.A1(new_n291_), .A2(KEYINPUT2), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n288_), .B(new_n289_), .C1(new_n292_), .C2(new_n293_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n284_), .B1(new_n286_), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT1), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n284_), .A2(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n298_));
  NAND4_X1  g097(.A1(new_n297_), .A2(new_n298_), .A3(new_n287_), .A4(new_n290_), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n295_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT29), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT28), .ZN(new_n303_));
  XOR2_X1   g102(.A(G22gat), .B(G50gat), .Z(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n300_), .ZN(new_n307_));
  AOI211_X1 g106(.A(KEYINPUT95), .B(new_n243_), .C1(KEYINPUT29), .C2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G78gat), .B(G106gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT98), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G228gat), .A2(G233gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n308_), .B(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n306_), .A2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n308_), .B(new_n312_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(new_n305_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n283_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G227gat), .A2(G233gat), .ZN(new_n320_));
  INV_X1    g119(.A(G71gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(G99gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n225_), .B(new_n323_), .ZN(new_n324_));
  XOR2_X1   g123(.A(KEYINPUT92), .B(KEYINPUT31), .Z(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n324_), .B(new_n326_), .ZN(new_n327_));
  XOR2_X1   g126(.A(G127gat), .B(G134gat), .Z(new_n328_));
  XOR2_X1   g127(.A(G113gat), .B(G120gat), .Z(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT91), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G127gat), .B(G134gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G113gat), .B(G120gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  XOR2_X1   g133(.A(new_n331_), .B(new_n334_), .Z(new_n335_));
  XNOR2_X1  g134(.A(G15gat), .B(G43gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT90), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT30), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n335_), .B(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n327_), .B(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(KEYINPUT4), .B1(new_n307_), .B2(new_n335_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n330_), .A2(new_n334_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT99), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(new_n300_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT100), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n307_), .A2(new_n335_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT100), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n343_), .A2(new_n300_), .A3(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n345_), .A2(new_n346_), .A3(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n341_), .B1(new_n349_), .B2(KEYINPUT4), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G225gat), .A2(G233gat), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n351_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n349_), .A2(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G1gat), .B(G29gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(G85gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT0), .B(G57gat), .ZN(new_n358_));
  XOR2_X1   g157(.A(new_n357_), .B(new_n358_), .Z(new_n359_));
  NAND2_X1  g158(.A1(new_n355_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n359_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n361_), .B1(new_n352_), .B2(new_n354_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n340_), .A2(new_n360_), .A3(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(KEYINPUT105), .B1(new_n319_), .B2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT105), .ZN(new_n366_));
  NOR4_X1   g165(.A1(new_n283_), .A2(new_n363_), .A3(new_n366_), .A4(new_n318_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n365_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n340_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(KEYINPUT101), .A2(KEYINPUT33), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n360_), .A2(new_n370_), .ZN(new_n371_));
  NOR4_X1   g170(.A1(new_n352_), .A2(new_n361_), .A3(new_n354_), .A4(new_n370_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n350_), .A2(new_n353_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n361_), .B1(new_n349_), .B2(new_n351_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n376_), .A2(new_n272_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n371_), .A2(new_n373_), .A3(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n360_), .A2(new_n362_), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n267_), .A2(KEYINPUT32), .ZN(new_n380_));
  NOR3_X1   g179(.A1(new_n270_), .A2(new_n262_), .A3(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n381_), .B1(new_n380_), .B2(new_n279_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n379_), .A2(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n318_), .B1(new_n378_), .B2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n318_), .A2(new_n362_), .A3(new_n360_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n283_), .A2(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n369_), .B1(new_n384_), .B2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT104), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT104), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n389_), .B(new_n369_), .C1(new_n384_), .C2(new_n386_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n368_), .B1(new_n388_), .B2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G1gat), .B(G8gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(KEYINPUT81), .ZN(new_n393_));
  INV_X1    g192(.A(G15gat), .ZN(new_n394_));
  INV_X1    g193(.A(G22gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G15gat), .A2(G22gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G1gat), .A2(G8gat), .ZN(new_n398_));
  AOI22_X1  g197(.A1(new_n396_), .A2(new_n397_), .B1(KEYINPUT14), .B2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n393_), .B(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G29gat), .B(G36gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G43gat), .B(G50gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n401_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n405_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n404_), .B(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(new_n400_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n407_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G229gat), .A2(G233gat), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n411_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT15), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n406_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n409_), .A2(KEYINPUT15), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n416_), .A2(new_n417_), .A3(new_n400_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n413_), .B1(new_n401_), .B2(new_n406_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n414_), .A2(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G113gat), .B(G141gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G169gat), .B(G197gat), .ZN(new_n423_));
  XOR2_X1   g222(.A(new_n422_), .B(new_n423_), .Z(new_n424_));
  XOR2_X1   g223(.A(new_n424_), .B(KEYINPUT85), .Z(new_n425_));
  NAND2_X1  g224(.A1(new_n421_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT86), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n414_), .A2(new_n420_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n427_), .B1(new_n428_), .B2(new_n424_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n424_), .ZN(new_n430_));
  NOR3_X1   g229(.A1(new_n421_), .A2(KEYINPUT86), .A3(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n426_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n391_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(G85gat), .ZN(new_n435_));
  INV_X1    g234(.A(G92gat), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(G85gat), .A2(G92gat), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G99gat), .A2(G106gat), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT67), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n441_), .A2(KEYINPUT6), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT6), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n443_), .A2(KEYINPUT67), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n440_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(KEYINPUT67), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n441_), .A2(KEYINPUT6), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n446_), .A2(new_n447_), .A3(G99gat), .A4(G106gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n445_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT69), .ZN(new_n450_));
  NOR2_X1   g249(.A1(G99gat), .A2(G106gat), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n450_), .B1(new_n451_), .B2(KEYINPUT68), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT7), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT68), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n454_), .B1(new_n453_), .B2(KEYINPUT69), .ZN(new_n455_));
  AOI22_X1  g254(.A1(new_n452_), .A2(new_n453_), .B1(new_n451_), .B2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n439_), .B1(new_n449_), .B2(new_n456_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(KEYINPUT70), .A2(KEYINPUT8), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(KEYINPUT70), .A2(KEYINPUT8), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n457_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n438_), .B1(new_n437_), .B2(KEYINPUT9), .ZN(new_n462_));
  XOR2_X1   g261(.A(KEYINPUT66), .B(G92gat), .Z(new_n463_));
  NOR2_X1   g262(.A1(new_n463_), .A2(new_n435_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(KEYINPUT65), .B(KEYINPUT9), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n462_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  XOR2_X1   g265(.A(KEYINPUT64), .B(G106gat), .Z(new_n467_));
  XNOR2_X1  g266(.A(KEYINPUT10), .B(G99gat), .ZN(new_n468_));
  OR2_X1    g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n449_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n466_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n454_), .B1(G99gat), .B2(G106gat), .ZN(new_n472_));
  AOI21_X1  g271(.A(KEYINPUT7), .B1(new_n472_), .B2(new_n450_), .ZN(new_n473_));
  AOI21_X1  g272(.A(KEYINPUT68), .B1(new_n450_), .B2(KEYINPUT7), .ZN(new_n474_));
  OR2_X1    g273(.A1(G99gat), .A2(G106gat), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n448_), .B(new_n445_), .C1(new_n473_), .C2(new_n476_), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n477_), .A2(KEYINPUT70), .A3(KEYINPUT8), .A4(new_n439_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n461_), .A2(new_n471_), .A3(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(G64gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(G57gat), .ZN(new_n481_));
  INV_X1    g280(.A(G57gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(G64gat), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n481_), .A2(new_n483_), .A3(KEYINPUT11), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT71), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G57gat), .B(G64gat), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT71), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n486_), .A2(new_n487_), .A3(KEYINPUT11), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n485_), .A2(new_n488_), .ZN(new_n489_));
  XOR2_X1   g288(.A(G71gat), .B(G78gat), .Z(new_n490_));
  OAI21_X1  g289(.A(new_n490_), .B1(KEYINPUT11), .B2(new_n486_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n489_), .A2(new_n491_), .ZN(new_n492_));
  OR2_X1    g291(.A1(new_n486_), .A2(KEYINPUT11), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n493_), .A2(new_n485_), .A3(new_n488_), .A4(new_n490_), .ZN(new_n494_));
  AND2_X1   g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n479_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT12), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n495_), .A2(new_n461_), .A3(new_n471_), .A4(new_n478_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G230gat), .A2(G233gat), .ZN(new_n501_));
  AND2_X1   g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n471_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n460_), .ZN(new_n504_));
  AOI211_X1 g303(.A(new_n458_), .B(new_n504_), .C1(new_n477_), .C2(new_n439_), .ZN(new_n505_));
  AND4_X1   g304(.A1(KEYINPUT70), .A2(new_n477_), .A3(KEYINPUT8), .A4(new_n439_), .ZN(new_n506_));
  OAI21_X1  g305(.A(KEYINPUT72), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT72), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n461_), .A2(new_n508_), .A3(new_n478_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n503_), .B1(new_n507_), .B2(new_n509_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n495_), .A2(new_n498_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  OAI211_X1 g311(.A(new_n499_), .B(new_n502_), .C1(new_n510_), .C2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n497_), .A2(new_n500_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n501_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n513_), .A2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G120gat), .B(G148gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT5), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G176gat), .B(G204gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT73), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n517_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT74), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n513_), .A2(new_n516_), .A3(new_n521_), .ZN(new_n526_));
  AND3_X1   g325(.A1(new_n524_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n525_), .B1(new_n524_), .B2(new_n526_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  OR2_X1    g328(.A1(new_n529_), .A2(KEYINPUT13), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(KEYINPUT13), .ZN(new_n531_));
  AND2_X1   g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT75), .ZN(new_n533_));
  OR2_X1    g332(.A1(new_n479_), .A2(new_n409_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G232gat), .A2(G233gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT34), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT35), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n534_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n416_), .A2(new_n417_), .ZN(new_n542_));
  NOR3_X1   g341(.A1(new_n510_), .A2(KEYINPUT78), .A3(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT78), .ZN(new_n544_));
  AND3_X1   g343(.A1(new_n461_), .A2(new_n508_), .A3(new_n478_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n508_), .B1(new_n461_), .B2(new_n478_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n471_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n406_), .B(KEYINPUT15), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n544_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n541_), .B1(new_n543_), .B2(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n537_), .A2(new_n538_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(KEYINPUT78), .B1(new_n510_), .B2(new_n542_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n547_), .A2(new_n548_), .A3(new_n544_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n551_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n555_), .A2(new_n556_), .A3(new_n541_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G190gat), .B(G218gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G134gat), .B(G162gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  OR2_X1    g359(.A1(new_n560_), .A2(KEYINPUT36), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n561_), .B(KEYINPUT79), .Z(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n552_), .A2(new_n557_), .A3(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT80), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT80), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n552_), .A2(new_n557_), .A3(new_n566_), .A4(new_n563_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n560_), .B(KEYINPUT36), .Z(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n570_), .B1(new_n552_), .B2(new_n557_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(KEYINPUT37), .B1(new_n568_), .B2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT37), .ZN(new_n574_));
  AOI211_X1 g373(.A(new_n574_), .B(new_n571_), .C1(new_n565_), .C2(new_n567_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n573_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(G127gat), .B(G155gat), .Z(new_n578_));
  XNOR2_X1  g377(.A(G183gat), .B(G211gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  XOR2_X1   g379(.A(KEYINPUT83), .B(KEYINPUT16), .Z(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(KEYINPUT17), .ZN(new_n583_));
  NAND2_X1  g382(.A1(G231gat), .A2(G233gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT82), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  AND3_X1   g385(.A1(new_n583_), .A2(KEYINPUT84), .A3(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n586_), .B1(new_n583_), .B2(KEYINPUT84), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(new_n495_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n496_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(new_n400_), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n582_), .A2(KEYINPUT17), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n590_), .A2(new_n401_), .A3(new_n591_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n593_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n577_), .A2(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n434_), .A2(new_n533_), .A3(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n379_), .ZN(new_n600_));
  NOR3_X1   g399(.A1(new_n599_), .A2(G1gat), .A3(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(G1gat), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n532_), .A2(new_n433_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(new_n596_), .ZN(new_n606_));
  NOR3_X1   g405(.A1(new_n372_), .A2(new_n376_), .A3(new_n272_), .ZN(new_n607_));
  AOI22_X1  g406(.A1(new_n607_), .A2(new_n371_), .B1(new_n379_), .B2(new_n382_), .ZN(new_n608_));
  OAI22_X1  g407(.A1(new_n608_), .A2(new_n318_), .B1(new_n283_), .B2(new_n385_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n389_), .B1(new_n609_), .B2(new_n369_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n390_), .ZN(new_n611_));
  OAI22_X1  g410(.A1(new_n610_), .A2(new_n611_), .B1(new_n365_), .B2(new_n367_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n556_), .B1(new_n555_), .B2(new_n541_), .ZN(new_n613_));
  AOI211_X1 g412(.A(new_n551_), .B(new_n540_), .C1(new_n553_), .C2(new_n554_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n566_), .B1(new_n615_), .B2(new_n563_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n567_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n572_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n612_), .A2(KEYINPUT107), .A3(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT107), .ZN(new_n620_));
  INV_X1    g419(.A(new_n618_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n620_), .B1(new_n391_), .B2(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n606_), .B1(new_n619_), .B2(new_n622_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n623_), .A2(new_n379_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n603_), .B1(new_n604_), .B2(new_n624_), .ZN(G1324gat));
  INV_X1    g424(.A(KEYINPUT40), .ZN(new_n626_));
  INV_X1    g425(.A(new_n606_), .ZN(new_n627_));
  AOI21_X1  g426(.A(KEYINPUT107), .B1(new_n612_), .B2(new_n618_), .ZN(new_n628_));
  NOR3_X1   g427(.A1(new_n391_), .A2(new_n621_), .A3(new_n620_), .ZN(new_n629_));
  OAI211_X1 g428(.A(new_n283_), .B(new_n627_), .C1(new_n628_), .C2(new_n629_), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n630_), .A2(KEYINPUT108), .A3(G8gat), .ZN(new_n631_));
  AOI21_X1  g430(.A(KEYINPUT108), .B1(new_n630_), .B2(G8gat), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT39), .ZN(new_n633_));
  NOR3_X1   g432(.A1(new_n631_), .A2(new_n632_), .A3(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n633_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n283_), .ZN(new_n636_));
  NOR3_X1   g435(.A1(new_n599_), .A2(G8gat), .A3(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n635_), .A2(new_n638_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n626_), .B1(new_n634_), .B2(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n637_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n632_), .A2(new_n633_), .ZN(new_n642_));
  OAI211_X1 g441(.A(KEYINPUT40), .B(new_n641_), .C1(new_n642_), .C2(new_n631_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n640_), .A2(new_n643_), .ZN(G1325gat));
  INV_X1    g443(.A(new_n599_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n645_), .A2(new_n394_), .A3(new_n340_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n623_), .A2(new_n340_), .ZN(new_n647_));
  AND3_X1   g446(.A1(new_n647_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n648_));
  AOI21_X1  g447(.A(KEYINPUT41), .B1(new_n647_), .B2(G15gat), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n646_), .B1(new_n648_), .B2(new_n649_), .ZN(G1326gat));
  NAND3_X1  g449(.A1(new_n645_), .A2(new_n395_), .A3(new_n318_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT42), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n623_), .A2(new_n318_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n652_), .B1(new_n653_), .B2(G22gat), .ZN(new_n654_));
  AOI211_X1 g453(.A(KEYINPUT42), .B(new_n395_), .C1(new_n623_), .C2(new_n318_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n651_), .B1(new_n654_), .B2(new_n655_), .ZN(G1327gat));
  NAND2_X1  g455(.A1(new_n621_), .A2(new_n597_), .ZN(new_n657_));
  NOR4_X1   g456(.A1(new_n391_), .A2(new_n433_), .A3(new_n532_), .A4(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(G29gat), .B1(new_n658_), .B2(new_n379_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT43), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n612_), .A2(new_n660_), .A3(new_n577_), .ZN(new_n661_));
  OAI21_X1  g460(.A(KEYINPUT43), .B1(new_n391_), .B2(new_n576_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NOR3_X1   g462(.A1(new_n532_), .A2(new_n596_), .A3(new_n433_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n663_), .A2(KEYINPUT44), .A3(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(KEYINPUT44), .B1(new_n663_), .B2(new_n664_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n379_), .A2(G29gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n659_), .B1(new_n668_), .B2(new_n669_), .ZN(G1328gat));
  INV_X1    g469(.A(G36gat), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n658_), .A2(new_n671_), .A3(new_n283_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n672_), .B(new_n673_), .Z(new_n674_));
  NOR3_X1   g473(.A1(new_n666_), .A2(new_n636_), .A3(new_n667_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n674_), .B1(new_n675_), .B2(new_n671_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT46), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  OAI211_X1 g477(.A(new_n674_), .B(KEYINPUT46), .C1(new_n675_), .C2(new_n671_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(G1329gat));
  AOI21_X1  g479(.A(new_n660_), .B1(new_n612_), .B2(new_n577_), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n391_), .A2(KEYINPUT43), .A3(new_n576_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n664_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(G43gat), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n369_), .A2(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n685_), .A2(new_n665_), .A3(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT110), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n685_), .A2(KEYINPUT110), .A3(new_n665_), .A4(new_n687_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n658_), .A2(new_n340_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(new_n686_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n690_), .A2(new_n691_), .A3(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(KEYINPUT47), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT47), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n690_), .A2(new_n696_), .A3(new_n691_), .A4(new_n693_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(G1330gat));
  AOI21_X1  g497(.A(G50gat), .B1(new_n658_), .B2(new_n318_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n318_), .A2(G50gat), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n668_), .B2(new_n700_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT111), .ZN(G1331gat));
  NAND2_X1  g501(.A1(new_n433_), .A2(new_n596_), .ZN(new_n703_));
  AOI211_X1 g502(.A(new_n533_), .B(new_n703_), .C1(new_n619_), .C2(new_n622_), .ZN(new_n704_));
  OAI21_X1  g503(.A(G57gat), .B1(new_n600_), .B2(KEYINPUT113), .ZN(new_n705_));
  OAI211_X1 g504(.A(new_n704_), .B(new_n705_), .C1(KEYINPUT113), .C2(G57gat), .ZN(new_n706_));
  INV_X1    g505(.A(new_n532_), .ZN(new_n707_));
  NOR3_X1   g506(.A1(new_n577_), .A2(new_n707_), .A3(new_n597_), .ZN(new_n708_));
  OR2_X1    g507(.A1(new_n708_), .A2(KEYINPUT112), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n391_), .A2(new_n432_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(KEYINPUT112), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n709_), .A2(new_n710_), .A3(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n482_), .B1(new_n712_), .B2(new_n600_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n706_), .A2(new_n713_), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT114), .Z(G1332gat));
  INV_X1    g514(.A(new_n712_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n716_), .A2(new_n480_), .A3(new_n283_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT48), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n704_), .A2(new_n283_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n718_), .B1(new_n719_), .B2(G64gat), .ZN(new_n720_));
  AOI211_X1 g519(.A(KEYINPUT48), .B(new_n480_), .C1(new_n704_), .C2(new_n283_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n717_), .B1(new_n720_), .B2(new_n721_), .ZN(G1333gat));
  NAND3_X1  g521(.A1(new_n716_), .A2(new_n321_), .A3(new_n340_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n704_), .A2(new_n340_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(KEYINPUT115), .B(KEYINPUT49), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n724_), .A2(G71gat), .A3(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n724_), .B2(G71gat), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n723_), .B1(new_n726_), .B2(new_n727_), .ZN(G1334gat));
  INV_X1    g527(.A(G78gat), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n716_), .A2(new_n729_), .A3(new_n318_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT50), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n704_), .A2(new_n318_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n731_), .B1(new_n732_), .B2(G78gat), .ZN(new_n733_));
  AOI211_X1 g532(.A(KEYINPUT50), .B(new_n729_), .C1(new_n704_), .C2(new_n318_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n730_), .B1(new_n733_), .B2(new_n734_), .ZN(G1335gat));
  NOR3_X1   g534(.A1(new_n707_), .A2(new_n596_), .A3(new_n432_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n663_), .A2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT116), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n736_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT116), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n739_), .A2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT117), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n739_), .A2(KEYINPUT117), .A3(new_n742_), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n745_), .A2(new_n379_), .A3(new_n746_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n533_), .A2(new_n657_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n710_), .A2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n379_), .A2(new_n435_), .ZN(new_n750_));
  OAI22_X1  g549(.A1(new_n747_), .A2(new_n435_), .B1(new_n749_), .B2(new_n750_), .ZN(G1336gat));
  NOR2_X1   g550(.A1(new_n636_), .A2(new_n463_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n745_), .A2(new_n746_), .A3(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n436_), .B1(new_n749_), .B2(new_n636_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n753_), .A2(new_n754_), .ZN(G1337gat));
  OR3_X1    g554(.A1(new_n749_), .A2(new_n468_), .A3(new_n369_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n369_), .B1(new_n739_), .B2(new_n742_), .ZN(new_n757_));
  INV_X1    g556(.A(G99gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n756_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(KEYINPUT51), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT51), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n761_), .B(new_n756_), .C1(new_n757_), .C2(new_n758_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(G1338gat));
  INV_X1    g562(.A(new_n318_), .ZN(new_n764_));
  OR3_X1    g563(.A1(new_n749_), .A2(new_n467_), .A3(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n741_), .A2(new_n318_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n766_), .A2(new_n767_), .A3(G106gat), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n766_), .B2(G106gat), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n765_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g570(.A1(new_n428_), .A2(new_n427_), .A3(new_n424_), .ZN(new_n772_));
  OAI21_X1  g571(.A(KEYINPUT86), .B1(new_n421_), .B2(new_n430_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n418_), .A2(new_n407_), .A3(new_n413_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n411_), .A2(new_n412_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(new_n776_), .A3(new_n430_), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n774_), .A2(new_n526_), .A3(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT55), .ZN(new_n779_));
  OAI21_X1  g578(.A(KEYINPUT118), .B1(new_n513_), .B2(new_n779_), .ZN(new_n780_));
  AOI22_X1  g579(.A1(new_n547_), .A2(new_n511_), .B1(new_n498_), .B2(new_n497_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT118), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n781_), .A2(new_n782_), .A3(KEYINPUT55), .A4(new_n502_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n513_), .A2(new_n779_), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n500_), .B(new_n499_), .C1(new_n510_), .C2(new_n512_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n515_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n780_), .A2(new_n783_), .A3(new_n784_), .A4(new_n786_), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n787_), .A2(KEYINPUT56), .A3(new_n523_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT56), .B1(new_n787_), .B2(new_n523_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n778_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT58), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  OAI211_X1 g591(.A(KEYINPUT58), .B(new_n778_), .C1(new_n788_), .C2(new_n789_), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n792_), .B(new_n793_), .C1(new_n573_), .C2(new_n575_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n432_), .A2(new_n526_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n787_), .A2(new_n523_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT56), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n787_), .A2(KEYINPUT56), .A3(new_n523_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n795_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n774_), .A2(new_n777_), .ZN(new_n801_));
  NOR3_X1   g600(.A1(new_n801_), .A2(new_n527_), .A3(new_n528_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n618_), .B1(new_n800_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT57), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n618_), .B(KEYINPUT57), .C1(new_n800_), .C2(new_n802_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n794_), .A2(new_n805_), .A3(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(KEYINPUT119), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT119), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n794_), .A2(new_n805_), .A3(new_n809_), .A4(new_n806_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n808_), .A2(new_n597_), .A3(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT120), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n703_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n576_), .A2(new_n813_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n814_), .B(KEYINPUT54), .ZN(new_n815_));
  AND3_X1   g614(.A1(new_n811_), .A2(new_n812_), .A3(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n812_), .B1(new_n811_), .B2(new_n815_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n319_), .A2(new_n379_), .A3(new_n340_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(G113gat), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n822_), .A2(new_n823_), .A3(new_n432_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n807_), .A2(new_n597_), .ZN(new_n825_));
  AND2_X1   g624(.A1(new_n815_), .A2(new_n825_), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n826_), .A2(KEYINPUT59), .A3(new_n819_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n827_), .B1(new_n821_), .B2(KEYINPUT59), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n828_), .A2(new_n432_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n824_), .B1(new_n829_), .B2(new_n823_), .ZN(G1340gat));
  INV_X1    g629(.A(G120gat), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n831_), .B1(new_n707_), .B2(KEYINPUT60), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n822_), .B(new_n832_), .C1(KEYINPUT60), .C2(new_n831_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n533_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n828_), .A2(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n833_), .B1(new_n835_), .B2(new_n831_), .ZN(G1341gat));
  INV_X1    g635(.A(G127gat), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n822_), .A2(new_n837_), .A3(new_n596_), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n828_), .A2(new_n596_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n838_), .B1(new_n839_), .B2(new_n837_), .ZN(G1342gat));
  INV_X1    g639(.A(G134gat), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n841_), .B1(new_n821_), .B2(new_n618_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(KEYINPUT121), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT121), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n844_), .B(new_n841_), .C1(new_n821_), .C2(new_n618_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n576_), .A2(new_n841_), .ZN(new_n846_));
  AOI22_X1  g645(.A1(new_n843_), .A2(new_n845_), .B1(new_n828_), .B2(new_n846_), .ZN(G1343gat));
  NAND2_X1  g646(.A1(new_n811_), .A2(new_n815_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(KEYINPUT120), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n811_), .A2(new_n812_), .A3(new_n815_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n764_), .A2(new_n340_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n636_), .A2(new_n852_), .A3(new_n379_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n851_), .A2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n432_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g655(.A1(new_n854_), .A2(new_n834_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g657(.A(KEYINPUT122), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n854_), .A2(new_n859_), .A3(new_n596_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n853_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n818_), .A2(new_n596_), .A3(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT122), .ZN(new_n863_));
  XNOR2_X1  g662(.A(KEYINPUT61), .B(G155gat), .ZN(new_n864_));
  AND3_X1   g663(.A1(new_n860_), .A2(new_n863_), .A3(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n864_), .B1(new_n860_), .B2(new_n863_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n865_), .A2(new_n866_), .ZN(G1346gat));
  AOI21_X1  g666(.A(G162gat), .B1(new_n854_), .B2(new_n621_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n577_), .A2(G162gat), .ZN(new_n869_));
  XOR2_X1   g668(.A(new_n869_), .B(KEYINPUT123), .Z(new_n870_));
  AOI21_X1  g669(.A(new_n868_), .B1(new_n854_), .B2(new_n870_), .ZN(G1347gat));
  NOR2_X1   g670(.A1(new_n636_), .A2(new_n379_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n340_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n826_), .A2(new_n318_), .A3(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n217_), .B1(new_n874_), .B2(new_n432_), .ZN(new_n875_));
  OR2_X1    g674(.A1(new_n875_), .A2(KEYINPUT62), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n874_), .A2(new_n203_), .A3(new_n432_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n875_), .A2(KEYINPUT62), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n876_), .A2(new_n877_), .A3(new_n878_), .ZN(G1348gat));
  NAND2_X1  g678(.A1(new_n874_), .A2(new_n532_), .ZN(new_n880_));
  AND2_X1   g679(.A1(new_n880_), .A2(new_n202_), .ZN(new_n881_));
  OR2_X1    g680(.A1(new_n881_), .A2(KEYINPUT124), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(KEYINPUT124), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n851_), .A2(new_n318_), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n533_), .A2(new_n218_), .A3(new_n873_), .ZN(new_n885_));
  AOI22_X1  g684(.A1(new_n882_), .A2(new_n883_), .B1(new_n884_), .B2(new_n885_), .ZN(G1349gat));
  NOR2_X1   g685(.A1(new_n873_), .A2(new_n597_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n209_), .B1(new_n884_), .B2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n247_), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n826_), .A2(new_n318_), .A3(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n888_), .A2(new_n890_), .ZN(G1350gat));
  NOR2_X1   g690(.A1(new_n618_), .A2(new_n246_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(KEYINPUT125), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n874_), .A2(new_n893_), .ZN(new_n894_));
  AND2_X1   g693(.A1(new_n874_), .A2(new_n577_), .ZN(new_n895_));
  INV_X1    g694(.A(G190gat), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n894_), .B1(new_n895_), .B2(new_n896_), .ZN(G1351gat));
  AND2_X1   g696(.A1(new_n872_), .A2(new_n852_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n849_), .A2(new_n850_), .A3(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT126), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  NAND4_X1  g700(.A1(new_n849_), .A2(KEYINPUT126), .A3(new_n850_), .A4(new_n898_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n433_), .B1(new_n901_), .B2(new_n902_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(new_n228_), .ZN(G1352gat));
  AOI21_X1  g703(.A(new_n533_), .B1(new_n901_), .B2(new_n902_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(new_n230_), .ZN(G1353gat));
  XNOR2_X1  g705(.A(KEYINPUT63), .B(G211gat), .ZN(new_n907_));
  AOI211_X1 g706(.A(new_n597_), .B(new_n907_), .C1(new_n901_), .C2(new_n902_), .ZN(new_n908_));
  AOI21_X1  g707(.A(KEYINPUT126), .B1(new_n818_), .B2(new_n898_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n902_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n596_), .B1(new_n909_), .B2(new_n910_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n908_), .B1(new_n911_), .B2(new_n912_), .ZN(G1354gat));
  NAND2_X1  g712(.A1(new_n577_), .A2(G218gat), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n914_), .B1(new_n901_), .B2(new_n902_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n618_), .B1(new_n901_), .B2(new_n902_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT127), .ZN(new_n917_));
  AOI21_X1  g716(.A(G218gat), .B1(new_n916_), .B2(new_n917_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n621_), .B1(new_n909_), .B2(new_n910_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(KEYINPUT127), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n915_), .B1(new_n918_), .B2(new_n920_), .ZN(G1355gat));
endmodule


