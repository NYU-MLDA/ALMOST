//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 1 1 1 0 0 1 1 0 1 0 0 0 0 0 1 1 0 1 0 0 0 0 1 0 0 0 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 0 1 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n650_, new_n651_, new_n652_, new_n653_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n860_, new_n862_,
    new_n863_, new_n864_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n871_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n883_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n897_, new_n899_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_;
  INV_X1    g000(.A(KEYINPUT97), .ZN(new_n202_));
  XOR2_X1   g001(.A(G190gat), .B(G218gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT73), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G134gat), .B(G162gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT36), .ZN(new_n207_));
  OR3_X1    g006(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT66), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT6), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n212_), .B1(G99gat), .B2(G106gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G99gat), .A2(G106gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n214_), .A2(KEYINPUT6), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n211_), .B1(new_n213_), .B2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(KEYINPUT6), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n212_), .A2(G99gat), .A3(G106gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n217_), .A2(new_n218_), .A3(KEYINPUT66), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n210_), .B1(new_n216_), .B2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G85gat), .B(G92gat), .ZN(new_n221_));
  OR2_X1    g020(.A1(new_n221_), .A2(KEYINPUT8), .ZN(new_n222_));
  INV_X1    g021(.A(new_n209_), .ZN(new_n223_));
  NOR3_X1   g022(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n217_), .A2(new_n218_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n221_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT8), .ZN(new_n228_));
  OAI22_X1  g027(.A1(new_n220_), .A2(new_n222_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT9), .ZN(new_n230_));
  NAND2_X1  g029(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n230_), .B(G92gat), .C1(new_n232_), .C2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT65), .ZN(new_n235_));
  OAI211_X1 g034(.A(new_n234_), .B(new_n235_), .C1(new_n230_), .C2(new_n221_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n230_), .A2(G92gat), .ZN(new_n237_));
  INV_X1    g036(.A(new_n233_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n237_), .B1(new_n238_), .B2(new_n231_), .ZN(new_n239_));
  AND2_X1   g038(.A1(G85gat), .A2(G92gat), .ZN(new_n240_));
  NOR2_X1   g039(.A1(G85gat), .A2(G92gat), .ZN(new_n241_));
  NOR3_X1   g040(.A1(new_n240_), .A2(new_n241_), .A3(new_n230_), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT65), .B1(new_n239_), .B2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n216_), .A2(new_n219_), .ZN(new_n244_));
  XOR2_X1   g043(.A(KEYINPUT10), .B(G99gat), .Z(new_n245_));
  INV_X1    g044(.A(G106gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n236_), .A2(new_n243_), .A3(new_n244_), .A4(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n229_), .A2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G43gat), .B(G50gat), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G29gat), .B(G36gat), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT70), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(G36gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(G29gat), .ZN(new_n256_));
  INV_X1    g055(.A(G29gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(G36gat), .ZN(new_n258_));
  AND3_X1   g057(.A1(new_n256_), .A2(new_n258_), .A3(new_n253_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n251_), .B1(new_n254_), .B2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n256_), .A2(new_n258_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT70), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n252_), .A2(new_n253_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n262_), .A2(new_n263_), .A3(new_n250_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n260_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G232gat), .A2(G233gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT34), .ZN(new_n267_));
  OAI22_X1  g066(.A1(new_n249_), .A2(new_n265_), .B1(KEYINPUT35), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  XOR2_X1   g068(.A(KEYINPUT71), .B(KEYINPUT15), .Z(new_n270_));
  AND3_X1   g069(.A1(new_n260_), .A2(new_n270_), .A3(new_n264_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n270_), .B1(new_n260_), .B2(new_n264_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  AND3_X1   g072(.A1(new_n273_), .A2(KEYINPUT72), .A3(new_n249_), .ZN(new_n274_));
  AOI21_X1  g073(.A(KEYINPUT72), .B1(new_n273_), .B2(new_n249_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n269_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n267_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT35), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n276_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n279_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n273_), .A2(new_n249_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT72), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n273_), .A2(KEYINPUT72), .A3(new_n249_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n281_), .B1(new_n286_), .B2(new_n269_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n207_), .B1(new_n280_), .B2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n276_), .A2(new_n279_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n286_), .A2(new_n281_), .A3(new_n269_), .ZN(new_n290_));
  XOR2_X1   g089(.A(KEYINPUT74), .B(KEYINPUT36), .Z(new_n291_));
  AND2_X1   g090(.A1(new_n206_), .A2(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n289_), .A2(new_n290_), .A3(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n288_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT37), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n295_), .B1(new_n293_), .B2(KEYINPUT75), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  OAI211_X1 g096(.A(new_n288_), .B(new_n293_), .C1(KEYINPUT75), .C2(new_n295_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT77), .ZN(new_n300_));
  XOR2_X1   g099(.A(G71gat), .B(G78gat), .Z(new_n301_));
  XNOR2_X1  g100(.A(G57gat), .B(G64gat), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n301_), .B1(KEYINPUT11), .B2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT67), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n304_), .B1(new_n302_), .B2(KEYINPUT11), .ZN(new_n305_));
  INV_X1    g104(.A(G64gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(G57gat), .ZN(new_n307_));
  INV_X1    g106(.A(G57gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(G64gat), .ZN(new_n309_));
  AND4_X1   g108(.A1(new_n304_), .A2(new_n307_), .A3(new_n309_), .A4(KEYINPUT11), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n303_), .B1(new_n305_), .B2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n307_), .A2(new_n309_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT11), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT67), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n302_), .A2(new_n304_), .A3(KEYINPUT11), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n312_), .A2(new_n313_), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n314_), .A2(new_n315_), .A3(new_n316_), .A4(new_n301_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n311_), .A2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G1gat), .B(G8gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT76), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G15gat), .B(G22gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G1gat), .A2(G8gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(KEYINPUT14), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n321_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n320_), .A2(new_n324_), .ZN(new_n325_));
  OR2_X1    g124(.A1(new_n319_), .A2(KEYINPUT76), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n319_), .A2(KEYINPUT76), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n326_), .A2(new_n323_), .A3(new_n321_), .A4(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n325_), .A2(new_n328_), .ZN(new_n329_));
  AND2_X1   g128(.A1(G231gat), .A2(G233gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n329_), .A2(new_n330_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n318_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n333_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n318_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n335_), .A2(new_n336_), .A3(new_n331_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT68), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n334_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  XOR2_X1   g138(.A(G127gat), .B(G155gat), .Z(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(KEYINPUT16), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G183gat), .B(G211gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT17), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n339_), .A2(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n338_), .B1(new_n334_), .B2(new_n337_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n300_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n347_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n349_), .A2(KEYINPUT77), .A3(new_n345_), .A4(new_n339_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  AND2_X1   g150(.A1(new_n343_), .A2(new_n344_), .ZN(new_n352_));
  OR3_X1    g151(.A1(new_n352_), .A2(new_n345_), .A3(KEYINPUT78), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n334_), .A2(new_n337_), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT78), .B1(new_n352_), .B2(new_n345_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n353_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(KEYINPUT79), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT79), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n353_), .A2(new_n358_), .A3(new_n354_), .A4(new_n355_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n357_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n351_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n299_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(KEYINPUT80), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT13), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n249_), .A2(new_n336_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT12), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n367_), .B1(new_n229_), .B2(new_n248_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n318_), .A2(new_n338_), .ZN(new_n370_));
  AOI21_X1  g169(.A(KEYINPUT68), .B1(new_n311_), .B2(new_n317_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n369_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n229_), .A2(new_n318_), .A3(new_n248_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G230gat), .A2(G233gat), .ZN(new_n374_));
  AND3_X1   g173(.A1(new_n373_), .A2(KEYINPUT69), .A3(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(KEYINPUT69), .B1(new_n373_), .B2(new_n374_), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n368_), .B(new_n372_), .C1(new_n375_), .C2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n366_), .A2(new_n373_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n374_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n377_), .A2(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G120gat), .B(G148gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT5), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G176gat), .B(G204gat), .ZN(new_n384_));
  XOR2_X1   g183(.A(new_n383_), .B(new_n384_), .Z(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  AND2_X1   g185(.A1(new_n381_), .A2(new_n386_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n381_), .A2(new_n386_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n365_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  OR2_X1    g188(.A1(new_n381_), .A2(new_n386_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n381_), .A2(new_n386_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n390_), .A2(KEYINPUT13), .A3(new_n391_), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n389_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT80), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n299_), .A2(new_n394_), .A3(new_n362_), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n364_), .A2(KEYINPUT81), .A3(new_n393_), .A4(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G8gat), .B(G36gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G64gat), .B(G92gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G183gat), .A2(G190gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(KEYINPUT23), .ZN(new_n404_));
  OR2_X1    g203(.A1(G183gat), .A2(G190gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(G169gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n406_), .A2(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(KEYINPUT25), .B(G183gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(KEYINPUT26), .B(G190gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(G169gat), .ZN(new_n413_));
  INV_X1    g212(.A(G176gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  OR2_X1    g214(.A1(new_n415_), .A2(KEYINPUT24), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n412_), .A2(new_n404_), .A3(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G169gat), .A2(G176gat), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n415_), .A2(KEYINPUT24), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT84), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n415_), .A2(KEYINPUT84), .A3(KEYINPUT24), .A4(new_n418_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n409_), .B1(new_n417_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT85), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT21), .ZN(new_n427_));
  XNOR2_X1  g226(.A(KEYINPUT88), .B(G204gat), .ZN(new_n428_));
  INV_X1    g227(.A(G197gat), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(G197gat), .A2(G204gat), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n427_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  XOR2_X1   g231(.A(G211gat), .B(G218gat), .Z(new_n433_));
  NAND2_X1  g232(.A1(new_n428_), .A2(new_n429_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n427_), .B1(G197gat), .B2(G204gat), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n433_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n430_), .A2(new_n431_), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n433_), .A2(KEYINPUT21), .ZN(new_n438_));
  AOI22_X1  g237(.A1(new_n432_), .A2(new_n436_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n409_), .B(KEYINPUT85), .C1(new_n417_), .C2(new_n423_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n426_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n432_), .A2(new_n436_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n437_), .A2(new_n438_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n412_), .A2(new_n404_), .A3(new_n416_), .A4(new_n419_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT91), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(new_n409_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n445_), .A2(KEYINPUT91), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n444_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n441_), .A2(KEYINPUT20), .A3(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G226gat), .A2(G233gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(KEYINPUT19), .ZN(new_n452_));
  OR2_X1    g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n426_), .A2(new_n440_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(new_n444_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n439_), .A2(new_n445_), .A3(new_n409_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(KEYINPUT20), .A3(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(new_n452_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n402_), .B1(new_n453_), .B2(new_n458_), .ZN(new_n459_));
  OR3_X1    g258(.A1(new_n444_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n452_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n455_), .A2(new_n460_), .A3(KEYINPUT20), .A4(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n450_), .A2(new_n452_), .ZN(new_n463_));
  AND3_X1   g262(.A1(new_n462_), .A2(new_n463_), .A3(new_n402_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT27), .ZN(new_n465_));
  NOR3_X1   g264(.A1(new_n459_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n402_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n465_), .B1(new_n464_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT96), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  OAI211_X1 g269(.A(KEYINPUT96), .B(new_n465_), .C1(new_n464_), .C2(new_n467_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n466_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(G141gat), .ZN(new_n473_));
  INV_X1    g272(.A(G148gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G141gat), .A2(G148gat), .ZN(new_n476_));
  NOR2_X1   g275(.A1(G155gat), .A2(G162gat), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT87), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G155gat), .A2(G162gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT1), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n475_), .B(new_n476_), .C1(new_n479_), .C2(new_n481_), .ZN(new_n482_));
  OR3_X1    g281(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT2), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n476_), .A2(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n483_), .A2(new_n485_), .A3(new_n486_), .A4(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n477_), .B(KEYINPUT87), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n488_), .A2(new_n489_), .A3(new_n480_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n482_), .A2(new_n490_), .ZN(new_n491_));
  OAI21_X1  g290(.A(KEYINPUT28), .B1(new_n491_), .B2(KEYINPUT29), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT28), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT29), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n482_), .A2(new_n493_), .A3(new_n494_), .A4(new_n490_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n492_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G228gat), .A2(G233gat), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n497_), .A2(KEYINPUT89), .ZN(new_n498_));
  XOR2_X1   g297(.A(new_n496_), .B(new_n498_), .Z(new_n499_));
  NAND2_X1  g298(.A1(new_n497_), .A2(KEYINPUT89), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n494_), .B1(new_n482_), .B2(new_n490_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n500_), .B1(new_n439_), .B2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G78gat), .B(G106gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT90), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n502_), .A2(new_n505_), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n504_), .B(new_n500_), .C1(new_n439_), .C2(new_n501_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G22gat), .B(G50gat), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n506_), .A2(new_n507_), .A3(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n509_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  AND3_X1   g311(.A1(new_n499_), .A2(new_n510_), .A3(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n499_), .B1(new_n512_), .B2(new_n510_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  XOR2_X1   g314(.A(G127gat), .B(G134gat), .Z(new_n516_));
  XOR2_X1   g315(.A(G113gat), .B(G120gat), .Z(new_n517_));
  XOR2_X1   g316(.A(new_n516_), .B(new_n517_), .Z(new_n518_));
  NAND2_X1  g317(.A1(new_n491_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G225gat), .A2(G233gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n516_), .B(new_n517_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n521_), .A2(new_n482_), .A3(new_n490_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n519_), .A2(new_n520_), .A3(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT93), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n519_), .A2(KEYINPUT4), .A3(new_n522_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n520_), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n525_), .B(new_n526_), .C1(KEYINPUT4), .C2(new_n519_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n524_), .A2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G1gat), .B(G29gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(G85gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(KEYINPUT0), .B(G57gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n528_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n532_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n524_), .A2(new_n534_), .A3(new_n527_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G15gat), .B(G43gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G71gat), .B(G99gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n454_), .B(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(new_n518_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G227gat), .A2(G233gat), .ZN(new_n543_));
  XOR2_X1   g342(.A(new_n543_), .B(KEYINPUT86), .Z(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT30), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT31), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n542_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n542_), .A2(new_n547_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n472_), .A2(new_n515_), .A3(new_n537_), .A4(new_n550_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n515_), .A2(new_n536_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n464_), .A2(new_n467_), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n524_), .A2(new_n527_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT94), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n554_), .A2(new_n555_), .A3(KEYINPUT33), .A4(new_n534_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n519_), .A2(new_n522_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT95), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT95), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n519_), .A2(new_n559_), .A3(new_n522_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n558_), .A2(new_n526_), .A3(new_n560_), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n525_), .B(new_n520_), .C1(KEYINPUT4), .C2(new_n519_), .ZN(new_n562_));
  AND3_X1   g361(.A1(new_n561_), .A2(new_n532_), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT33), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n535_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  OAI21_X1  g364(.A(KEYINPUT94), .B1(new_n535_), .B2(new_n564_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n553_), .A2(new_n556_), .A3(new_n565_), .A4(new_n566_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n402_), .A2(KEYINPUT32), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n462_), .A2(new_n463_), .A3(new_n569_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n453_), .A2(new_n458_), .ZN(new_n571_));
  OAI211_X1 g370(.A(new_n536_), .B(new_n570_), .C1(new_n571_), .C2(new_n569_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n567_), .A2(new_n572_), .ZN(new_n573_));
  AOI22_X1  g372(.A1(new_n472_), .A2(new_n552_), .B1(new_n573_), .B2(new_n515_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n551_), .B1(new_n574_), .B2(new_n550_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n329_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(new_n265_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n329_), .A2(new_n264_), .A3(new_n260_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G229gat), .A2(G233gat), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n273_), .A2(new_n576_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n583_), .A2(new_n578_), .A3(new_n580_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  XOR2_X1   g384(.A(G113gat), .B(G141gat), .Z(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT82), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G169gat), .B(G197gat), .ZN(new_n588_));
  XOR2_X1   g387(.A(new_n587_), .B(new_n588_), .Z(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n585_), .A2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n582_), .A2(new_n584_), .A3(new_n589_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n593_), .B(KEYINPUT83), .Z(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n396_), .A2(new_n575_), .A3(new_n595_), .ZN(new_n596_));
  AOI211_X1 g395(.A(KEYINPUT80), .B(new_n361_), .C1(new_n297_), .C2(new_n298_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n394_), .B1(new_n299_), .B2(new_n362_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(KEYINPUT81), .B1(new_n599_), .B2(new_n393_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n202_), .B1(new_n596_), .B2(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n364_), .A2(new_n393_), .A3(new_n395_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT81), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n472_), .A2(new_n552_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n573_), .A2(new_n515_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n550_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n594_), .B1(new_n609_), .B2(new_n551_), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n604_), .A2(new_n610_), .A3(KEYINPUT97), .A4(new_n396_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n601_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT98), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n601_), .A2(KEYINPUT98), .A3(new_n611_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n537_), .A2(G1gat), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n614_), .A2(new_n615_), .A3(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT38), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n393_), .A2(new_n593_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n620_), .A2(new_n361_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n575_), .A2(new_n294_), .A3(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(G1gat), .B1(new_n622_), .B2(new_n537_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n617_), .A2(new_n618_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n619_), .A2(new_n623_), .A3(new_n624_), .ZN(G1324gat));
  NOR2_X1   g424(.A1(new_n472_), .A2(G8gat), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n614_), .A2(new_n615_), .A3(new_n626_), .ZN(new_n627_));
  OAI21_X1  g426(.A(KEYINPUT99), .B1(new_n622_), .B2(new_n472_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n294_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n629_), .B1(new_n609_), .B2(new_n551_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT99), .ZN(new_n631_));
  INV_X1    g430(.A(new_n472_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n630_), .A2(new_n631_), .A3(new_n632_), .A4(new_n621_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n628_), .A2(new_n633_), .A3(G8gat), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT100), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT100), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n628_), .A2(new_n633_), .A3(new_n636_), .A4(G8gat), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n635_), .A2(KEYINPUT39), .A3(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT39), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n634_), .A2(KEYINPUT100), .A3(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n627_), .A2(new_n638_), .A3(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n641_), .B(new_n642_), .ZN(G1325gat));
  OR3_X1    g442(.A1(new_n612_), .A2(G15gat), .A3(new_n608_), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n644_), .A2(KEYINPUT102), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(KEYINPUT102), .ZN(new_n646_));
  OAI21_X1  g445(.A(G15gat), .B1(new_n622_), .B2(new_n608_), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n647_), .B(KEYINPUT41), .Z(new_n648_));
  NAND3_X1  g447(.A1(new_n645_), .A2(new_n646_), .A3(new_n648_), .ZN(G1326gat));
  OAI21_X1  g448(.A(G22gat), .B1(new_n622_), .B2(new_n515_), .ZN(new_n650_));
  XOR2_X1   g449(.A(KEYINPUT103), .B(KEYINPUT42), .Z(new_n651_));
  XNOR2_X1  g450(.A(new_n650_), .B(new_n651_), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n515_), .A2(G22gat), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n652_), .B1(new_n612_), .B2(new_n653_), .ZN(G1327gat));
  NOR2_X1   g453(.A1(new_n620_), .A2(new_n362_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT43), .ZN(new_n656_));
  INV_X1    g455(.A(new_n299_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n550_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n551_), .ZN(new_n659_));
  OAI211_X1 g458(.A(new_n656_), .B(new_n657_), .C1(new_n658_), .C2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n656_), .B1(new_n575_), .B2(new_n657_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n655_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT44), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  OAI211_X1 g465(.A(KEYINPUT44), .B(new_n655_), .C1(new_n661_), .C2(new_n662_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  NOR3_X1   g467(.A1(new_n666_), .A2(new_n668_), .A3(new_n537_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n362_), .A2(new_n294_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n610_), .A2(new_n393_), .A3(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n536_), .A2(new_n257_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT104), .ZN(new_n673_));
  OAI22_X1  g472(.A1(new_n669_), .A2(new_n257_), .B1(new_n671_), .B2(new_n673_), .ZN(G1328gat));
  NAND2_X1  g473(.A1(new_n632_), .A2(new_n255_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n671_), .A2(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n676_), .B(new_n677_), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n666_), .A2(new_n668_), .A3(new_n472_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n678_), .B1(new_n679_), .B2(new_n255_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT46), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  OAI211_X1 g481(.A(KEYINPUT46), .B(new_n678_), .C1(new_n679_), .C2(new_n255_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(G1329gat));
  AND2_X1   g483(.A1(new_n550_), .A2(G43gat), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n665_), .A2(new_n667_), .A3(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT106), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n665_), .A2(KEYINPUT106), .A3(new_n667_), .A4(new_n685_), .ZN(new_n689_));
  XOR2_X1   g488(.A(KEYINPUT107), .B(G43gat), .Z(new_n690_));
  OAI21_X1  g489(.A(new_n690_), .B1(new_n671_), .B2(new_n608_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n688_), .A2(new_n689_), .A3(new_n691_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g492(.A(new_n671_), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n513_), .A2(new_n514_), .ZN(new_n695_));
  AOI21_X1  g494(.A(G50gat), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n666_), .A2(new_n668_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n695_), .A2(G50gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n696_), .B1(new_n697_), .B2(new_n698_), .ZN(G1331gat));
  NAND2_X1  g498(.A1(new_n575_), .A2(new_n294_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n393_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n701_), .A2(new_n362_), .A3(new_n594_), .ZN(new_n702_));
  OR2_X1    g501(.A1(new_n700_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n704_), .A2(G57gat), .A3(new_n536_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT109), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n393_), .A2(new_n593_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n575_), .A2(new_n707_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n708_), .A2(new_n599_), .ZN(new_n709_));
  OR2_X1    g508(.A1(new_n709_), .A2(KEYINPUT108), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(KEYINPUT108), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n710_), .A2(new_n536_), .A3(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n706_), .B1(new_n308_), .B2(new_n712_), .ZN(G1332gat));
  OAI21_X1  g512(.A(G64gat), .B1(new_n703_), .B2(new_n472_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT48), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n709_), .A2(new_n306_), .A3(new_n632_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1333gat));
  INV_X1    g516(.A(new_n709_), .ZN(new_n718_));
  OR3_X1    g517(.A1(new_n718_), .A2(G71gat), .A3(new_n608_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n704_), .A2(new_n550_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT49), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n720_), .A2(new_n721_), .A3(G71gat), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n721_), .B1(new_n720_), .B2(G71gat), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n719_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT110), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  OAI211_X1 g526(.A(KEYINPUT110), .B(new_n719_), .C1(new_n723_), .C2(new_n724_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1334gat));
  OAI21_X1  g528(.A(G78gat), .B1(new_n703_), .B2(new_n515_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT50), .ZN(new_n731_));
  OR2_X1    g530(.A1(new_n515_), .A2(G78gat), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n731_), .B1(new_n718_), .B2(new_n732_), .ZN(G1335gat));
  NAND2_X1  g532(.A1(new_n708_), .A2(new_n670_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(G85gat), .B1(new_n735_), .B2(new_n536_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n661_), .A2(new_n662_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n707_), .A2(new_n361_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n537_), .B1(new_n238_), .B2(new_n231_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n736_), .B1(new_n739_), .B2(new_n740_), .ZN(G1336gat));
  NAND3_X1  g540(.A1(new_n739_), .A2(G92gat), .A3(new_n632_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n735_), .A2(new_n632_), .ZN(new_n743_));
  INV_X1    g542(.A(G92gat), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n743_), .A2(KEYINPUT111), .A3(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(KEYINPUT111), .B1(new_n743_), .B2(new_n744_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n742_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT112), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  OAI211_X1 g549(.A(KEYINPUT112), .B(new_n742_), .C1(new_n746_), .C2(new_n747_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(G1337gat));
  NAND2_X1  g551(.A1(new_n550_), .A2(new_n245_), .ZN(new_n753_));
  OR2_X1    g552(.A1(new_n734_), .A2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT51), .ZN(new_n755_));
  NOR3_X1   g554(.A1(new_n737_), .A2(new_n608_), .A3(new_n738_), .ZN(new_n756_));
  INV_X1    g555(.A(G99gat), .ZN(new_n757_));
  OAI221_X1 g556(.A(new_n754_), .B1(KEYINPUT113), .B2(new_n755_), .C1(new_n756_), .C2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n755_), .A2(KEYINPUT113), .ZN(new_n759_));
  XOR2_X1   g558(.A(new_n759_), .B(KEYINPUT114), .Z(new_n760_));
  XOR2_X1   g559(.A(new_n758_), .B(new_n760_), .Z(G1338gat));
  XNOR2_X1  g560(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  NOR3_X1   g562(.A1(new_n734_), .A2(G106gat), .A3(new_n515_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT115), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n246_), .B1(new_n739_), .B2(new_n695_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT52), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n765_), .A2(new_n767_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n766_), .A2(KEYINPUT52), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n763_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n769_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n771_), .A2(new_n767_), .A3(new_n765_), .A4(new_n762_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(G1339gat));
  NAND4_X1  g572(.A1(new_n393_), .A2(new_n299_), .A3(new_n594_), .A4(new_n362_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(KEYINPUT117), .A2(KEYINPUT54), .ZN(new_n775_));
  OR2_X1    g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n775_), .ZN(new_n777_));
  AOI22_X1  g576(.A1(new_n776_), .A2(new_n777_), .B1(KEYINPUT117), .B2(KEYINPUT54), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT57), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n579_), .A2(new_n580_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n583_), .A2(new_n578_), .A3(new_n581_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n780_), .A2(new_n781_), .A3(new_n590_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n592_), .A2(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n783_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n368_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n786_));
  AOI22_X1  g585(.A1(new_n377_), .A2(new_n785_), .B1(new_n786_), .B2(new_n379_), .ZN(new_n787_));
  OAI21_X1  g586(.A(KEYINPUT119), .B1(new_n377_), .B2(new_n785_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n376_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n373_), .A2(KEYINPUT69), .A3(new_n374_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  OR2_X1    g590(.A1(new_n370_), .A2(new_n371_), .ZN(new_n792_));
  AOI22_X1  g591(.A1(new_n792_), .A2(new_n369_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT119), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n791_), .A2(new_n793_), .A3(new_n794_), .A4(KEYINPUT55), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n787_), .A2(new_n788_), .A3(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(new_n385_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT56), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT120), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT56), .B1(new_n796_), .B2(new_n385_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT120), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n796_), .A2(KEYINPUT56), .A3(new_n385_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT121), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n796_), .A2(KEYINPUT121), .A3(KEYINPUT56), .A4(new_n385_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n801_), .A2(new_n803_), .A3(new_n806_), .A4(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n391_), .A2(new_n593_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT118), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n809_), .B(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n784_), .B1(new_n808_), .B2(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n779_), .B1(new_n813_), .B2(new_n629_), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n806_), .A2(new_n807_), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT120), .B1(new_n797_), .B2(new_n798_), .ZN(new_n816_));
  AOI211_X1 g615(.A(new_n800_), .B(KEYINPUT56), .C1(new_n796_), .C2(new_n385_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n811_), .B1(new_n815_), .B2(new_n818_), .ZN(new_n819_));
  OAI211_X1 g618(.A(KEYINPUT57), .B(new_n294_), .C1(new_n819_), .C2(new_n784_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n387_), .A2(new_n783_), .ZN(new_n821_));
  AND3_X1   g620(.A1(new_n796_), .A2(KEYINPUT56), .A3(new_n385_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n821_), .B1(new_n822_), .B2(new_n802_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT58), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n299_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n799_), .A2(new_n804_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n826_), .A2(KEYINPUT122), .A3(KEYINPUT58), .A4(new_n821_), .ZN(new_n827_));
  OAI211_X1 g626(.A(KEYINPUT58), .B(new_n821_), .C1(new_n822_), .C2(new_n802_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT122), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n825_), .A2(new_n827_), .A3(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n814_), .A2(new_n820_), .A3(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n778_), .B1(new_n832_), .B2(new_n361_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n632_), .A2(new_n695_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n834_), .A2(new_n536_), .A3(new_n550_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n833_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(G113gat), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n836_), .A2(new_n837_), .A3(new_n593_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT59), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n839_), .B1(new_n833_), .B2(new_n835_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n835_), .ZN(new_n841_));
  AND3_X1   g640(.A1(new_n825_), .A2(new_n827_), .A3(new_n830_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n294_), .B1(new_n819_), .B2(new_n784_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(new_n779_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n362_), .B1(new_n844_), .B2(new_n820_), .ZN(new_n845_));
  OAI211_X1 g644(.A(KEYINPUT59), .B(new_n841_), .C1(new_n845_), .C2(new_n778_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n594_), .B1(new_n840_), .B2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n838_), .B1(new_n847_), .B2(new_n837_), .ZN(G1340gat));
  INV_X1    g647(.A(G120gat), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(new_n393_), .B2(KEYINPUT60), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n836_), .B(new_n850_), .C1(KEYINPUT60), .C2(new_n849_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n393_), .B1(new_n840_), .B2(new_n846_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT123), .ZN(new_n853_));
  OAI21_X1  g652(.A(G120gat), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  AOI211_X1 g653(.A(KEYINPUT123), .B(new_n393_), .C1(new_n840_), .C2(new_n846_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n851_), .B1(new_n854_), .B2(new_n855_), .ZN(G1341gat));
  AOI21_X1  g655(.A(G127gat), .B1(new_n836_), .B2(new_n362_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n840_), .A2(new_n846_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n361_), .A2(KEYINPUT124), .ZN(new_n859_));
  MUX2_X1   g658(.A(KEYINPUT124), .B(new_n859_), .S(G127gat), .Z(new_n860_));
  AOI21_X1  g659(.A(new_n857_), .B1(new_n858_), .B2(new_n860_), .ZN(G1342gat));
  INV_X1    g660(.A(G134gat), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n836_), .A2(new_n862_), .A3(new_n629_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n299_), .B1(new_n840_), .B2(new_n846_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n864_), .B2(new_n862_), .ZN(G1343gat));
  NOR4_X1   g664(.A1(new_n632_), .A2(new_n515_), .A3(new_n537_), .A4(new_n550_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n833_), .A2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n593_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g669(.A1(new_n868_), .A2(new_n701_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g671(.A(KEYINPUT125), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n868_), .A2(new_n873_), .A3(new_n362_), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n362_), .B(new_n866_), .C1(new_n845_), .C2(new_n778_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(KEYINPUT125), .ZN(new_n876_));
  XNOR2_X1  g675(.A(KEYINPUT61), .B(G155gat), .ZN(new_n877_));
  AND3_X1   g676(.A1(new_n874_), .A2(new_n876_), .A3(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n877_), .B1(new_n874_), .B2(new_n876_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1346gat));
  INV_X1    g679(.A(new_n868_), .ZN(new_n881_));
  OR3_X1    g680(.A1(new_n881_), .A2(G162gat), .A3(new_n294_), .ZN(new_n882_));
  OAI21_X1  g681(.A(G162gat), .B1(new_n881_), .B2(new_n299_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(G1347gat));
  INV_X1    g683(.A(KEYINPUT62), .ZN(new_n885_));
  INV_X1    g684(.A(new_n593_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n608_), .A2(new_n695_), .A3(new_n536_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  NOR4_X1   g687(.A1(new_n833_), .A2(new_n472_), .A3(new_n886_), .A4(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT22), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n885_), .B1(new_n889_), .B2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(G169gat), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n413_), .B1(new_n889_), .B2(new_n885_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n891_), .B2(new_n893_), .ZN(G1348gat));
  NOR2_X1   g693(.A1(new_n833_), .A2(new_n472_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n887_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n896_), .A2(new_n393_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(new_n414_), .ZN(G1349gat));
  NAND3_X1  g697(.A1(new_n895_), .A2(new_n362_), .A3(new_n887_), .ZN(new_n899_));
  MUX2_X1   g698(.A(new_n410_), .B(G183gat), .S(new_n899_), .Z(G1350gat));
  OAI21_X1  g699(.A(G190gat), .B1(new_n896_), .B2(new_n299_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n629_), .A2(new_n411_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n896_), .B2(new_n902_), .ZN(G1351gat));
  NAND2_X1  g702(.A1(new_n608_), .A2(new_n552_), .ZN(new_n904_));
  NOR3_X1   g703(.A1(new_n833_), .A2(new_n472_), .A3(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(new_n593_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(KEYINPUT126), .B(G197gat), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n906_), .B(new_n907_), .ZN(G1352gat));
  NAND2_X1  g707(.A1(new_n905_), .A2(new_n701_), .ZN(new_n909_));
  MUX2_X1   g708(.A(new_n428_), .B(G204gat), .S(new_n909_), .Z(G1353gat));
  INV_X1    g709(.A(new_n904_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(KEYINPUT63), .B(G211gat), .ZN(new_n912_));
  NAND4_X1  g711(.A1(new_n895_), .A2(new_n362_), .A3(new_n911_), .A4(new_n912_), .ZN(new_n913_));
  NOR4_X1   g712(.A1(new_n833_), .A2(new_n361_), .A3(new_n472_), .A4(new_n904_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n913_), .B1(new_n914_), .B2(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(KEYINPUT127), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT127), .ZN(new_n918_));
  OAI211_X1 g717(.A(new_n913_), .B(new_n918_), .C1(new_n914_), .C2(new_n915_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n917_), .A2(new_n919_), .ZN(G1354gat));
  INV_X1    g719(.A(G218gat), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n905_), .A2(new_n921_), .A3(new_n629_), .ZN(new_n922_));
  AND2_X1   g721(.A1(new_n905_), .A2(new_n657_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n922_), .B1(new_n923_), .B2(new_n921_), .ZN(G1355gat));
endmodule


