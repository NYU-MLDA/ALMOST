//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 1 1 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 0 0 1 1 1 0 1 0 0 0 1 1 0 1 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n765_, new_n766_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n891_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n917_, new_n919_, new_n920_, new_n921_, new_n923_, new_n924_,
    new_n926_, new_n927_, new_n928_, new_n930_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_;
  INV_X1    g000(.A(KEYINPUT85), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G227gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT83), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT84), .ZN(new_n205_));
  OR2_X1    g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G71gat), .B(G99gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n204_), .A2(new_n205_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n206_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n207_), .B1(new_n206_), .B2(new_n208_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT22), .B(G169gat), .ZN(new_n215_));
  INV_X1    g014(.A(G176gat), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n214_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G183gat), .A2(G190gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT23), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  OR2_X1    g019(.A1(G183gat), .A2(G190gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n220_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n217_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT26), .B(G190gat), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT82), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT25), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n226_), .B1(new_n227_), .B2(G183gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT25), .B(G183gat), .ZN(new_n229_));
  OAI211_X1 g028(.A(new_n225_), .B(new_n228_), .C1(new_n229_), .C2(new_n226_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n218_), .B(KEYINPUT23), .ZN(new_n232_));
  OR2_X1    g031(.A1(G169gat), .A2(G176gat), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n233_), .A2(KEYINPUT24), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n233_), .A2(KEYINPUT24), .A3(new_n213_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n232_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n224_), .B1(new_n231_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT30), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n237_), .A2(new_n238_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n212_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G15gat), .B(G43gat), .ZN(new_n243_));
  AND3_X1   g042(.A1(new_n232_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n244_));
  AOI22_X1  g043(.A1(new_n244_), .A2(new_n230_), .B1(new_n217_), .B2(new_n223_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT30), .ZN(new_n246_));
  OAI211_X1 g045(.A(new_n246_), .B(new_n239_), .C1(new_n210_), .C2(new_n211_), .ZN(new_n247_));
  AND3_X1   g046(.A1(new_n242_), .A2(new_n243_), .A3(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n243_), .B1(new_n242_), .B2(new_n247_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n202_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n242_), .A2(new_n247_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n243_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n242_), .A2(new_n247_), .A3(new_n243_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n253_), .A2(KEYINPUT85), .A3(new_n254_), .ZN(new_n255_));
  XOR2_X1   g054(.A(G127gat), .B(G134gat), .Z(new_n256_));
  XOR2_X1   g055(.A(G113gat), .B(G120gat), .Z(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT31), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n250_), .A2(new_n255_), .A3(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n259_), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n253_), .A2(KEYINPUT85), .A3(new_n254_), .A4(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  XOR2_X1   g062(.A(G155gat), .B(G162gat), .Z(new_n264_));
  INV_X1    g063(.A(KEYINPUT1), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n267_));
  NOR2_X1   g066(.A1(G141gat), .A2(G148gat), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G141gat), .A2(G148gat), .ZN(new_n270_));
  AND2_X1   g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n266_), .A2(KEYINPUT86), .A3(new_n267_), .A4(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT86), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G155gat), .B(G162gat), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n274_), .A2(KEYINPUT1), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n269_), .A2(new_n267_), .A3(new_n270_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n273_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n268_), .B(KEYINPUT3), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n270_), .B(KEYINPUT2), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  AOI22_X1  g079(.A1(new_n272_), .A2(new_n277_), .B1(new_n264_), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT29), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  XOR2_X1   g082(.A(G22gat), .B(G50gat), .Z(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT28), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n283_), .B(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G78gat), .B(G106gat), .ZN(new_n287_));
  XOR2_X1   g086(.A(new_n287_), .B(KEYINPUT92), .Z(new_n288_));
  XNOR2_X1  g087(.A(G211gat), .B(G218gat), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  XOR2_X1   g089(.A(KEYINPUT88), .B(G197gat), .Z(new_n291_));
  INV_X1    g090(.A(G204gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT21), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n294_), .B1(G197gat), .B2(G204gat), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n290_), .B1(new_n293_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT89), .ZN(new_n297_));
  NOR2_X1   g096(.A1(G197gat), .A2(G204gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT88), .B(G197gat), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n298_), .B1(new_n299_), .B2(G204gat), .ZN(new_n300_));
  OAI211_X1 g099(.A(new_n296_), .B(new_n297_), .C1(KEYINPUT21), .C2(new_n300_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n299_), .A2(G204gat), .ZN(new_n302_));
  INV_X1    g101(.A(new_n295_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n289_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n300_), .A2(KEYINPUT21), .ZN(new_n305_));
  OAI21_X1  g104(.A(KEYINPUT89), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n301_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT90), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n289_), .B(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n300_), .ZN(new_n310_));
  NOR3_X1   g109(.A1(new_n309_), .A2(new_n310_), .A3(new_n294_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n307_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n272_), .A2(new_n277_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n280_), .A2(new_n264_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT29), .ZN(new_n317_));
  INV_X1    g116(.A(G233gat), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT87), .ZN(new_n319_));
  OR2_X1    g118(.A1(new_n319_), .A2(G228gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(G228gat), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n318_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  XOR2_X1   g121(.A(new_n322_), .B(KEYINPUT91), .Z(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n313_), .A2(new_n317_), .A3(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n311_), .B1(new_n301_), .B2(new_n306_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n281_), .A2(new_n282_), .ZN(new_n327_));
  OAI22_X1  g126(.A1(new_n326_), .A2(new_n327_), .B1(KEYINPUT91), .B2(new_n322_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n288_), .B1(new_n325_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT93), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n286_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT94), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n325_), .A2(new_n328_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n288_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n335_), .A2(new_n329_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT94), .ZN(new_n337_));
  OAI211_X1 g136(.A(new_n337_), .B(new_n286_), .C1(new_n329_), .C2(new_n330_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n332_), .A2(new_n336_), .A3(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n336_), .B1(new_n332_), .B2(new_n338_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n263_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  OR2_X1    g141(.A1(new_n335_), .A2(new_n329_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n322_), .A2(KEYINPUT91), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n344_), .B1(new_n313_), .B2(new_n317_), .ZN(new_n345_));
  NOR3_X1   g144(.A1(new_n326_), .A2(new_n327_), .A3(new_n323_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n334_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT93), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n337_), .B1(new_n348_), .B2(new_n286_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n338_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n343_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  AND2_X1   g150(.A1(new_n260_), .A2(new_n262_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n351_), .A2(new_n352_), .A3(new_n339_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n342_), .A2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT20), .B1(new_n326_), .B2(new_n245_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G226gat), .A2(G233gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT19), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT98), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n236_), .B1(new_n229_), .B2(new_n225_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n232_), .A2(new_n221_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT96), .ZN(new_n363_));
  AND2_X1   g162(.A1(new_n363_), .A2(new_n217_), .ZN(new_n364_));
  OR2_X1    g163(.A1(new_n362_), .A2(KEYINPUT96), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n361_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  AND3_X1   g165(.A1(new_n326_), .A2(new_n360_), .A3(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n360_), .B1(new_n326_), .B2(new_n366_), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n356_), .B(new_n359_), .C1(new_n367_), .C2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n307_), .A2(new_n312_), .A3(new_n245_), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n370_), .B(KEYINPUT20), .C1(new_n326_), .C2(new_n366_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n358_), .B(KEYINPUT95), .ZN(new_n372_));
  AND3_X1   g171(.A1(new_n371_), .A2(KEYINPUT97), .A3(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(KEYINPUT97), .B1(new_n371_), .B2(new_n372_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n369_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G8gat), .B(G36gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT18), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(G64gat), .ZN(new_n378_));
  INV_X1    g177(.A(G92gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n375_), .A2(new_n381_), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n369_), .B(new_n380_), .C1(new_n373_), .C2(new_n374_), .ZN(new_n383_));
  AOI21_X1  g182(.A(KEYINPUT27), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G225gat), .A2(G233gat), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT4), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT100), .ZN(new_n388_));
  INV_X1    g187(.A(new_n258_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n388_), .B1(new_n316_), .B2(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n281_), .A2(KEYINPUT100), .A3(new_n258_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n316_), .A2(KEYINPUT99), .A3(new_n389_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT99), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n394_), .B1(new_n281_), .B2(new_n258_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n387_), .B1(new_n392_), .B2(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(KEYINPUT4), .B1(new_n316_), .B2(new_n389_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n386_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  AND2_X1   g198(.A1(new_n392_), .A2(new_n396_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(new_n385_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G1gat), .B(G29gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(KEYINPUT0), .ZN(new_n404_));
  INV_X1    g203(.A(G57gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(G85gat), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n402_), .A2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n399_), .A2(new_n401_), .A3(new_n407_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT27), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n326_), .A2(new_n366_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n358_), .B1(new_n413_), .B2(new_n355_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n414_), .B1(new_n372_), .B2(new_n371_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n412_), .B1(new_n415_), .B2(new_n381_), .ZN(new_n416_));
  AND2_X1   g215(.A1(new_n416_), .A2(new_n383_), .ZN(new_n417_));
  NOR3_X1   g216(.A1(new_n384_), .A2(new_n411_), .A3(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n380_), .A2(KEYINPUT32), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT102), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n421_), .B(new_n369_), .C1(new_n374_), .C2(new_n373_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n415_), .A2(KEYINPUT32), .A3(new_n380_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n411_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT33), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n402_), .A2(new_n425_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n399_), .A2(KEYINPUT33), .A3(new_n401_), .A4(new_n407_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n382_), .A2(new_n426_), .A3(new_n383_), .A4(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n385_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT101), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT101), .ZN(new_n431_));
  OAI211_X1 g230(.A(new_n431_), .B(new_n385_), .C1(new_n397_), .C2(new_n398_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n400_), .A2(new_n386_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n430_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n407_), .B1(new_n434_), .B2(KEYINPUT33), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n424_), .B1(new_n428_), .B2(new_n435_), .ZN(new_n436_));
  NOR3_X1   g235(.A1(new_n340_), .A2(new_n352_), .A3(new_n341_), .ZN(new_n437_));
  AOI22_X1  g236(.A1(new_n354_), .A2(new_n418_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(G64gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(G57gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n405_), .A2(G64gat), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n440_), .A2(new_n441_), .A3(KEYINPUT11), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT67), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G57gat), .B(G64gat), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT67), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n444_), .A2(new_n445_), .A3(KEYINPUT11), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n440_), .A2(new_n441_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT11), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  XOR2_X1   g248(.A(G71gat), .B(G78gat), .Z(new_n450_));
  AND4_X1   g249(.A1(new_n443_), .A2(new_n446_), .A3(new_n449_), .A4(new_n450_), .ZN(new_n451_));
  AOI22_X1  g250(.A1(new_n443_), .A2(new_n446_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT12), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT7), .ZN(new_n454_));
  INV_X1    g253(.A(G99gat), .ZN(new_n455_));
  INV_X1    g254(.A(G106gat), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n454_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G99gat), .A2(G106gat), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT6), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n457_), .A2(new_n460_), .A3(new_n461_), .A4(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(G85gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(new_n379_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G85gat), .A2(G92gat), .ZN(new_n466_));
  AND2_X1   g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n463_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(KEYINPUT8), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT8), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n463_), .A2(new_n470_), .A3(new_n467_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT65), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND4_X1  g273(.A1(KEYINPUT65), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  OR2_X1    g275(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n477_));
  NAND2_X1  g276(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n477_), .A2(new_n466_), .A3(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n476_), .A2(new_n465_), .A3(new_n479_), .ZN(new_n480_));
  AND2_X1   g279(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n481_));
  NOR2_X1   g280(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n482_));
  NOR3_X1   g281(.A1(new_n481_), .A2(new_n482_), .A3(G106gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n460_), .A2(new_n461_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  AOI22_X1  g284(.A1(new_n469_), .A2(new_n471_), .B1(new_n480_), .B2(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT68), .B1(new_n453_), .B2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT12), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n450_), .B1(KEYINPUT11), .B2(new_n444_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n445_), .B1(new_n444_), .B2(KEYINPUT11), .ZN(new_n490_));
  AND4_X1   g289(.A1(new_n445_), .A2(new_n440_), .A3(new_n441_), .A4(KEYINPUT11), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n489_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n443_), .A2(new_n446_), .A3(new_n449_), .A4(new_n450_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n488_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT68), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n480_), .A2(new_n485_), .ZN(new_n496_));
  AND3_X1   g295(.A1(new_n463_), .A2(new_n470_), .A3(new_n467_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n470_), .B1(new_n463_), .B2(new_n467_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n496_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n494_), .A2(new_n495_), .A3(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n487_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(KEYINPUT66), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n451_), .A2(new_n452_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT66), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n496_), .B(new_n504_), .C1(new_n497_), .C2(new_n498_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n502_), .A2(new_n503_), .A3(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n503_), .B1(new_n502_), .B2(new_n505_), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n501_), .B(new_n506_), .C1(KEYINPUT12), .C2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G230gat), .A2(G233gat), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT69), .B1(new_n508_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n507_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(new_n506_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(new_n510_), .ZN(new_n514_));
  AND3_X1   g313(.A1(new_n494_), .A2(new_n495_), .A3(new_n499_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n495_), .B1(new_n494_), .B2(new_n499_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n506_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n502_), .A2(new_n505_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n503_), .ZN(new_n520_));
  AOI21_X1  g319(.A(KEYINPUT12), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT69), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n518_), .A2(new_n522_), .A3(new_n523_), .A4(new_n509_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n511_), .A2(new_n514_), .A3(new_n524_), .ZN(new_n525_));
  XOR2_X1   g324(.A(KEYINPUT70), .B(KEYINPUT5), .Z(new_n526_));
  XNOR2_X1  g325(.A(G120gat), .B(G148gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G176gat), .B(G204gat), .ZN(new_n529_));
  XOR2_X1   g328(.A(new_n528_), .B(new_n529_), .Z(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n525_), .A2(new_n531_), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n511_), .A2(new_n514_), .A3(new_n524_), .A4(new_n530_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n534_), .B1(KEYINPUT71), .B2(KEYINPUT13), .ZN(new_n535_));
  XOR2_X1   g334(.A(KEYINPUT71), .B(KEYINPUT13), .Z(new_n536_));
  AOI21_X1  g335(.A(new_n536_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n535_), .A2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G113gat), .B(G141gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(G197gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(KEYINPUT80), .B(G169gat), .ZN(new_n541_));
  XOR2_X1   g340(.A(new_n540_), .B(new_n541_), .Z(new_n542_));
  XNOR2_X1  g341(.A(G15gat), .B(G22gat), .ZN(new_n543_));
  INV_X1    g342(.A(G1gat), .ZN(new_n544_));
  INV_X1    g343(.A(G8gat), .ZN(new_n545_));
  OAI21_X1  g344(.A(KEYINPUT14), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n543_), .A2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G1gat), .B(G8gat), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n547_), .B(new_n548_), .Z(new_n549_));
  XNOR2_X1  g348(.A(G29gat), .B(G36gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G43gat), .B(G50gat), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n551_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n549_), .A2(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n547_), .B(new_n548_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n556_), .A2(new_n553_), .A3(new_n552_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT79), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G229gat), .A2(G233gat), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n559_), .A2(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n554_), .B(KEYINPUT15), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(new_n556_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n564_), .A2(new_n560_), .A3(new_n555_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n542_), .B1(new_n562_), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n562_), .A2(new_n565_), .A3(new_n542_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n567_), .A2(KEYINPUT81), .A3(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT81), .ZN(new_n570_));
  AND3_X1   g369(.A1(new_n562_), .A2(new_n565_), .A3(new_n542_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n570_), .B1(new_n571_), .B2(new_n566_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n569_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NOR3_X1   g373(.A1(new_n438_), .A2(new_n538_), .A3(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G232gat), .A2(G233gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT34), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT35), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n502_), .A2(new_n554_), .A3(new_n505_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n578_), .A2(new_n579_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n581_), .A2(KEYINPUT73), .A3(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n563_), .A2(KEYINPUT72), .A3(new_n499_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n563_), .A2(new_n499_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT72), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n583_), .A2(new_n584_), .A3(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(KEYINPUT73), .B1(new_n581_), .B2(new_n582_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n580_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n580_), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n581_), .A2(new_n585_), .A3(new_n591_), .A4(new_n582_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n590_), .A2(new_n592_), .ZN(new_n593_));
  XOR2_X1   g392(.A(G134gat), .B(G162gat), .Z(new_n594_));
  XNOR2_X1  g393(.A(G190gat), .B(G218gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT36), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n596_), .A2(new_n597_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n593_), .A2(new_n598_), .A3(new_n600_), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n590_), .A2(new_n597_), .A3(new_n596_), .A4(new_n592_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(KEYINPUT74), .B(KEYINPUT37), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  AND3_X1   g403(.A1(new_n601_), .A2(new_n602_), .A3(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n604_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G183gat), .B(G211gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G127gat), .B(G155gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n612_), .A2(KEYINPUT17), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n612_), .A2(KEYINPUT17), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT75), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n556_), .B(new_n616_), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n617_), .A2(new_n520_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(G231gat), .A2(G233gat), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n617_), .A2(new_n520_), .ZN(new_n621_));
  AND3_X1   g420(.A1(new_n618_), .A2(new_n620_), .A3(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n620_), .B1(new_n618_), .B2(new_n621_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n615_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n624_), .A2(KEYINPUT77), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n622_), .A2(new_n623_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(new_n613_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n624_), .A2(KEYINPUT77), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n625_), .A2(new_n627_), .A3(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n607_), .A2(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT78), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n575_), .A2(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n632_), .A2(new_n544_), .A3(new_n411_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT38), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n535_), .A2(new_n537_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n567_), .A2(new_n568_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n636_), .A2(new_n629_), .A3(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n601_), .A2(new_n602_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n638_), .A2(new_n640_), .A3(new_n438_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n544_), .B1(new_n641_), .B2(new_n411_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n635_), .A2(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n643_), .B1(new_n634_), .B2(new_n633_), .ZN(G1324gat));
  INV_X1    g443(.A(KEYINPUT40), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n384_), .A2(new_n417_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n641_), .A2(new_n647_), .ZN(new_n648_));
  OR2_X1    g447(.A1(new_n648_), .A2(KEYINPUT103), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n545_), .B1(new_n648_), .B2(KEYINPUT103), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT39), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(KEYINPUT104), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n651_), .A2(KEYINPUT104), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n649_), .A2(new_n650_), .A3(new_n652_), .A4(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n632_), .A2(new_n545_), .A3(new_n647_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n652_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n645_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n657_), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n659_), .A2(KEYINPUT40), .A3(new_n655_), .A4(new_n654_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(G1325gat));
  INV_X1    g460(.A(G15gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n662_), .B1(new_n641_), .B2(new_n352_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT41), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n632_), .A2(new_n662_), .A3(new_n352_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1326gat));
  INV_X1    g465(.A(G22gat), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n340_), .A2(new_n341_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n667_), .B1(new_n641_), .B2(new_n669_), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT42), .Z(new_n671_));
  NAND3_X1  g470(.A1(new_n632_), .A2(new_n667_), .A3(new_n669_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1327gat));
  NOR2_X1   g472(.A1(new_n629_), .A2(new_n639_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n575_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(G29gat), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n411_), .A2(new_n676_), .ZN(new_n677_));
  XOR2_X1   g476(.A(new_n677_), .B(KEYINPUT107), .Z(new_n678_));
  NAND2_X1  g477(.A1(new_n675_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n411_), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n351_), .A2(new_n352_), .A3(new_n339_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n352_), .B1(new_n351_), .B2(new_n339_), .ZN(new_n682_));
  OAI211_X1 g481(.A(new_n646_), .B(new_n680_), .C1(new_n681_), .C2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n436_), .A2(new_n437_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n607_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(KEYINPUT43), .B1(new_n685_), .B2(KEYINPUT105), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT105), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT43), .ZN(new_n688_));
  OAI211_X1 g487(.A(new_n687_), .B(new_n688_), .C1(new_n438_), .C2(new_n607_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n625_), .A2(new_n627_), .A3(new_n628_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n636_), .A2(new_n690_), .A3(new_n637_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n686_), .A2(new_n689_), .A3(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n693_), .A2(new_n694_), .A3(KEYINPUT44), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n680_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n679_), .B1(new_n699_), .B2(new_n676_), .ZN(G1328gat));
  NOR2_X1   g499(.A1(new_n646_), .A2(G36gat), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n575_), .A2(new_n674_), .A3(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(KEYINPUT108), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT108), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n575_), .A2(new_n704_), .A3(new_n674_), .A4(new_n701_), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n703_), .A2(KEYINPUT45), .A3(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(KEYINPUT45), .B1(new_n703_), .B2(new_n705_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n646_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n709_));
  INV_X1    g508(.A(G36gat), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n708_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT46), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n708_), .B(KEYINPUT46), .C1(new_n709_), .C2(new_n710_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(G1329gat));
  NAND2_X1  g514(.A1(new_n352_), .A2(G43gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n716_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n717_));
  XOR2_X1   g516(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n718_));
  XNOR2_X1  g517(.A(KEYINPUT109), .B(G43gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n719_), .B1(new_n675_), .B2(new_n352_), .ZN(new_n720_));
  OR3_X1    g519(.A1(new_n717_), .A2(new_n718_), .A3(new_n720_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n718_), .B1(new_n717_), .B2(new_n720_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1330gat));
  AOI21_X1  g522(.A(G50gat), .B1(new_n675_), .B2(new_n669_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n697_), .A2(new_n698_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n669_), .A2(G50gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n724_), .B1(new_n725_), .B2(new_n726_), .ZN(G1331gat));
  NOR2_X1   g526(.A1(new_n438_), .A2(new_n640_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n574_), .A2(new_n629_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n636_), .A2(new_n729_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n728_), .A2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  OAI21_X1  g531(.A(G57gat), .B1(new_n732_), .B2(new_n680_), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n438_), .A2(new_n636_), .A3(new_n637_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n734_), .A2(new_n631_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n735_), .A2(new_n405_), .A3(new_n411_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n733_), .A2(new_n736_), .ZN(G1332gat));
  AOI21_X1  g536(.A(new_n439_), .B1(new_n731_), .B2(new_n647_), .ZN(new_n738_));
  XOR2_X1   g537(.A(KEYINPUT111), .B(KEYINPUT48), .Z(new_n739_));
  XNOR2_X1  g538(.A(new_n738_), .B(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n735_), .A2(new_n439_), .A3(new_n647_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(G1333gat));
  INV_X1    g541(.A(G71gat), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n735_), .A2(new_n743_), .A3(new_n352_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n731_), .B2(new_n352_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT112), .ZN(new_n746_));
  OR2_X1    g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n746_), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n747_), .A2(KEYINPUT49), .A3(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(KEYINPUT49), .B1(new_n747_), .B2(new_n748_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n744_), .B1(new_n749_), .B2(new_n750_), .ZN(G1334gat));
  INV_X1    g550(.A(G78gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n752_), .B1(new_n731_), .B2(new_n669_), .ZN(new_n753_));
  XOR2_X1   g552(.A(new_n753_), .B(KEYINPUT50), .Z(new_n754_));
  NAND2_X1  g553(.A1(new_n669_), .A2(new_n752_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT113), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n735_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n754_), .A2(new_n757_), .ZN(G1335gat));
  NOR3_X1   g557(.A1(new_n636_), .A2(new_n629_), .A3(new_n637_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n686_), .A2(new_n689_), .A3(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(G85gat), .B1(new_n760_), .B2(new_n680_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n734_), .A2(new_n674_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n762_), .A2(new_n464_), .A3(new_n411_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(G1336gat));
  OAI21_X1  g563(.A(G92gat), .B1(new_n760_), .B2(new_n646_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n762_), .A2(new_n379_), .A3(new_n647_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(G1337gat));
  OAI21_X1  g566(.A(G99gat), .B1(new_n760_), .B2(new_n263_), .ZN(new_n768_));
  NOR3_X1   g567(.A1(new_n263_), .A2(new_n482_), .A3(new_n481_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n762_), .A2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g571(.A1(new_n762_), .A2(new_n456_), .A3(new_n669_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n686_), .A2(new_n669_), .A3(new_n689_), .A4(new_n759_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n774_), .A2(new_n775_), .A3(G106gat), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n774_), .B2(G106gat), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n773_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  XOR2_X1   g577(.A(KEYINPUT114), .B(KEYINPUT53), .Z(new_n779_));
  XNOR2_X1  g578(.A(new_n778_), .B(new_n779_), .ZN(G1339gat));
  NOR2_X1   g579(.A1(new_n647_), .A2(new_n680_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n782_), .A2(new_n353_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n784_));
  INV_X1    g583(.A(new_n607_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n559_), .A2(new_n560_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n560_), .B1(new_n549_), .B2(new_n554_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n542_), .B1(new_n564_), .B2(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n571_), .B1(new_n786_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(new_n533_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT55), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n511_), .A2(new_n791_), .A3(new_n524_), .ZN(new_n792_));
  NOR3_X1   g591(.A1(new_n517_), .A2(new_n521_), .A3(new_n510_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT55), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n510_), .B1(new_n517_), .B2(new_n521_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT116), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT116), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n508_), .A2(new_n797_), .A3(new_n510_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n792_), .A2(new_n794_), .A3(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n531_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT56), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n800_), .A2(KEYINPUT56), .A3(new_n531_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n790_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(KEYINPUT117), .B(KEYINPUT58), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n785_), .B1(new_n805_), .B2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(KEYINPUT118), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n789_), .A2(new_n533_), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT56), .B1(new_n800_), .B2(new_n531_), .ZN(new_n811_));
  AOI22_X1  g610(.A1(new_n796_), .A2(new_n798_), .B1(KEYINPUT55), .B2(new_n793_), .ZN(new_n812_));
  AOI211_X1 g611(.A(new_n802_), .B(new_n530_), .C1(new_n812_), .C2(new_n792_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n810_), .B1(new_n811_), .B2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n607_), .B1(new_n814_), .B2(new_n806_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT118), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n805_), .A2(KEYINPUT58), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n809_), .A2(new_n817_), .A3(new_n818_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n533_), .B(new_n637_), .C1(new_n811_), .C2(new_n813_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n534_), .A2(new_n789_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(KEYINPUT57), .B1(new_n822_), .B2(new_n639_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT57), .ZN(new_n824_));
  AOI211_X1 g623(.A(new_n824_), .B(new_n640_), .C1(new_n820_), .C2(new_n821_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n823_), .A2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n629_), .B1(new_n819_), .B2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT115), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n574_), .A2(new_n629_), .A3(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n729_), .A2(KEYINPUT115), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n636_), .A2(new_n829_), .A3(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(KEYINPUT54), .B1(new_n831_), .B2(new_n785_), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n830_), .A2(new_n829_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT54), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n833_), .A2(new_n834_), .A3(new_n607_), .A4(new_n636_), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n832_), .A2(new_n835_), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n783_), .B(new_n784_), .C1(new_n827_), .C2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT119), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n818_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n839_));
  AOI211_X1 g638(.A(KEYINPUT118), .B(new_n607_), .C1(new_n814_), .C2(new_n806_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n838_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n809_), .A2(KEYINPUT119), .A3(new_n817_), .A4(new_n818_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n841_), .A2(new_n842_), .A3(new_n826_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n836_), .B1(new_n843_), .B2(new_n690_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n783_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT59), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n573_), .B(new_n837_), .C1(new_n846_), .C2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(G113gat), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n637_), .A2(new_n533_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n850_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n821_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n639_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n824_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n822_), .A2(KEYINPUT57), .A3(new_n639_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n856_), .B1(new_n819_), .B2(new_n838_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n629_), .B1(new_n857_), .B2(new_n842_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n783_), .B1(new_n858_), .B2(new_n836_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n637_), .ZN(new_n860_));
  OR3_X1    g659(.A1(new_n859_), .A2(G113gat), .A3(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n849_), .A2(new_n861_), .ZN(G1340gat));
  OAI211_X1 g661(.A(new_n538_), .B(new_n837_), .C1(new_n846_), .C2(new_n847_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(G120gat), .ZN(new_n864_));
  INV_X1    g663(.A(G120gat), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n865_), .A2(KEYINPUT60), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(new_n636_), .B2(KEYINPUT60), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT121), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n866_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n846_), .B(new_n869_), .C1(new_n868_), .C2(new_n867_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n864_), .A2(new_n870_), .ZN(G1341gat));
  OAI211_X1 g670(.A(new_n629_), .B(new_n837_), .C1(new_n846_), .C2(new_n847_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(G127gat), .ZN(new_n873_));
  OR3_X1    g672(.A1(new_n859_), .A2(G127gat), .A3(new_n690_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(G1342gat));
  NOR3_X1   g674(.A1(new_n844_), .A2(new_n639_), .A3(new_n845_), .ZN(new_n876_));
  OAI21_X1  g675(.A(KEYINPUT122), .B1(new_n876_), .B2(G134gat), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT122), .ZN(new_n878_));
  INV_X1    g677(.A(G134gat), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n878_), .B(new_n879_), .C1(new_n859_), .C2(new_n639_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n837_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n881_), .B1(new_n859_), .B2(KEYINPUT59), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n607_), .A2(new_n879_), .ZN(new_n883_));
  AOI22_X1  g682(.A1(new_n877_), .A2(new_n880_), .B1(new_n882_), .B2(new_n883_), .ZN(G1343gat));
  NAND2_X1  g683(.A1(new_n843_), .A2(new_n690_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n836_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n782_), .A2(new_n342_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n887_), .A2(new_n637_), .A3(new_n888_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g689(.A1(new_n887_), .A2(new_n538_), .A3(new_n888_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(G148gat), .ZN(G1345gat));
  NOR3_X1   g691(.A1(new_n844_), .A2(new_n342_), .A3(new_n782_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(KEYINPUT61), .B(G155gat), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(KEYINPUT123), .ZN(new_n895_));
  AND3_X1   g694(.A1(new_n893_), .A2(new_n629_), .A3(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n895_), .B1(new_n893_), .B2(new_n629_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n896_), .A2(new_n897_), .ZN(G1346gat));
  INV_X1    g697(.A(G162gat), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n893_), .A2(new_n899_), .A3(new_n640_), .ZN(new_n900_));
  AND2_X1   g699(.A1(new_n893_), .A2(new_n785_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(new_n899_), .ZN(G1347gat));
  NOR2_X1   g701(.A1(new_n646_), .A2(new_n411_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n352_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(KEYINPUT124), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  OAI211_X1 g705(.A(new_n668_), .B(new_n906_), .C1(new_n827_), .C2(new_n836_), .ZN(new_n907_));
  OAI21_X1  g706(.A(G169gat), .B1(new_n907_), .B2(new_n860_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT62), .ZN(new_n909_));
  OR2_X1    g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n907_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n911_), .A2(new_n215_), .A3(new_n637_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n908_), .A2(new_n909_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n910_), .A2(new_n912_), .A3(new_n913_), .ZN(G1348gat));
  AOI21_X1  g713(.A(G176gat), .B1(new_n911_), .B2(new_n538_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n844_), .A2(new_n669_), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n905_), .A2(new_n216_), .A3(new_n636_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n915_), .B1(new_n916_), .B2(new_n917_), .ZN(G1349gat));
  NOR3_X1   g717(.A1(new_n907_), .A2(new_n690_), .A3(new_n229_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n916_), .A2(new_n629_), .A3(new_n906_), .ZN(new_n920_));
  INV_X1    g719(.A(G183gat), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n919_), .B1(new_n920_), .B2(new_n921_), .ZN(G1350gat));
  OAI21_X1  g721(.A(G190gat), .B1(new_n907_), .B2(new_n607_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n640_), .A2(new_n225_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n923_), .B1(new_n907_), .B2(new_n924_), .ZN(G1351gat));
  NAND2_X1  g724(.A1(new_n903_), .A2(new_n682_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n844_), .A2(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(new_n637_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g728(.A1(new_n927_), .A2(new_n538_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g730(.A(new_n690_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n932_));
  INV_X1    g731(.A(new_n932_), .ZN(new_n933_));
  NOR3_X1   g732(.A1(new_n844_), .A2(new_n926_), .A3(new_n933_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n935_));
  INV_X1    g734(.A(new_n935_), .ZN(new_n936_));
  OAI21_X1  g735(.A(KEYINPUT125), .B1(new_n934_), .B2(new_n936_), .ZN(new_n937_));
  INV_X1    g736(.A(new_n926_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n887_), .A2(new_n938_), .A3(new_n932_), .ZN(new_n939_));
  INV_X1    g738(.A(KEYINPUT125), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n939_), .A2(new_n940_), .A3(new_n935_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n934_), .A2(new_n936_), .ZN(new_n942_));
  AND3_X1   g741(.A1(new_n937_), .A2(new_n941_), .A3(new_n942_), .ZN(G1354gat));
  AND3_X1   g742(.A1(new_n927_), .A2(G218gat), .A3(new_n785_), .ZN(new_n944_));
  NAND3_X1  g743(.A1(new_n887_), .A2(new_n640_), .A3(new_n938_), .ZN(new_n945_));
  AOI21_X1  g744(.A(G218gat), .B1(new_n945_), .B2(KEYINPUT126), .ZN(new_n946_));
  INV_X1    g745(.A(KEYINPUT126), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n927_), .A2(new_n947_), .A3(new_n640_), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n944_), .B1(new_n946_), .B2(new_n948_), .ZN(G1355gat));
endmodule


