//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 0 1 0 0 1 1 1 1 1 0 1 1 1 0 0 0 0 1 0 1 1 0 0 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 0 1 0 1 1 0 1 1 0 1 1 1 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n677_, new_n678_,
    new_n679_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n773_, new_n774_, new_n775_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n874_, new_n875_,
    new_n876_, new_n878_, new_n879_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n900_, new_n902_, new_n903_, new_n904_, new_n905_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_;
  INV_X1    g000(.A(KEYINPUT75), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT13), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NOR2_X1   g003(.A1(KEYINPUT75), .A2(KEYINPUT13), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT71), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT68), .ZN(new_n208_));
  OR2_X1    g007(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n209_), .A2(KEYINPUT64), .A3(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n212_));
  AND2_X1   g011(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n212_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n211_), .A2(new_n215_), .ZN(new_n216_));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G106gat), .Z(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G99gat), .A2(G106gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT6), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT6), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(G99gat), .A3(G106gat), .ZN(new_n222_));
  AND3_X1   g021(.A1(new_n220_), .A2(new_n222_), .A3(KEYINPUT67), .ZN(new_n223_));
  AOI21_X1  g022(.A(KEYINPUT67), .B1(new_n220_), .B2(new_n222_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT66), .ZN(new_n226_));
  OAI211_X1 g025(.A(G85gat), .B(G92gat), .C1(new_n226_), .C2(KEYINPUT9), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n226_), .B(KEYINPUT9), .C1(G85gat), .C2(G92gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n226_), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  AND4_X1   g030(.A1(new_n208_), .A2(new_n218_), .A3(new_n225_), .A4(new_n231_), .ZN(new_n232_));
  AOI22_X1  g031(.A1(new_n216_), .A2(new_n217_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n208_), .B1(new_n233_), .B2(new_n225_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n232_), .A2(new_n234_), .ZN(new_n235_));
  XOR2_X1   g034(.A(G85gat), .B(G92gat), .Z(new_n236_));
  INV_X1    g035(.A(KEYINPUT8), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT69), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(KEYINPUT7), .ZN(new_n240_));
  NOR2_X1   g039(.A1(G99gat), .A2(G106gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(KEYINPUT69), .B(KEYINPUT7), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n242_), .B1(new_n243_), .B2(new_n241_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n238_), .B1(new_n225_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT7), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(KEYINPUT69), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n241_), .B1(new_n240_), .B2(new_n248_), .ZN(new_n249_));
  AOI211_X1 g048(.A(G99gat), .B(G106gat), .C1(new_n239_), .C2(KEYINPUT7), .ZN(new_n250_));
  OAI21_X1  g049(.A(KEYINPUT70), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n220_), .A2(new_n222_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT70), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n253_), .B(new_n242_), .C1(new_n243_), .C2(new_n241_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n251_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(new_n236_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n246_), .B1(new_n256_), .B2(KEYINPUT8), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n207_), .B1(new_n235_), .B2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n246_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n236_), .ZN(new_n260_));
  AOI22_X1  g059(.A1(new_n244_), .A2(KEYINPUT70), .B1(new_n220_), .B2(new_n222_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n260_), .B1(new_n261_), .B2(new_n254_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n259_), .B1(new_n262_), .B2(new_n237_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n218_), .A2(new_n225_), .A3(new_n231_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT68), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n233_), .A2(new_n208_), .A3(new_n225_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n263_), .A2(new_n267_), .A3(KEYINPUT71), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G57gat), .B(G64gat), .ZN(new_n269_));
  OR2_X1    g068(.A1(new_n269_), .A2(KEYINPUT11), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(KEYINPUT11), .ZN(new_n271_));
  XOR2_X1   g070(.A(G71gat), .B(G78gat), .Z(new_n272_));
  NAND3_X1  g071(.A1(new_n270_), .A2(new_n271_), .A3(new_n272_), .ZN(new_n273_));
  OR2_X1    g072(.A1(new_n271_), .A2(new_n272_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT72), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n258_), .A2(new_n268_), .A3(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n263_), .A2(new_n267_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n275_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n278_), .A2(KEYINPUT12), .A3(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n277_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n258_), .A2(new_n268_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n276_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT12), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G230gat), .A2(G233gat), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n282_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT73), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n285_), .A2(new_n290_), .A3(new_n277_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n276_), .B1(new_n258_), .B2(new_n268_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n288_), .B1(new_n292_), .B2(KEYINPUT73), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G120gat), .B(G148gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT5), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G176gat), .B(G204gat), .ZN(new_n297_));
  XOR2_X1   g096(.A(new_n296_), .B(new_n297_), .Z(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n289_), .A2(new_n294_), .A3(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT74), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n289_), .A2(new_n294_), .A3(KEYINPUT74), .A4(new_n299_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n289_), .A2(new_n294_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(new_n298_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n206_), .B1(new_n304_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n204_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n304_), .A2(new_n306_), .A3(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n311_), .B(KEYINPUT76), .Z(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT105), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G228gat), .A2(G233gat), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  OR2_X1    g115(.A1(G141gat), .A2(G148gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT3), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT94), .ZN(new_n319_));
  NAND3_X1  g118(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n320_), .B1(new_n317_), .B2(KEYINPUT3), .ZN(new_n321_));
  AOI21_X1  g120(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n319_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT92), .ZN(new_n325_));
  INV_X1    g124(.A(G155gat), .ZN(new_n326_));
  INV_X1    g125(.A(G162gat), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n325_), .A2(new_n326_), .A3(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(KEYINPUT92), .B1(G155gat), .B2(G162gat), .ZN(new_n329_));
  AND2_X1   g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G155gat), .A2(G162gat), .ZN(new_n331_));
  AND2_X1   g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(KEYINPUT1), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n328_), .A2(new_n333_), .A3(new_n329_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT93), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n328_), .A2(new_n333_), .A3(KEYINPUT93), .A4(new_n329_), .ZN(new_n337_));
  OAI211_X1 g136(.A(new_n336_), .B(new_n337_), .C1(KEYINPUT1), .C2(new_n331_), .ZN(new_n338_));
  XOR2_X1   g137(.A(G141gat), .B(G148gat), .Z(new_n339_));
  AOI22_X1  g138(.A1(new_n324_), .A2(new_n332_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT29), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  XOR2_X1   g141(.A(G197gat), .B(G204gat), .Z(new_n343_));
  XOR2_X1   g142(.A(G211gat), .B(G218gat), .Z(new_n344_));
  NAND3_X1  g143(.A1(new_n343_), .A2(new_n344_), .A3(KEYINPUT21), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT96), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT21), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G197gat), .B(G204gat), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n344_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(G197gat), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n351_), .A2(KEYINPUT95), .A3(G204gat), .ZN(new_n352_));
  OAI211_X1 g151(.A(KEYINPUT21), .B(new_n352_), .C1(new_n343_), .C2(KEYINPUT95), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n347_), .B1(new_n350_), .B2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n350_), .A2(new_n353_), .A3(new_n347_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n346_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n316_), .B1(new_n342_), .B2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n356_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n345_), .B1(new_n359_), .B2(new_n354_), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n360_), .B(new_n315_), .C1(new_n341_), .C2(new_n340_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n358_), .A2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G78gat), .B(G106gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n363_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n358_), .A2(new_n361_), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n364_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n340_), .A2(new_n341_), .ZN(new_n368_));
  XOR2_X1   g167(.A(G22gat), .B(G50gat), .Z(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT28), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n368_), .B(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n365_), .B1(new_n358_), .B2(new_n361_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n371_), .B1(new_n372_), .B2(KEYINPUT97), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n367_), .A2(new_n373_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n364_), .A2(new_n371_), .A3(KEYINPUT97), .A4(new_n366_), .ZN(new_n375_));
  AND2_X1   g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G1gat), .B(G29gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(G85gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(KEYINPUT0), .B(G57gat), .ZN(new_n379_));
  XOR2_X1   g178(.A(new_n378_), .B(new_n379_), .Z(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n324_), .A2(new_n332_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n338_), .A2(new_n339_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G127gat), .B(G134gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G113gat), .B(G120gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT89), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  OR2_X1    g188(.A1(new_n385_), .A2(new_n386_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT90), .ZN(new_n391_));
  OR2_X1    g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n390_), .A2(new_n391_), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n389_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n384_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G225gat), .A2(G233gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n390_), .A2(new_n387_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n340_), .A2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n395_), .A2(new_n396_), .A3(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT101), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT101), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n395_), .A2(new_n398_), .A3(new_n401_), .A4(new_n396_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n389_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n340_), .A2(new_n404_), .ZN(new_n405_));
  AND3_X1   g204(.A1(new_n382_), .A2(new_n383_), .A3(new_n397_), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT4), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT4), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n395_), .A2(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n396_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n381_), .B1(new_n403_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n396_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n408_), .B1(new_n395_), .B2(new_n398_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n405_), .A2(KEYINPUT4), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n412_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n415_), .A2(new_n380_), .A3(new_n400_), .A4(new_n402_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT102), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n411_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n417_), .B1(new_n411_), .B2(new_n416_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n376_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G226gat), .A2(G233gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(KEYINPUT19), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G183gat), .A2(G190gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(KEYINPUT23), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT23), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n427_), .A2(G183gat), .A3(G190gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n426_), .A2(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(G183gat), .A2(G190gat), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n429_), .A2(new_n431_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(G169gat), .ZN(new_n434_));
  AND2_X1   g233(.A1(new_n432_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  OR3_X1    g235(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n437_));
  AOI21_X1  g236(.A(KEYINPUT87), .B1(new_n426_), .B2(new_n428_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT87), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n439_), .B1(new_n425_), .B2(KEYINPUT23), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n437_), .B1(new_n438_), .B2(new_n440_), .ZN(new_n441_));
  OR2_X1    g240(.A1(new_n441_), .A2(KEYINPUT98), .ZN(new_n442_));
  XNOR2_X1  g241(.A(KEYINPUT26), .B(G190gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(KEYINPUT25), .B(G183gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT24), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n446_), .B1(G169gat), .B2(G176gat), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n447_), .B1(G169gat), .B2(G176gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n445_), .A2(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n449_), .B1(new_n441_), .B2(KEYINPUT98), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n442_), .A2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n357_), .A2(new_n436_), .A3(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT20), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n431_), .B1(new_n438_), .B2(new_n440_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(new_n434_), .ZN(new_n455_));
  INV_X1    g254(.A(G190gat), .ZN(new_n456_));
  OAI21_X1  g255(.A(KEYINPUT86), .B1(new_n456_), .B2(KEYINPUT26), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n457_), .B(new_n444_), .C1(new_n443_), .C2(KEYINPUT86), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n458_), .A2(new_n429_), .A3(new_n448_), .A4(new_n437_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n455_), .A2(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n453_), .B1(new_n360_), .B2(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n424_), .B1(new_n452_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n460_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n453_), .B1(new_n357_), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT99), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n466_), .B1(new_n442_), .B2(new_n450_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n442_), .A2(new_n450_), .A3(new_n466_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n435_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n465_), .B1(new_n470_), .B2(new_n357_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n463_), .B1(new_n471_), .B2(new_n423_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT104), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G8gat), .B(G36gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT18), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G64gat), .B(G92gat), .ZN(new_n476_));
  XOR2_X1   g275(.A(new_n475_), .B(new_n476_), .Z(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT103), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n472_), .A2(new_n473_), .A3(new_n479_), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT20), .B1(new_n360_), .B2(new_n460_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n469_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n436_), .B1(new_n482_), .B2(new_n467_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n481_), .B1(new_n483_), .B2(new_n360_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n462_), .B1(new_n484_), .B2(new_n424_), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT104), .B1(new_n485_), .B2(new_n478_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT100), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n482_), .A2(new_n467_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n357_), .A2(new_n436_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n487_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n360_), .A2(new_n435_), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n491_), .B(KEYINPUT100), .C1(new_n467_), .C2(new_n482_), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n490_), .A2(new_n492_), .A3(new_n424_), .A4(new_n461_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n471_), .A2(new_n423_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n493_), .A2(new_n494_), .A3(new_n477_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n480_), .A2(new_n486_), .A3(KEYINPUT27), .A4(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT27), .ZN(new_n497_));
  AND3_X1   g296(.A1(new_n493_), .A2(new_n494_), .A3(new_n477_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n477_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n497_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n496_), .A2(new_n500_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n314_), .B1(new_n421_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n374_), .A2(new_n375_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n420_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n503_), .B1(new_n504_), .B2(new_n418_), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n505_), .A2(KEYINPUT105), .A3(new_n500_), .A4(new_n496_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT33), .ZN(new_n507_));
  OR2_X1    g306(.A1(new_n416_), .A2(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n412_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n395_), .A2(new_n412_), .A3(new_n398_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(new_n381_), .ZN(new_n511_));
  OAI21_X1  g310(.A(KEYINPUT33), .B1(new_n509_), .B2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(new_n416_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n493_), .A2(new_n494_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n477_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n508_), .A2(new_n513_), .A3(new_n516_), .A4(new_n495_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n411_), .A2(new_n416_), .ZN(new_n518_));
  AND2_X1   g317(.A1(new_n477_), .A2(KEYINPUT32), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n472_), .A2(new_n519_), .ZN(new_n520_));
  OAI211_X1 g319(.A(new_n518_), .B(new_n520_), .C1(new_n514_), .C2(new_n519_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n517_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(new_n503_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n502_), .A2(new_n506_), .A3(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n394_), .B(KEYINPUT31), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT91), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n460_), .B(KEYINPUT30), .ZN(new_n528_));
  XNOR2_X1  g327(.A(KEYINPUT88), .B(G43gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G227gat), .A2(G233gat), .ZN(new_n531_));
  XOR2_X1   g330(.A(new_n531_), .B(G15gat), .Z(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(G71gat), .ZN(new_n533_));
  INV_X1    g332(.A(G99gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n530_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n529_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n528_), .B(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(new_n535_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n527_), .B1(new_n537_), .B2(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n525_), .A2(new_n526_), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n537_), .A2(new_n540_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n541_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n524_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT107), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n496_), .A2(new_n500_), .A3(new_n503_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT106), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT106), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n496_), .A2(new_n500_), .A3(new_n550_), .A4(new_n503_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n549_), .A2(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n544_), .B1(new_n420_), .B2(new_n419_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n547_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n555_));
  AOI211_X1 g354(.A(KEYINPUT107), .B(new_n553_), .C1(new_n549_), .C2(new_n551_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n546_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G29gat), .B(G36gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT78), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G43gat), .B(G50gat), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n559_), .A2(new_n561_), .ZN(new_n562_));
  OR2_X1    g361(.A1(new_n558_), .A2(KEYINPUT78), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n558_), .A2(KEYINPUT78), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n563_), .A2(new_n564_), .A3(new_n560_), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n562_), .A2(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT15), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G15gat), .B(G22gat), .ZN(new_n568_));
  INV_X1    g367(.A(G1gat), .ZN(new_n569_));
  INV_X1    g368(.A(G8gat), .ZN(new_n570_));
  OAI21_X1  g369(.A(KEYINPUT14), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n568_), .A2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G1gat), .B(G8gat), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n572_), .B(new_n573_), .Z(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n567_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n566_), .A2(new_n574_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G229gat), .A2(G233gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT83), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n576_), .A2(new_n577_), .A3(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT84), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT82), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n562_), .A2(new_n565_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n575_), .A2(new_n583_), .ZN(new_n584_));
  AND3_X1   g383(.A1(new_n577_), .A2(new_n582_), .A3(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n582_), .B1(new_n577_), .B2(new_n584_), .ZN(new_n586_));
  OAI211_X1 g385(.A(G229gat), .B(G233gat), .C1(new_n585_), .C2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n580_), .A2(new_n581_), .A3(new_n587_), .ZN(new_n588_));
  XOR2_X1   g387(.A(G113gat), .B(G141gat), .Z(new_n589_));
  XNOR2_X1  g388(.A(G169gat), .B(G197gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n580_), .A2(new_n587_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n591_), .B1(new_n592_), .B2(KEYINPUT84), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n580_), .A2(new_n587_), .A3(new_n591_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT85), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n580_), .A2(new_n587_), .A3(KEYINPUT85), .A4(new_n591_), .ZN(new_n597_));
  AOI22_X1  g396(.A1(new_n588_), .A2(new_n593_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n557_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT79), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n601_), .B1(new_n283_), .B2(new_n583_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n567_), .A2(new_n278_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT80), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n258_), .A2(new_n268_), .A3(KEYINPUT79), .A4(new_n566_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(G232gat), .A2(G233gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT35), .ZN(new_n608_));
  XOR2_X1   g407(.A(KEYINPUT77), .B(KEYINPUT34), .Z(new_n609_));
  XOR2_X1   g408(.A(new_n608_), .B(new_n609_), .Z(new_n610_));
  NAND4_X1  g409(.A1(new_n604_), .A2(new_n605_), .A3(new_n606_), .A4(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n602_), .A2(new_n606_), .A3(new_n603_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT35), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G190gat), .B(G218gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G134gat), .B(G162gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  AOI22_X1  g415(.A1(new_n612_), .A2(new_n613_), .B1(KEYINPUT36), .B2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n610_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n618_), .B1(new_n612_), .B2(KEYINPUT80), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n611_), .A2(new_n617_), .A3(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n616_), .A2(KEYINPUT36), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n621_), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n611_), .A2(new_n617_), .A3(new_n619_), .A4(new_n623_), .ZN(new_n624_));
  AND3_X1   g423(.A1(new_n622_), .A2(KEYINPUT37), .A3(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(KEYINPUT37), .B1(new_n622_), .B2(new_n624_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G127gat), .B(G155gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT16), .ZN(new_n628_));
  XOR2_X1   g427(.A(G183gat), .B(G211gat), .Z(new_n629_));
  XNOR2_X1  g428(.A(new_n628_), .B(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT17), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(G231gat), .A2(G233gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n574_), .B(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n632_), .B1(new_n276_), .B2(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n635_), .B1(new_n276_), .B2(new_n634_), .ZN(new_n636_));
  AOI211_X1 g435(.A(new_n631_), .B(new_n630_), .C1(new_n634_), .C2(new_n279_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n637_), .B1(new_n279_), .B2(new_n634_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n636_), .A2(new_n638_), .ZN(new_n639_));
  NOR3_X1   g438(.A1(new_n625_), .A2(new_n626_), .A3(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT81), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n313_), .A2(new_n600_), .A3(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n419_), .A2(new_n420_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  OR3_X1    g443(.A1(new_n642_), .A2(G1gat), .A3(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT38), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n310_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n599_), .B1(new_n648_), .B2(new_n307_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT108), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n311_), .A2(KEYINPUT108), .A3(new_n599_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n622_), .A2(new_n624_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n654_), .A2(new_n639_), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n557_), .A2(new_n651_), .A3(new_n652_), .A4(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(G1gat), .B1(new_n656_), .B2(new_n644_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n645_), .A2(new_n646_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n647_), .A2(new_n657_), .A3(new_n658_), .ZN(G1324gat));
  INV_X1    g458(.A(new_n501_), .ZN(new_n660_));
  OAI21_X1  g459(.A(G8gat), .B1(new_n656_), .B2(new_n660_), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n661_), .A2(KEYINPUT39), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n661_), .A2(KEYINPUT39), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n501_), .A2(new_n570_), .ZN(new_n665_));
  OAI22_X1  g464(.A1(new_n663_), .A2(new_n664_), .B1(new_n642_), .B2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT40), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  OAI221_X1 g467(.A(KEYINPUT40), .B1(new_n642_), .B2(new_n665_), .C1(new_n663_), .C2(new_n664_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(G1325gat));
  OAI21_X1  g469(.A(G15gat), .B1(new_n656_), .B2(new_n545_), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n671_), .B(KEYINPUT109), .Z(new_n672_));
  OR2_X1    g471(.A1(new_n672_), .A2(KEYINPUT41), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(KEYINPUT41), .ZN(new_n674_));
  OR3_X1    g473(.A1(new_n642_), .A2(G15gat), .A3(new_n545_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n673_), .A2(new_n674_), .A3(new_n675_), .ZN(G1326gat));
  OAI21_X1  g475(.A(G22gat), .B1(new_n656_), .B2(new_n503_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT42), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n503_), .A2(G22gat), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n678_), .B1(new_n642_), .B2(new_n679_), .ZN(G1327gat));
  INV_X1    g479(.A(new_n311_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n654_), .A2(new_n639_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n600_), .A2(new_n683_), .ZN(new_n684_));
  OR3_X1    g483(.A1(new_n684_), .A2(G29gat), .A3(new_n644_), .ZN(new_n685_));
  AND3_X1   g484(.A1(new_n651_), .A2(new_n652_), .A3(new_n639_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT37), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n653_), .A2(new_n688_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n622_), .A2(KEYINPUT37), .A3(new_n624_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  AND3_X1   g490(.A1(new_n557_), .A2(new_n687_), .A3(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n687_), .B1(new_n557_), .B2(new_n691_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n686_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  OAI211_X1 g495(.A(KEYINPUT44), .B(new_n686_), .C1(new_n692_), .C2(new_n693_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n696_), .A2(new_n643_), .A3(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT110), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n698_), .A2(new_n699_), .A3(G29gat), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n698_), .B2(G29gat), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n685_), .B1(new_n700_), .B2(new_n701_), .ZN(G1328gat));
  INV_X1    g501(.A(KEYINPUT46), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n703_), .A2(KEYINPUT111), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n696_), .A2(new_n501_), .A3(new_n697_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(G36gat), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n703_), .A2(KEYINPUT111), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n660_), .A2(G36gat), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n683_), .A2(new_n557_), .A3(new_n599_), .A4(new_n709_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n710_), .A2(KEYINPUT45), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n710_), .A2(KEYINPUT45), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n708_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n705_), .B1(new_n707_), .B2(new_n714_), .ZN(new_n715_));
  AOI211_X1 g514(.A(new_n704_), .B(new_n713_), .C1(new_n706_), .C2(G36gat), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1329gat));
  NAND4_X1  g516(.A1(new_n696_), .A2(G43gat), .A3(new_n544_), .A4(new_n697_), .ZN(new_n718_));
  INV_X1    g517(.A(G43gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n719_), .B1(new_n684_), .B2(new_n545_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g521(.A1(new_n696_), .A2(G50gat), .A3(new_n376_), .A4(new_n697_), .ZN(new_n723_));
  INV_X1    g522(.A(G50gat), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n724_), .B1(new_n684_), .B2(new_n503_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n723_), .A2(new_n725_), .ZN(G1331gat));
  AND2_X1   g525(.A1(new_n557_), .A2(new_n655_), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n727_), .A2(new_n598_), .A3(new_n312_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(G57gat), .B1(new_n729_), .B2(new_n644_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n557_), .A2(new_n598_), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT112), .Z(new_n732_));
  AND2_X1   g531(.A1(new_n641_), .A2(new_n681_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n644_), .A2(G57gat), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n730_), .B1(new_n734_), .B2(new_n735_), .ZN(G1332gat));
  NAND4_X1  g535(.A1(new_n727_), .A2(new_n598_), .A3(new_n312_), .A4(new_n501_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(G64gat), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n738_), .A2(KEYINPUT113), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(KEYINPUT113), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT48), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n739_), .A2(KEYINPUT48), .A3(new_n740_), .ZN(new_n744_));
  OR3_X1    g543(.A1(new_n734_), .A2(G64gat), .A3(new_n660_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n743_), .A2(new_n744_), .A3(new_n745_), .ZN(G1333gat));
  OR3_X1    g545(.A1(new_n734_), .A2(G71gat), .A3(new_n545_), .ZN(new_n747_));
  OAI21_X1  g546(.A(G71gat), .B1(new_n729_), .B2(new_n545_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n748_), .A2(KEYINPUT49), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n748_), .A2(KEYINPUT49), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n747_), .B1(new_n749_), .B2(new_n750_), .ZN(G1334gat));
  NOR2_X1   g550(.A1(new_n503_), .A2(G78gat), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT114), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n727_), .A2(new_n598_), .A3(new_n312_), .A4(new_n376_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT50), .ZN(new_n755_));
  AND3_X1   g554(.A1(new_n754_), .A2(new_n755_), .A3(G78gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n754_), .B2(G78gat), .ZN(new_n757_));
  OAI22_X1  g556(.A1(new_n734_), .A2(new_n753_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT115), .ZN(G1335gat));
  NOR2_X1   g558(.A1(new_n313_), .A2(new_n682_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n732_), .A2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(G85gat), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n762_), .A2(new_n763_), .A3(new_n643_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n639_), .ZN(new_n765_));
  NOR3_X1   g564(.A1(new_n311_), .A2(new_n599_), .A3(new_n765_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n766_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT116), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  OAI211_X1 g568(.A(KEYINPUT116), .B(new_n766_), .C1(new_n692_), .C2(new_n693_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n644_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n764_), .B1(new_n763_), .B2(new_n771_), .ZN(G1336gat));
  INV_X1    g571(.A(G92gat), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n762_), .A2(new_n773_), .A3(new_n501_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n660_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n774_), .B1(new_n773_), .B2(new_n775_), .ZN(G1337gat));
  NAND4_X1  g575(.A1(new_n732_), .A2(new_n544_), .A3(new_n216_), .A4(new_n760_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n545_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n777_), .B1(new_n778_), .B2(new_n534_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT51), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT51), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n781_), .B(new_n777_), .C1(new_n778_), .C2(new_n534_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(G1338gat));
  OAI211_X1 g582(.A(new_n376_), .B(new_n766_), .C1(new_n692_), .C2(new_n693_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n785_));
  AND3_X1   g584(.A1(new_n784_), .A2(new_n785_), .A3(G106gat), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n785_), .B1(new_n784_), .B2(G106gat), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n376_), .A2(new_n217_), .ZN(new_n788_));
  OAI22_X1  g587(.A1(new_n786_), .A2(new_n787_), .B1(new_n761_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT53), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n791_));
  OAI221_X1 g590(.A(new_n791_), .B1(new_n761_), .B2(new_n788_), .C1(new_n787_), .C2(new_n786_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n792_), .ZN(G1339gat));
  INV_X1    g592(.A(KEYINPUT54), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n640_), .A2(new_n794_), .A3(new_n598_), .A4(new_n311_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n598_), .B1(new_n648_), .B2(new_n307_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n689_), .A2(new_n765_), .A3(new_n690_), .ZN(new_n797_));
  OAI21_X1  g596(.A(KEYINPUT54), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n795_), .A2(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n598_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n288_), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT12), .B1(new_n283_), .B2(new_n284_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n801_), .B1(new_n802_), .B2(new_n281_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(KEYINPUT117), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n277_), .B(new_n280_), .C1(new_n292_), .C2(KEYINPUT12), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n805_), .B1(new_n806_), .B2(new_n801_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n282_), .A2(new_n287_), .A3(KEYINPUT55), .A4(new_n288_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT117), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n806_), .A2(new_n809_), .A3(new_n801_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n804_), .A2(new_n807_), .A3(new_n808_), .A4(new_n810_), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n811_), .A2(KEYINPUT56), .A3(new_n298_), .ZN(new_n812_));
  AOI21_X1  g611(.A(KEYINPUT56), .B1(new_n811_), .B2(new_n298_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n800_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT118), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n800_), .B(KEYINPUT118), .C1(new_n812_), .C2(new_n813_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n304_), .A2(new_n306_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n579_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n579_), .B1(new_n566_), .B2(new_n574_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n591_), .B1(new_n576_), .B2(new_n820_), .ZN(new_n821_));
  AOI22_X1  g620(.A1(new_n596_), .A2(new_n597_), .B1(new_n819_), .B2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n818_), .A2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n816_), .A2(new_n817_), .A3(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT57), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n654_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n304_), .A2(new_n822_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n813_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n811_), .A2(KEYINPUT56), .A3(new_n298_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n828_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT119), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n832_), .A2(KEYINPUT58), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n831_), .A2(new_n834_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n812_), .A2(new_n813_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n833_), .B1(new_n836_), .B2(new_n828_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n835_), .A2(new_n691_), .A3(new_n837_), .ZN(new_n838_));
  AOI22_X1  g637(.A1(new_n814_), .A2(new_n815_), .B1(new_n818_), .B2(new_n822_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n654_), .B1(new_n839_), .B2(new_n817_), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n827_), .B(new_n838_), .C1(new_n840_), .C2(KEYINPUT57), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n799_), .B1(new_n841_), .B2(new_n639_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n552_), .A2(new_n544_), .A3(new_n643_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(G113gat), .B1(new_n844_), .B2(new_n599_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT59), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n846_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n843_), .ZN(new_n848_));
  AOI22_X1  g647(.A1(new_n831_), .A2(new_n834_), .B1(new_n690_), .B2(new_n689_), .ZN(new_n849_));
  AOI22_X1  g648(.A1(new_n824_), .A2(new_n826_), .B1(new_n849_), .B2(new_n837_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n824_), .A2(new_n653_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n825_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n765_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n853_));
  OAI211_X1 g652(.A(KEYINPUT59), .B(new_n848_), .C1(new_n853_), .C2(new_n799_), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n847_), .A2(KEYINPUT120), .A3(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(KEYINPUT120), .B1(new_n847_), .B2(new_n854_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n599_), .A2(G113gat), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n845_), .B1(new_n857_), .B2(new_n858_), .ZN(G1340gat));
  INV_X1    g658(.A(G120gat), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n860_), .B1(new_n311_), .B2(KEYINPUT60), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n844_), .B(new_n861_), .C1(KEYINPUT60), .C2(new_n860_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n313_), .B1(new_n847_), .B2(new_n854_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(new_n863_), .B2(new_n860_), .ZN(G1341gat));
  AOI21_X1  g663(.A(G127gat), .B1(new_n844_), .B2(new_n765_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n765_), .A2(G127gat), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(KEYINPUT121), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n865_), .B1(new_n857_), .B2(new_n867_), .ZN(G1342gat));
  AOI21_X1  g667(.A(G134gat), .B1(new_n844_), .B2(new_n654_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n691_), .ZN(new_n870_));
  XOR2_X1   g669(.A(KEYINPUT122), .B(G134gat), .Z(new_n871_));
  NOR2_X1   g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n869_), .B1(new_n857_), .B2(new_n872_), .ZN(G1343gat));
  NOR2_X1   g672(.A1(new_n842_), .A2(new_n544_), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n644_), .A2(new_n501_), .A3(new_n503_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n874_), .A2(new_n599_), .A3(new_n875_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g676(.A1(new_n874_), .A2(new_n312_), .A3(new_n875_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(KEYINPUT123), .B(G148gat), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n878_), .B(new_n879_), .ZN(G1345gat));
  NAND3_X1  g679(.A1(new_n874_), .A2(new_n765_), .A3(new_n875_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(KEYINPUT61), .B(G155gat), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n881_), .B(new_n882_), .ZN(G1346gat));
  NAND2_X1  g682(.A1(new_n874_), .A2(new_n875_), .ZN(new_n884_));
  OAI21_X1  g683(.A(G162gat), .B1(new_n884_), .B2(new_n870_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n654_), .A2(new_n327_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n885_), .B1(new_n884_), .B2(new_n886_), .ZN(G1347gat));
  NOR3_X1   g686(.A1(new_n660_), .A2(new_n553_), .A3(new_n376_), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n599_), .B(new_n888_), .C1(new_n853_), .C2(new_n799_), .ZN(new_n889_));
  OAI21_X1  g688(.A(G169gat), .B1(new_n889_), .B2(KEYINPUT62), .ZN(new_n890_));
  OAI21_X1  g689(.A(KEYINPUT62), .B1(new_n889_), .B2(KEYINPUT22), .ZN(new_n891_));
  MUX2_X1   g690(.A(G169gat), .B(new_n890_), .S(new_n891_), .Z(G1348gat));
  INV_X1    g691(.A(new_n888_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n842_), .A2(new_n893_), .ZN(new_n894_));
  AND3_X1   g693(.A1(new_n894_), .A2(G176gat), .A3(new_n312_), .ZN(new_n895_));
  AOI21_X1  g694(.A(G176gat), .B1(new_n894_), .B2(new_n681_), .ZN(new_n896_));
  OR2_X1    g695(.A1(new_n896_), .A2(KEYINPUT124), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(KEYINPUT124), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n895_), .B1(new_n897_), .B2(new_n898_), .ZN(G1349gat));
  NAND2_X1  g698(.A1(new_n894_), .A2(new_n765_), .ZN(new_n900_));
  MUX2_X1   g699(.A(new_n444_), .B(G183gat), .S(new_n900_), .Z(G1350gat));
  INV_X1    g700(.A(new_n894_), .ZN(new_n902_));
  OAI21_X1  g701(.A(G190gat), .B1(new_n902_), .B2(new_n870_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n654_), .A2(new_n443_), .ZN(new_n904_));
  XOR2_X1   g703(.A(new_n904_), .B(KEYINPUT125), .Z(new_n905_));
  OAI21_X1  g704(.A(new_n903_), .B1(new_n902_), .B2(new_n905_), .ZN(G1351gat));
  NOR2_X1   g705(.A1(new_n660_), .A2(new_n421_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n874_), .A2(new_n907_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n599_), .B1(KEYINPUT126), .B2(G197gat), .ZN(new_n909_));
  NAND2_X1  g708(.A1(KEYINPUT126), .A2(G197gat), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(KEYINPUT127), .ZN(new_n911_));
  OR3_X1    g710(.A1(new_n908_), .A2(new_n909_), .A3(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n911_), .B1(new_n908_), .B2(new_n909_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(G1352gat));
  NAND3_X1  g713(.A1(new_n874_), .A2(new_n312_), .A3(new_n907_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(G204gat), .ZN(G1353gat));
  XNOR2_X1  g715(.A(KEYINPUT63), .B(G211gat), .ZN(new_n917_));
  OR2_X1    g716(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n874_), .A2(new_n765_), .A3(new_n907_), .ZN(new_n919_));
  MUX2_X1   g718(.A(new_n917_), .B(new_n918_), .S(new_n919_), .Z(G1354gat));
  OAI21_X1  g719(.A(G218gat), .B1(new_n908_), .B2(new_n870_), .ZN(new_n921_));
  OR2_X1    g720(.A1(new_n653_), .A2(G218gat), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n921_), .B1(new_n908_), .B2(new_n922_), .ZN(G1355gat));
endmodule


