//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 1 1 0 0 1 1 1 1 1 0 0 1 0 0 1 0 1 0 1 0 0 1 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 0 1 0 1 0 0 1 1 0 0 0 1 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n628_, new_n629_,
    new_n630_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n712_, new_n713_, new_n714_, new_n715_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n845_, new_n846_, new_n848_, new_n849_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n856_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n893_, new_n895_,
    new_n896_, new_n898_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT29), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT3), .ZN(new_n209_));
  INV_X1    g008(.A(G141gat), .ZN(new_n210_));
  INV_X1    g009(.A(G148gat), .ZN(new_n211_));
  NAND4_X1  g010(.A1(new_n209_), .A2(new_n210_), .A3(new_n211_), .A4(KEYINPUT79), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT79), .ZN(new_n213_));
  OAI22_X1  g012(.A1(new_n213_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n214_));
  AND2_X1   g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G141gat), .A2(G148gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT2), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT2), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(G141gat), .A3(G148gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  AOI21_X1  g019(.A(KEYINPUT80), .B1(new_n215_), .B2(new_n220_), .ZN(new_n221_));
  AND4_X1   g020(.A1(KEYINPUT80), .A2(new_n220_), .A3(new_n214_), .A4(new_n212_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n208_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n207_), .B1(KEYINPUT1), .B2(new_n205_), .ZN(new_n224_));
  OR2_X1    g023(.A1(new_n205_), .A2(KEYINPUT1), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(G141gat), .A2(G148gat), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  AND3_X1   g027(.A1(new_n226_), .A2(new_n216_), .A3(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n204_), .B1(new_n223_), .B2(new_n230_), .ZN(new_n231_));
  XOR2_X1   g030(.A(G197gat), .B(G204gat), .Z(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT21), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G197gat), .B(G204gat), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT21), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G211gat), .B(G218gat), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT83), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(G218gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(G211gat), .ZN(new_n241_));
  INV_X1    g040(.A(G211gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(G218gat), .ZN(new_n243_));
  AND3_X1   g042(.A1(new_n241_), .A2(new_n243_), .A3(new_n238_), .ZN(new_n244_));
  OAI211_X1 g043(.A(new_n233_), .B(new_n236_), .C1(new_n239_), .C2(new_n244_), .ZN(new_n245_));
  OR2_X1    g044(.A1(new_n237_), .A2(new_n238_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n244_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n234_), .A2(new_n235_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n246_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  AND2_X1   g048(.A1(new_n245_), .A2(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n203_), .B1(new_n231_), .B2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n245_), .A2(new_n249_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT80), .ZN(new_n253_));
  AND2_X1   g052(.A1(new_n217_), .A2(new_n219_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n212_), .A2(new_n214_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n253_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n220_), .A2(KEYINPUT80), .A3(new_n214_), .A4(new_n212_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n229_), .B1(new_n258_), .B2(new_n208_), .ZN(new_n259_));
  OAI211_X1 g058(.A(new_n202_), .B(new_n252_), .C1(new_n259_), .C2(new_n204_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G78gat), .B(G106gat), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n251_), .A2(new_n260_), .A3(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT84), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT84), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n251_), .A2(new_n265_), .A3(new_n260_), .A4(new_n262_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n251_), .A2(new_n260_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(new_n261_), .ZN(new_n268_));
  AND3_X1   g067(.A1(new_n264_), .A2(new_n266_), .A3(new_n268_), .ZN(new_n269_));
  XOR2_X1   g068(.A(G22gat), .B(G50gat), .Z(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  XOR2_X1   g070(.A(KEYINPUT81), .B(KEYINPUT28), .Z(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n273_), .B1(new_n259_), .B2(new_n204_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n208_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n275_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n276_));
  NOR4_X1   g075(.A1(new_n276_), .A2(new_n229_), .A3(KEYINPUT29), .A4(new_n272_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n271_), .B1(new_n274_), .B2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n223_), .A2(new_n204_), .A3(new_n230_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(new_n272_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n259_), .A2(new_n204_), .A3(new_n273_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n280_), .A2(new_n270_), .A3(new_n281_), .ZN(new_n282_));
  AND3_X1   g081(.A1(new_n278_), .A2(new_n282_), .A3(KEYINPUT82), .ZN(new_n283_));
  AOI21_X1  g082(.A(KEYINPUT82), .B1(new_n278_), .B2(new_n282_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  OAI21_X1  g084(.A(KEYINPUT85), .B1(new_n269_), .B2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n264_), .A2(new_n266_), .A3(new_n268_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT85), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n287_), .B(new_n288_), .C1(new_n283_), .C2(new_n284_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n286_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n278_), .A2(new_n282_), .ZN(new_n291_));
  AND3_X1   g090(.A1(new_n268_), .A2(new_n263_), .A3(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT86), .ZN(new_n293_));
  AND2_X1   g092(.A1(new_n290_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT76), .ZN(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT25), .B(G183gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT26), .B(G190gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT24), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n299_), .B1(G169gat), .B2(G176gat), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT75), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n301_), .B1(G169gat), .B2(G176gat), .ZN(new_n302_));
  INV_X1    g101(.A(G169gat), .ZN(new_n303_));
  INV_X1    g102(.A(G176gat), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n303_), .A2(new_n304_), .A3(KEYINPUT75), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n300_), .A2(new_n302_), .A3(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n295_), .B1(new_n298_), .B2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G183gat), .A2(G190gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT23), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n305_), .A2(new_n302_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n309_), .B1(new_n310_), .B2(KEYINPUT24), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n307_), .A2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n298_), .A2(new_n306_), .A3(new_n295_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(G183gat), .ZN(new_n315_));
  INV_X1    g114(.A(G190gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n303_), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT22), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n319_), .A2(new_n304_), .A3(G169gat), .ZN(new_n320_));
  AOI22_X1  g119(.A1(new_n309_), .A2(new_n317_), .B1(new_n318_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n314_), .A2(new_n322_), .ZN(new_n323_));
  XOR2_X1   g122(.A(new_n323_), .B(KEYINPUT30), .Z(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(KEYINPUT77), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G71gat), .B(G99gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(G43gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G227gat), .A2(G233gat), .ZN(new_n328_));
  INV_X1    g127(.A(G15gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n327_), .B(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n323_), .B(KEYINPUT30), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT77), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n331_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n325_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT78), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G127gat), .B(G134gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G113gat), .B(G120gat), .ZN(new_n338_));
  AND2_X1   g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n337_), .A2(new_n338_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n336_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n337_), .ZN(new_n342_));
  XOR2_X1   g141(.A(G113gat), .B(G120gat), .Z(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n337_), .A2(new_n338_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n344_), .A2(KEYINPUT78), .A3(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n341_), .A2(new_n346_), .ZN(new_n347_));
  XOR2_X1   g146(.A(new_n347_), .B(KEYINPUT31), .Z(new_n348_));
  NAND3_X1  g147(.A1(new_n324_), .A2(KEYINPUT77), .A3(new_n331_), .ZN(new_n349_));
  AND3_X1   g148(.A1(new_n335_), .A2(new_n348_), .A3(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n348_), .B1(new_n335_), .B2(new_n349_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n344_), .A2(new_n345_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n223_), .A2(new_n230_), .A3(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n347_), .B1(new_n276_), .B2(new_n229_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n355_), .A2(new_n356_), .A3(KEYINPUT4), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT90), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n355_), .A2(new_n356_), .A3(KEYINPUT90), .A4(KEYINPUT4), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  XOR2_X1   g160(.A(KEYINPUT92), .B(KEYINPUT4), .Z(new_n362_));
  OAI211_X1 g161(.A(new_n347_), .B(new_n362_), .C1(new_n276_), .C2(new_n229_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G225gat), .A2(G233gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT91), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n361_), .A2(new_n367_), .ZN(new_n368_));
  AND2_X1   g167(.A1(new_n355_), .A2(new_n356_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(new_n364_), .ZN(new_n370_));
  XOR2_X1   g169(.A(G1gat), .B(G29gat), .Z(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n371_), .B(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G57gat), .B(G85gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n368_), .A2(new_n370_), .A3(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n366_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n370_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n375_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n377_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT27), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT88), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G226gat), .A2(G233gat), .ZN(new_n384_));
  XOR2_X1   g183(.A(new_n384_), .B(KEYINPUT19), .Z(new_n385_));
  NAND3_X1  g184(.A1(new_n299_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n386_));
  AND3_X1   g185(.A1(new_n306_), .A2(new_n309_), .A3(new_n386_), .ZN(new_n387_));
  XOR2_X1   g186(.A(KEYINPUT26), .B(G190gat), .Z(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT87), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT87), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n297_), .A2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n389_), .A2(new_n296_), .A3(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n387_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(new_n322_), .ZN(new_n394_));
  OAI211_X1 g193(.A(KEYINPUT20), .B(new_n385_), .C1(new_n394_), .C2(new_n252_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n250_), .B1(new_n314_), .B2(new_n322_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n383_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n313_), .ZN(new_n398_));
  NOR3_X1   g197(.A1(new_n398_), .A2(new_n307_), .A3(new_n311_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n252_), .B1(new_n399_), .B2(new_n321_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n385_), .A2(KEYINPUT20), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n321_), .B1(new_n387_), .B2(new_n392_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n401_), .B1(new_n250_), .B2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n400_), .A2(new_n403_), .A3(KEYINPUT88), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n397_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n314_), .A2(new_n250_), .A3(new_n322_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n394_), .A2(new_n252_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n406_), .A2(KEYINPUT20), .A3(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n385_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  XOR2_X1   g209(.A(G8gat), .B(G36gat), .Z(new_n411_));
  XNOR2_X1  g210(.A(G64gat), .B(G92gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  AND3_X1   g214(.A1(new_n405_), .A2(new_n410_), .A3(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n415_), .B1(new_n405_), .B2(new_n410_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n382_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n415_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(KEYINPUT96), .B(KEYINPUT20), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n421_), .B1(new_n250_), .B2(new_n402_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n385_), .B1(new_n400_), .B2(new_n422_), .ZN(new_n423_));
  OAI22_X1  g222(.A1(new_n423_), .A2(KEYINPUT97), .B1(new_n408_), .B2(new_n409_), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n423_), .A2(KEYINPUT97), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n419_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  AOI22_X1  g225(.A1(new_n397_), .A2(new_n404_), .B1(new_n409_), .B2(new_n408_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(new_n415_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n426_), .A2(KEYINPUT27), .A3(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n418_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n294_), .A2(new_n353_), .A3(new_n381_), .A4(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT98), .ZN(new_n433_));
  OAI211_X1 g232(.A(KEYINPUT32), .B(new_n415_), .C1(new_n424_), .C2(new_n425_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n415_), .A2(KEYINPUT32), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n427_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n433_), .B1(new_n381_), .B2(new_n437_), .ZN(new_n438_));
  NOR3_X1   g237(.A1(new_n378_), .A2(new_n379_), .A3(new_n375_), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT33), .B1(new_n439_), .B2(KEYINPUT94), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT94), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT33), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n377_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n416_), .A2(new_n417_), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n363_), .A2(new_n364_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n361_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(KEYINPUT95), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT95), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n361_), .A2(new_n448_), .A3(new_n445_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n376_), .B1(new_n369_), .B2(new_n365_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n447_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n440_), .A2(new_n443_), .A3(new_n444_), .A4(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n377_), .A2(new_n380_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n453_), .A2(KEYINPUT98), .A3(new_n436_), .A4(new_n434_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n438_), .A2(new_n452_), .A3(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n430_), .B1(new_n290_), .B2(new_n293_), .ZN(new_n456_));
  AOI22_X1  g255(.A1(new_n294_), .A2(new_n455_), .B1(new_n456_), .B2(new_n381_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n432_), .B1(new_n457_), .B2(new_n353_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G15gat), .B(G22gat), .ZN(new_n459_));
  INV_X1    g258(.A(G1gat), .ZN(new_n460_));
  INV_X1    g259(.A(G8gat), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT14), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n459_), .A2(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G1gat), .B(G8gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G29gat), .B(G36gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G43gat), .B(G50gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n466_), .B(new_n467_), .ZN(new_n468_));
  XOR2_X1   g267(.A(new_n465_), .B(new_n468_), .Z(new_n469_));
  NAND2_X1  g268(.A1(G229gat), .A2(G233gat), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n468_), .B(KEYINPUT15), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(new_n465_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n465_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(new_n468_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n474_), .A2(new_n476_), .A3(new_n470_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n472_), .A2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G113gat), .B(G141gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(KEYINPUT74), .ZN(new_n480_));
  XOR2_X1   g279(.A(G169gat), .B(G197gat), .Z(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n478_), .B(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n458_), .A2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(KEYINPUT99), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G232gat), .A2(G233gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT34), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n487_), .A2(KEYINPUT35), .ZN(new_n488_));
  OR3_X1    g287(.A1(KEYINPUT66), .A2(G99gat), .A3(G106gat), .ZN(new_n489_));
  OR2_X1    g288(.A1(new_n489_), .A2(KEYINPUT7), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G99gat), .A2(G106gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT6), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n489_), .A2(KEYINPUT7), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n490_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  XOR2_X1   g293(.A(G85gat), .B(G92gat), .Z(new_n495_));
  NAND4_X1  g294(.A1(new_n494_), .A2(KEYINPUT67), .A3(KEYINPUT8), .A4(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n494_), .A2(new_n495_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(KEYINPUT67), .A2(KEYINPUT8), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT9), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n500_), .A2(G85gat), .A3(G92gat), .ZN(new_n501_));
  AND2_X1   g300(.A1(new_n492_), .A2(new_n501_), .ZN(new_n502_));
  XOR2_X1   g301(.A(KEYINPUT10), .B(G99gat), .Z(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT64), .B(G106gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n495_), .A2(KEYINPUT9), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n502_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT65), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  AND2_X1   g308(.A1(new_n505_), .A2(new_n506_), .ZN(new_n510_));
  AOI21_X1  g309(.A(KEYINPUT65), .B1(new_n510_), .B2(new_n502_), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n496_), .B(new_n499_), .C1(new_n509_), .C2(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n488_), .B1(new_n512_), .B2(new_n473_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n507_), .A2(new_n508_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n510_), .A2(KEYINPUT65), .A3(new_n502_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n516_), .A2(new_n468_), .A3(new_n496_), .A4(new_n499_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n487_), .A2(KEYINPUT35), .ZN(new_n518_));
  XOR2_X1   g317(.A(new_n518_), .B(KEYINPUT70), .Z(new_n519_));
  AND3_X1   g318(.A1(new_n513_), .A2(new_n517_), .A3(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n519_), .B1(new_n513_), .B2(new_n517_), .ZN(new_n521_));
  OAI21_X1  g320(.A(KEYINPUT71), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  XOR2_X1   g321(.A(G190gat), .B(G218gat), .Z(new_n523_));
  XNOR2_X1  g322(.A(G134gat), .B(G162gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n523_), .B(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT36), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n527_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n525_), .A2(new_n526_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n522_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n529_), .ZN(new_n531_));
  OAI221_X1 g330(.A(KEYINPUT71), .B1(new_n531_), .B2(new_n527_), .C1(new_n520_), .C2(new_n521_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT37), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(KEYINPUT72), .A3(new_n535_), .ZN(new_n536_));
  AND2_X1   g335(.A1(new_n535_), .A2(KEYINPUT72), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n535_), .A2(KEYINPUT72), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n533_), .A2(new_n538_), .A3(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n536_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G127gat), .B(G155gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT16), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G183gat), .B(G211gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G231gat), .A2(G233gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n465_), .B(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G57gat), .B(G64gat), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n550_), .A2(KEYINPUT11), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(KEYINPUT11), .ZN(new_n552_));
  XOR2_X1   g351(.A(G71gat), .B(G78gat), .Z(new_n553_));
  NAND3_X1  g352(.A1(new_n551_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n552_), .A2(new_n553_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n549_), .B(new_n556_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n547_), .B1(new_n557_), .B2(KEYINPUT73), .ZN(new_n558_));
  OAI21_X1  g357(.A(KEYINPUT17), .B1(new_n557_), .B2(new_n547_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  OAI211_X1 g359(.A(KEYINPUT17), .B(new_n547_), .C1(new_n557_), .C2(KEYINPUT73), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n543_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT68), .ZN(new_n564_));
  INV_X1    g363(.A(new_n556_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n512_), .A2(new_n565_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n516_), .A2(new_n496_), .A3(new_n499_), .A4(new_n556_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n566_), .A2(KEYINPUT12), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT12), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n512_), .A2(new_n569_), .A3(new_n565_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G230gat), .A2(G233gat), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n564_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n572_), .ZN(new_n574_));
  AOI211_X1 g373(.A(KEYINPUT68), .B(new_n574_), .C1(new_n568_), .C2(new_n570_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n573_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n566_), .A2(new_n567_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(new_n574_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(new_n578_), .ZN(new_n579_));
  XOR2_X1   g378(.A(G120gat), .B(G148gat), .Z(new_n580_));
  XNOR2_X1  g379(.A(G176gat), .B(G204gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n579_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n571_), .A2(new_n572_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(KEYINPUT68), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n574_), .B1(new_n568_), .B2(new_n570_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(new_n564_), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n588_), .A2(new_n578_), .A3(new_n590_), .A4(new_n584_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n586_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT13), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n586_), .A2(KEYINPUT13), .A3(new_n591_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n563_), .A2(new_n596_), .ZN(new_n597_));
  AND2_X1   g396(.A1(new_n485_), .A2(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n381_), .A2(G1gat), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT100), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n598_), .A2(KEYINPUT100), .A3(new_n599_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n602_), .A2(KEYINPUT38), .A3(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n290_), .A2(new_n293_), .ZN(new_n605_));
  NOR4_X1   g404(.A1(new_n605_), .A2(new_n352_), .A3(new_n453_), .A4(new_n430_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n455_), .A2(new_n294_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n456_), .A2(new_n381_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n606_), .B1(new_n609_), .B2(new_n352_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n610_), .A2(new_n533_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n483_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n562_), .ZN(new_n613_));
  NOR3_X1   g412(.A1(new_n596_), .A2(new_n612_), .A3(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n611_), .A2(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(G1gat), .B1(new_n615_), .B2(new_n381_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT101), .ZN(new_n617_));
  AOI21_X1  g416(.A(KEYINPUT38), .B1(new_n602_), .B2(new_n603_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT102), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n618_), .A2(new_n619_), .ZN(new_n621_));
  OAI211_X1 g420(.A(new_n604_), .B(new_n617_), .C1(new_n620_), .C2(new_n621_), .ZN(G1324gat));
  OAI21_X1  g421(.A(G8gat), .B1(new_n615_), .B2(new_n431_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT39), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n598_), .A2(new_n461_), .A3(new_n430_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n626_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g426(.A(G15gat), .B1(new_n615_), .B2(new_n352_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n628_), .B(KEYINPUT41), .Z(new_n629_));
  NAND3_X1  g428(.A1(new_n598_), .A2(new_n329_), .A3(new_n353_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(G1326gat));
  OAI21_X1  g430(.A(G22gat), .B1(new_n615_), .B2(new_n294_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT42), .ZN(new_n633_));
  INV_X1    g432(.A(G22gat), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n598_), .A2(new_n634_), .A3(new_n605_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n636_), .B(KEYINPUT103), .Z(G1327gat));
  NOR2_X1   g436(.A1(new_n596_), .A2(new_n612_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(new_n613_), .ZN(new_n639_));
  OAI21_X1  g438(.A(KEYINPUT43), .B1(new_n610_), .B2(new_n543_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT43), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n353_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n642_));
  OAI211_X1 g441(.A(new_n641_), .B(new_n542_), .C1(new_n642_), .C2(new_n606_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n639_), .B1(new_n640_), .B2(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(KEYINPUT104), .B1(new_n644_), .B2(KEYINPUT44), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NOR3_X1   g445(.A1(new_n644_), .A2(KEYINPUT104), .A3(KEYINPUT44), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n644_), .A2(KEYINPUT44), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  NOR3_X1   g449(.A1(new_n648_), .A2(new_n381_), .A3(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(G29gat), .ZN(new_n652_));
  INV_X1    g451(.A(new_n596_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n533_), .A2(new_n613_), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT105), .Z(new_n655_));
  AND2_X1   g454(.A1(new_n653_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n485_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n453_), .A2(new_n652_), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n658_), .B(KEYINPUT106), .Z(new_n659_));
  OAI22_X1  g458(.A1(new_n651_), .A2(new_n652_), .B1(new_n657_), .B2(new_n659_), .ZN(G1328gat));
  INV_X1    g459(.A(new_n657_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n431_), .A2(G36gat), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(KEYINPUT45), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT45), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n661_), .A2(new_n665_), .A3(new_n662_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n431_), .B1(new_n644_), .B2(KEYINPUT44), .ZN(new_n668_));
  OAI211_X1 g467(.A(KEYINPUT107), .B(new_n668_), .C1(new_n646_), .C2(new_n647_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(G36gat), .ZN(new_n670_));
  INV_X1    g469(.A(new_n647_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(new_n645_), .ZN(new_n672_));
  AOI21_X1  g471(.A(KEYINPUT107), .B1(new_n672_), .B2(new_n668_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n667_), .B1(new_n670_), .B2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT108), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n675_), .A2(KEYINPUT46), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n676_), .ZN(new_n677_));
  OAI221_X1 g476(.A(new_n667_), .B1(new_n675_), .B2(KEYINPUT46), .C1(new_n670_), .C2(new_n673_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1329gat));
  INV_X1    g478(.A(G43gat), .ZN(new_n680_));
  NOR4_X1   g479(.A1(new_n648_), .A2(new_n680_), .A3(new_n352_), .A4(new_n650_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n680_), .B1(new_n657_), .B2(new_n352_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  OR3_X1    g482(.A1(new_n681_), .A2(KEYINPUT47), .A3(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(KEYINPUT47), .B1(new_n681_), .B2(new_n683_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(G1330gat));
  OR3_X1    g485(.A1(new_n657_), .A2(G50gat), .A3(new_n294_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n648_), .A2(new_n650_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT109), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n688_), .A2(new_n689_), .A3(new_n605_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(G50gat), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n689_), .B1(new_n688_), .B2(new_n605_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n687_), .B1(new_n691_), .B2(new_n692_), .ZN(G1331gat));
  NAND2_X1  g492(.A1(new_n596_), .A2(new_n612_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n694_), .A2(new_n613_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n611_), .A2(new_n695_), .ZN(new_n696_));
  OAI21_X1  g495(.A(G57gat), .B1(new_n696_), .B2(new_n381_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n610_), .A2(new_n694_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n698_), .A2(new_n543_), .A3(new_n562_), .ZN(new_n699_));
  OR2_X1    g498(.A1(new_n381_), .A2(G57gat), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n697_), .B1(new_n699_), .B2(new_n700_), .ZN(G1332gat));
  OAI21_X1  g500(.A(G64gat), .B1(new_n696_), .B2(new_n431_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT48), .ZN(new_n703_));
  OR3_X1    g502(.A1(new_n699_), .A2(G64gat), .A3(new_n431_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT110), .ZN(G1333gat));
  OAI21_X1  g505(.A(G71gat), .B1(new_n696_), .B2(new_n352_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT49), .ZN(new_n708_));
  OR3_X1    g507(.A1(new_n699_), .A2(G71gat), .A3(new_n352_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT111), .Z(G1334gat));
  OAI21_X1  g510(.A(G78gat), .B1(new_n696_), .B2(new_n294_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT50), .ZN(new_n713_));
  OR3_X1    g512(.A1(new_n699_), .A2(G78gat), .A3(new_n294_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT112), .ZN(G1335gat));
  NAND2_X1  g515(.A1(new_n698_), .A2(new_n655_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT113), .ZN(new_n718_));
  AOI21_X1  g517(.A(G85gat), .B1(new_n718_), .B2(new_n453_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT114), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n596_), .A2(new_n612_), .A3(new_n613_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n721_), .B1(new_n640_), .B2(new_n643_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n722_), .A2(G85gat), .A3(new_n453_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n720_), .A2(new_n723_), .ZN(G1336gat));
  INV_X1    g523(.A(G92gat), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n718_), .A2(new_n725_), .A3(new_n430_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n722_), .ZN(new_n727_));
  OAI21_X1  g526(.A(G92gat), .B1(new_n727_), .B2(new_n431_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT115), .ZN(G1337gat));
  NAND3_X1  g529(.A1(new_n718_), .A2(new_n353_), .A3(new_n503_), .ZN(new_n731_));
  OAI21_X1  g530(.A(G99gat), .B1(new_n727_), .B2(new_n352_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT51), .ZN(G1338gat));
  XNOR2_X1  g533(.A(KEYINPUT118), .B(KEYINPUT52), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n721_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n643_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n641_), .B1(new_n458_), .B2(new_n542_), .ZN(new_n739_));
  OAI211_X1 g538(.A(new_n605_), .B(new_n737_), .C1(new_n738_), .C2(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(G106gat), .B1(new_n740_), .B2(KEYINPUT117), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT117), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n742_), .B1(new_n722_), .B2(new_n605_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n736_), .B1(new_n741_), .B2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT120), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  OAI211_X1 g545(.A(KEYINPUT120), .B(new_n736_), .C1(new_n741_), .C2(new_n743_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n740_), .A2(KEYINPUT117), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n722_), .A2(new_n742_), .A3(new_n605_), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n748_), .A2(new_n749_), .A3(G106gat), .A4(new_n735_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT119), .ZN(new_n751_));
  INV_X1    g550(.A(G106gat), .ZN(new_n752_));
  AOI211_X1 g551(.A(new_n294_), .B(new_n721_), .C1(new_n640_), .C2(new_n643_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n753_), .B2(new_n742_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT119), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n754_), .A2(new_n755_), .A3(new_n735_), .A4(new_n748_), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n746_), .A2(new_n747_), .A3(new_n751_), .A4(new_n756_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n605_), .A2(new_n504_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n718_), .A2(new_n758_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT116), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n757_), .A2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(KEYINPUT53), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT53), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n757_), .A2(new_n763_), .A3(new_n760_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n762_), .A2(new_n764_), .ZN(G1339gat));
  INV_X1    g564(.A(KEYINPUT54), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n597_), .A2(new_n766_), .A3(new_n612_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n766_), .B1(new_n597_), .B2(new_n612_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n591_), .A2(new_n483_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT56), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n568_), .A2(new_n574_), .A3(new_n570_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT55), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n774_), .B1(new_n587_), .B2(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n776_), .B1(new_n576_), .B2(new_n775_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n773_), .B1(new_n777_), .B2(new_n584_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n588_), .A2(new_n775_), .A3(new_n590_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n774_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n780_), .B1(new_n589_), .B2(KEYINPUT55), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n584_), .B1(new_n779_), .B2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT56), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n772_), .B1(new_n778_), .B2(new_n783_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n478_), .A2(new_n482_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n482_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n786_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT121), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n470_), .B1(new_n475_), .B2(new_n468_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n789_), .B1(new_n474_), .B2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n787_), .A2(new_n788_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n785_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n794_), .B1(new_n586_), .B2(new_n591_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n534_), .B1(new_n784_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT122), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n772_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n782_), .A2(KEYINPUT56), .ZN(new_n800_));
  AOI211_X1 g599(.A(new_n773_), .B(new_n584_), .C1(new_n779_), .C2(new_n781_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n799_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n795_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n804_), .A2(KEYINPUT122), .A3(new_n534_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT57), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n798_), .A2(new_n805_), .A3(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT123), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n808_), .B1(new_n591_), .B2(new_n793_), .ZN(new_n809_));
  AND3_X1   g608(.A1(new_n591_), .A2(new_n793_), .A3(new_n808_), .ZN(new_n810_));
  OAI22_X1  g609(.A1(new_n800_), .A2(new_n801_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT58), .ZN(new_n812_));
  AOI22_X1  g611(.A1(new_n811_), .A2(new_n812_), .B1(new_n536_), .B2(new_n541_), .ZN(new_n813_));
  OAI221_X1 g612(.A(KEYINPUT58), .B1(new_n810_), .B2(new_n809_), .C1(new_n800_), .C2(new_n801_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  OAI211_X1 g614(.A(KEYINPUT57), .B(new_n534_), .C1(new_n784_), .C2(new_n795_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT124), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n804_), .A2(KEYINPUT124), .A3(KEYINPUT57), .A4(new_n534_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n815_), .A2(new_n818_), .A3(new_n819_), .ZN(new_n820_));
  OAI211_X1 g619(.A(KEYINPUT125), .B(new_n613_), .C1(new_n807_), .C2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  AOI22_X1  g621(.A1(new_n814_), .A2(new_n813_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n798_), .A2(new_n805_), .A3(new_n806_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n824_), .A3(new_n819_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT125), .B1(new_n825_), .B2(new_n613_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n771_), .B1(new_n822_), .B2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT59), .ZN(new_n828_));
  NOR4_X1   g627(.A1(new_n605_), .A2(new_n352_), .A3(new_n381_), .A4(new_n430_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n827_), .A2(new_n828_), .A3(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n825_), .A2(new_n613_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n771_), .A2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(new_n829_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(KEYINPUT59), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n830_), .A2(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(G113gat), .B1(new_n835_), .B2(new_n612_), .ZN(new_n836_));
  OR3_X1    g635(.A1(new_n833_), .A2(G113gat), .A3(new_n612_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(G1340gat));
  OAI21_X1  g637(.A(G120gat), .B1(new_n835_), .B2(new_n653_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n833_), .ZN(new_n840_));
  INV_X1    g639(.A(G120gat), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n841_), .B1(new_n653_), .B2(KEYINPUT60), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n840_), .B(new_n842_), .C1(KEYINPUT60), .C2(new_n841_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n839_), .A2(new_n843_), .ZN(G1341gat));
  OAI21_X1  g643(.A(G127gat), .B1(new_n835_), .B2(new_n613_), .ZN(new_n845_));
  OR3_X1    g644(.A1(new_n833_), .A2(G127gat), .A3(new_n613_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(G1342gat));
  OAI21_X1  g646(.A(G134gat), .B1(new_n835_), .B2(new_n543_), .ZN(new_n848_));
  OR3_X1    g647(.A1(new_n833_), .A2(G134gat), .A3(new_n534_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(G1343gat));
  AOI21_X1  g649(.A(new_n353_), .B1(new_n771_), .B2(new_n831_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n456_), .A2(new_n453_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n853_), .A2(new_n612_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(new_n210_), .ZN(G1344gat));
  NOR2_X1   g654(.A1(new_n853_), .A2(new_n653_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(new_n211_), .ZN(G1345gat));
  NOR2_X1   g656(.A1(new_n853_), .A2(new_n613_), .ZN(new_n858_));
  XOR2_X1   g657(.A(KEYINPUT61), .B(G155gat), .Z(new_n859_));
  XNOR2_X1  g658(.A(new_n858_), .B(new_n859_), .ZN(G1346gat));
  INV_X1    g659(.A(G162gat), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n853_), .A2(new_n861_), .A3(new_n543_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n851_), .A2(new_n533_), .A3(new_n852_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n861_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT126), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n863_), .A2(KEYINPUT126), .A3(new_n861_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n862_), .B1(new_n866_), .B2(new_n867_), .ZN(G1347gat));
  NOR2_X1   g667(.A1(new_n431_), .A2(new_n453_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n869_), .A2(new_n294_), .A3(new_n353_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n827_), .A2(new_n319_), .A3(new_n483_), .A4(new_n871_), .ZN(new_n872_));
  AND3_X1   g671(.A1(new_n872_), .A2(KEYINPUT62), .A3(new_n303_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(KEYINPUT62), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT62), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n827_), .A2(new_n875_), .A3(new_n483_), .A4(new_n871_), .ZN(new_n876_));
  AND2_X1   g675(.A1(new_n876_), .A2(G169gat), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n873_), .B1(new_n874_), .B2(new_n877_), .ZN(G1348gat));
  NAND2_X1  g677(.A1(new_n832_), .A2(new_n871_), .ZN(new_n879_));
  NOR3_X1   g678(.A1(new_n879_), .A2(new_n304_), .A3(new_n653_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n827_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n881_), .A2(new_n870_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(new_n596_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n880_), .B1(new_n883_), .B2(new_n304_), .ZN(G1349gat));
  NOR2_X1   g683(.A1(new_n613_), .A2(new_n296_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n827_), .A2(new_n871_), .A3(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT127), .ZN(new_n887_));
  OR2_X1    g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n315_), .B1(new_n879_), .B2(new_n613_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n886_), .A2(new_n887_), .ZN(new_n890_));
  AND3_X1   g689(.A1(new_n888_), .A2(new_n889_), .A3(new_n890_), .ZN(G1350gat));
  NAND4_X1  g690(.A1(new_n882_), .A2(new_n389_), .A3(new_n391_), .A4(new_n533_), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n881_), .A2(new_n543_), .A3(new_n870_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n316_), .B2(new_n893_), .ZN(G1351gat));
  AND3_X1   g693(.A1(new_n851_), .A2(new_n605_), .A3(new_n869_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n483_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n596_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g698(.A(new_n613_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n895_), .A2(new_n900_), .ZN(new_n901_));
  OR2_X1    g700(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n901_), .B(new_n902_), .ZN(G1354gat));
  NAND3_X1  g702(.A1(new_n895_), .A2(new_n240_), .A3(new_n533_), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n895_), .A2(new_n542_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n905_), .B2(new_n240_), .ZN(G1355gat));
endmodule


