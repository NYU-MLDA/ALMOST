//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 0 1 1 0 0 0 1 0 0 0 0 0 1 0 0 0 1 1 0 0 1 1 1 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 0 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n727_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n777_, new_n778_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n897_, new_n898_, new_n900_,
    new_n902_, new_n903_, new_n905_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_, new_n924_, new_n926_, new_n927_, new_n929_, new_n930_,
    new_n931_, new_n933_, new_n934_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n946_, new_n947_, new_n948_, new_n950_, new_n951_, new_n952_;
  INV_X1    g000(.A(KEYINPUT102), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G8gat), .B(G36gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT18), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G64gat), .B(G92gat), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT32), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT91), .B(G204gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G197gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n210_), .B1(G197gat), .B2(G204gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT21), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G211gat), .B(G218gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(G204gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(G197gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(KEYINPUT90), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT92), .ZN(new_n219_));
  INV_X1    g018(.A(G197gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n209_), .A2(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n218_), .B1(new_n219_), .B2(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n222_), .B1(new_n219_), .B2(new_n221_), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n215_), .B1(new_n223_), .B2(KEYINPUT21), .ZN(new_n224_));
  NOR3_X1   g023(.A1(new_n211_), .A2(new_n212_), .A3(new_n214_), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(KEYINPUT94), .ZN(new_n228_));
  XOR2_X1   g027(.A(KEYINPUT22), .B(G169gat), .Z(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT95), .ZN(new_n230_));
  XOR2_X1   g029(.A(KEYINPUT83), .B(G176gat), .Z(new_n231_));
  AOI21_X1  g030(.A(new_n228_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n232_), .A2(KEYINPUT96), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(KEYINPUT96), .ZN(new_n234_));
  INV_X1    g033(.A(G183gat), .ZN(new_n235_));
  INV_X1    g034(.A(G190gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(KEYINPUT23), .B1(new_n235_), .B2(new_n236_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT81), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  OR3_X1    g039(.A1(new_n235_), .A2(new_n236_), .A3(KEYINPUT23), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  AOI22_X1  g041(.A1(new_n233_), .A2(new_n234_), .B1(new_n237_), .B2(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n235_), .A2(KEYINPUT25), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n235_), .A2(KEYINPUT25), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT26), .B(G190gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n241_), .A2(new_n238_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n227_), .A2(KEYINPUT24), .ZN(new_n252_));
  INV_X1    g051(.A(G169gat), .ZN(new_n253_));
  INV_X1    g052(.A(G176gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  MUX2_X1   g054(.A(KEYINPUT24), .B(new_n252_), .S(new_n255_), .Z(new_n256_));
  AND3_X1   g055(.A1(new_n250_), .A2(new_n251_), .A3(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n226_), .B1(new_n243_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G226gat), .A2(G233gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT19), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT20), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n224_), .A2(new_n225_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n244_), .B1(KEYINPUT80), .B2(new_n246_), .ZN(new_n264_));
  OAI211_X1 g063(.A(new_n264_), .B(new_n249_), .C1(KEYINPUT80), .C2(new_n246_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n242_), .A2(new_n256_), .A3(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n251_), .A2(new_n237_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n253_), .A2(KEYINPUT22), .ZN(new_n268_));
  OR3_X1    g067(.A1(new_n253_), .A2(KEYINPUT82), .A3(KEYINPUT22), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT82), .B1(new_n253_), .B2(KEYINPUT22), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n231_), .A2(new_n268_), .A3(new_n269_), .A4(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n267_), .A2(new_n271_), .A3(new_n227_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n266_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n262_), .B1(new_n263_), .B2(new_n274_), .ZN(new_n275_));
  AND3_X1   g074(.A1(new_n258_), .A2(new_n261_), .A3(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n262_), .B1(new_n226_), .B2(new_n273_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n242_), .A2(new_n237_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n234_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n232_), .A2(KEYINPUT96), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n278_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n257_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n281_), .A2(new_n263_), .A3(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n261_), .B1(new_n277_), .B2(new_n283_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n208_), .B1(new_n276_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT99), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  OAI211_X1 g086(.A(KEYINPUT99), .B(new_n208_), .C1(new_n276_), .C2(new_n284_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n277_), .A2(new_n283_), .A3(new_n261_), .ZN(new_n289_));
  AND2_X1   g088(.A1(new_n258_), .A2(new_n275_), .ZN(new_n290_));
  OAI211_X1 g089(.A(new_n289_), .B(new_n207_), .C1(new_n290_), .C2(new_n261_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n287_), .A2(new_n288_), .A3(new_n291_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(G155gat), .A2(G162gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT87), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G155gat), .A2(G162gat), .ZN(new_n296_));
  OR2_X1    g095(.A1(G141gat), .A2(G148gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT3), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT88), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G141gat), .A2(G148gat), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT2), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n304_));
  OAI211_X1 g103(.A(new_n303_), .B(new_n304_), .C1(new_n297_), .C2(KEYINPUT3), .ZN(new_n305_));
  OAI211_X1 g104(.A(new_n295_), .B(new_n296_), .C1(new_n300_), .C2(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n296_), .B(KEYINPUT1), .ZN(new_n307_));
  OAI211_X1 g106(.A(new_n297_), .B(new_n301_), .C1(new_n294_), .C2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  XOR2_X1   g108(.A(G127gat), .B(G134gat), .Z(new_n310_));
  XOR2_X1   g109(.A(G113gat), .B(G120gat), .Z(new_n311_));
  XOR2_X1   g110(.A(new_n310_), .B(new_n311_), .Z(new_n312_));
  NAND2_X1  g111(.A1(new_n309_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n312_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n314_), .A2(new_n306_), .A3(new_n308_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n313_), .A2(KEYINPUT4), .A3(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G225gat), .A2(G233gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT97), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT4), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n309_), .A2(new_n319_), .A3(new_n312_), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n316_), .A2(KEYINPUT98), .A3(new_n318_), .A4(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n318_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n313_), .A2(new_n315_), .A3(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n321_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n320_), .A2(new_n318_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(KEYINPUT98), .B1(new_n326_), .B2(new_n316_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n324_), .A2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G1gat), .B(G29gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(G85gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(KEYINPUT0), .B(G57gat), .ZN(new_n331_));
  XOR2_X1   g130(.A(new_n330_), .B(new_n331_), .Z(new_n332_));
  NAND3_X1  g131(.A1(new_n328_), .A2(KEYINPUT100), .A3(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT98), .ZN(new_n334_));
  INV_X1    g133(.A(new_n316_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n334_), .B1(new_n335_), .B2(new_n325_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n336_), .A2(new_n332_), .A3(new_n323_), .A4(new_n321_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT100), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n332_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n340_), .B1(new_n324_), .B2(new_n327_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n333_), .A2(new_n339_), .A3(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  XOR2_X1   g142(.A(new_n337_), .B(KEYINPUT33), .Z(new_n344_));
  INV_X1    g143(.A(new_n206_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n289_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n261_), .B1(new_n258_), .B2(new_n275_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n345_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  OAI211_X1 g147(.A(new_n206_), .B(new_n289_), .C1(new_n290_), .C2(new_n261_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n316_), .A2(new_n322_), .A3(new_n320_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n313_), .A2(new_n315_), .A3(new_n318_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n350_), .A2(new_n340_), .A3(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n348_), .A2(new_n349_), .A3(new_n352_), .ZN(new_n353_));
  OAI22_X1  g152(.A1(new_n292_), .A2(new_n343_), .B1(new_n344_), .B2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G78gat), .B(G106gat), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G228gat), .A2(G233gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n309_), .A2(KEYINPUT29), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n226_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n357_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n358_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n360_), .B1(new_n263_), .B2(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n356_), .B1(new_n359_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n359_), .A2(new_n362_), .A3(new_n356_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  OR3_X1    g165(.A1(new_n309_), .A2(KEYINPUT89), .A3(KEYINPUT29), .ZN(new_n367_));
  OAI21_X1  g166(.A(KEYINPUT89), .B1(new_n309_), .B2(KEYINPUT29), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G22gat), .B(G50gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT28), .ZN(new_n370_));
  AND3_X1   g169(.A1(new_n367_), .A2(new_n368_), .A3(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n370_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n373_), .B1(new_n363_), .B2(KEYINPUT93), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n366_), .A2(new_n374_), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n364_), .A2(KEYINPUT93), .A3(new_n365_), .A4(new_n373_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G227gat), .A2(G233gat), .ZN(new_n379_));
  INV_X1    g178(.A(G15gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(G71gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(KEYINPUT84), .B(G43gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(G99gat), .ZN(new_n385_));
  OR2_X1    g184(.A1(new_n383_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n383_), .A2(new_n385_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT85), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT85), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n386_), .A2(new_n390_), .A3(new_n387_), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n266_), .A2(KEYINPUT30), .A3(new_n272_), .ZN(new_n392_));
  AOI21_X1  g191(.A(KEYINPUT30), .B1(new_n266_), .B2(new_n272_), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n389_), .B(new_n391_), .C1(new_n392_), .C2(new_n393_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n392_), .A2(new_n393_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n391_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT86), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n394_), .A2(new_n397_), .A3(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT31), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT31), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n394_), .A2(new_n397_), .A3(new_n398_), .A4(new_n401_), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n400_), .A2(new_n312_), .A3(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n312_), .B1(new_n400_), .B2(new_n402_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n378_), .A2(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n345_), .B1(new_n276_), .B2(new_n284_), .ZN(new_n407_));
  AND3_X1   g206(.A1(new_n349_), .A2(new_n407_), .A3(KEYINPUT27), .ZN(new_n408_));
  AOI21_X1  g207(.A(KEYINPUT27), .B1(new_n348_), .B2(new_n349_), .ZN(new_n409_));
  NOR3_X1   g208(.A1(new_n408_), .A2(new_n409_), .A3(new_n342_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n377_), .A2(new_n405_), .ZN(new_n411_));
  OAI211_X1 g210(.A(new_n375_), .B(new_n376_), .C1(new_n403_), .C2(new_n404_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  AOI22_X1  g212(.A1(new_n354_), .A2(new_n406_), .B1(new_n410_), .B2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G113gat), .B(G141gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G169gat), .B(G197gat), .ZN(new_n416_));
  XOR2_X1   g215(.A(new_n415_), .B(new_n416_), .Z(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G1gat), .B(G8gat), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G15gat), .B(G22gat), .ZN(new_n421_));
  INV_X1    g220(.A(G8gat), .ZN(new_n422_));
  INV_X1    g221(.A(G1gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT75), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT75), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(G1gat), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n422_), .B1(new_n424_), .B2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT14), .ZN(new_n428_));
  OAI211_X1 g227(.A(KEYINPUT76), .B(new_n421_), .C1(new_n427_), .C2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(KEYINPUT75), .B(G1gat), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT14), .B1(new_n431_), .B2(new_n422_), .ZN(new_n432_));
  AOI21_X1  g231(.A(KEYINPUT76), .B1(new_n432_), .B2(new_n421_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n420_), .B1(new_n430_), .B2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G43gat), .B(G50gat), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G29gat), .B(G36gat), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n437_), .A2(KEYINPUT71), .ZN(new_n438_));
  INV_X1    g237(.A(G36gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(G29gat), .ZN(new_n440_));
  INV_X1    g239(.A(G29gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(G36gat), .ZN(new_n442_));
  AND3_X1   g241(.A1(new_n440_), .A2(new_n442_), .A3(KEYINPUT71), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n436_), .B1(new_n438_), .B2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n440_), .A2(new_n442_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT71), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n437_), .A2(KEYINPUT71), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n447_), .A2(new_n448_), .A3(new_n435_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n444_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT15), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT76), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n424_), .A2(new_n426_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n428_), .B1(new_n454_), .B2(G8gat), .ZN(new_n455_));
  INV_X1    g254(.A(new_n421_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n453_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n457_), .A2(new_n429_), .A3(new_n419_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n444_), .A2(KEYINPUT15), .A3(new_n449_), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n434_), .A2(new_n452_), .A3(new_n458_), .A4(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n450_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n462_), .B1(new_n434_), .B2(new_n458_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G229gat), .A2(G233gat), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NOR3_X1   g264(.A1(new_n461_), .A2(new_n463_), .A3(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT78), .ZN(new_n467_));
  AND3_X1   g266(.A1(new_n434_), .A2(new_n458_), .A3(new_n462_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n467_), .B1(new_n468_), .B2(new_n463_), .ZN(new_n469_));
  NOR3_X1   g268(.A1(new_n430_), .A2(new_n433_), .A3(new_n420_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n419_), .B1(new_n457_), .B2(new_n429_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n450_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n434_), .A2(new_n458_), .A3(new_n462_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n472_), .A2(KEYINPUT78), .A3(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n469_), .A2(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n466_), .B1(new_n475_), .B2(new_n465_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n418_), .B1(new_n476_), .B2(KEYINPUT79), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT79), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n464_), .B1(new_n469_), .B2(new_n474_), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n478_), .B(new_n417_), .C1(new_n479_), .C2(new_n466_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(KEYINPUT101), .B1(new_n414_), .B2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n354_), .A2(new_n406_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n410_), .A2(new_n413_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT101), .ZN(new_n486_));
  NOR3_X1   g285(.A1(new_n468_), .A2(new_n463_), .A3(new_n467_), .ZN(new_n487_));
  AOI21_X1  g286(.A(KEYINPUT78), .B1(new_n472_), .B2(new_n473_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n465_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n466_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n417_), .B1(new_n491_), .B2(new_n478_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n480_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n485_), .A2(new_n486_), .A3(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n482_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT37), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G85gat), .B(G92gat), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT9), .ZN(new_n501_));
  XOR2_X1   g300(.A(KEYINPUT10), .B(G99gat), .Z(new_n502_));
  INV_X1    g301(.A(G106gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G99gat), .A2(G106gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT6), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT6), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n507_), .A2(G99gat), .A3(G106gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(KEYINPUT64), .B(G92gat), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT9), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n510_), .A2(new_n511_), .A3(G85gat), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n501_), .A2(new_n504_), .A3(new_n509_), .A4(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT8), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n507_), .B1(G99gat), .B2(G106gat), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n505_), .A2(KEYINPUT6), .ZN(new_n516_));
  OAI21_X1  g315(.A(KEYINPUT65), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT65), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n506_), .A2(new_n508_), .A3(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT7), .ZN(new_n520_));
  INV_X1    g319(.A(G99gat), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n520_), .A2(new_n521_), .A3(new_n503_), .ZN(new_n522_));
  OAI21_X1  g321(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n523_));
  AND2_X1   g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n517_), .A2(new_n519_), .A3(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n514_), .B1(new_n525_), .B2(new_n500_), .ZN(new_n526_));
  AOI211_X1 g325(.A(KEYINPUT8), .B(new_n499_), .C1(new_n524_), .C2(new_n509_), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n450_), .B(new_n513_), .C1(new_n526_), .C2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT72), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n524_), .A2(new_n509_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n530_), .A2(new_n514_), .A3(new_n500_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n522_), .A2(new_n523_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n532_), .B1(KEYINPUT65), .B2(new_n509_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n499_), .B1(new_n533_), .B2(new_n519_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n531_), .B1(new_n534_), .B2(new_n514_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT72), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n535_), .A2(new_n536_), .A3(new_n450_), .A4(new_n513_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n529_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT74), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G232gat), .A2(G233gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT34), .ZN(new_n541_));
  XNOR2_X1  g340(.A(KEYINPUT70), .B(KEYINPUT35), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n539_), .B1(new_n541_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n459_), .ZN(new_n545_));
  AOI21_X1  g344(.A(KEYINPUT15), .B1(new_n444_), .B2(new_n449_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n513_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n544_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n538_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n541_), .A2(new_n543_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n538_), .A2(new_n549_), .A3(new_n551_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n553_), .A2(KEYINPUT73), .A3(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G190gat), .B(G218gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G134gat), .B(G162gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n558_), .A2(KEYINPUT36), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n555_), .A2(new_n560_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n553_), .A2(KEYINPUT73), .A3(new_n554_), .A4(new_n559_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n558_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT36), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n567_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n498_), .B1(new_n563_), .B2(new_n569_), .ZN(new_n570_));
  AOI211_X1 g369(.A(KEYINPUT37), .B(new_n568_), .C1(new_n561_), .C2(new_n562_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G176gat), .B(G204gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT69), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G120gat), .B(G148gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n576_), .B(new_n577_), .Z(new_n578_));
  OR2_X1    g377(.A1(new_n578_), .A2(KEYINPUT67), .ZN(new_n579_));
  NOR2_X1   g378(.A1(KEYINPUT66), .A2(G71gat), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(G78gat), .ZN(new_n582_));
  NAND2_X1  g381(.A1(KEYINPUT66), .A2(G71gat), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n581_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n583_), .ZN(new_n585_));
  OAI21_X1  g384(.A(G78gat), .B1(new_n585_), .B2(new_n580_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G57gat), .B(G64gat), .ZN(new_n587_));
  AOI22_X1  g386(.A1(new_n584_), .A2(new_n586_), .B1(KEYINPUT11), .B2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(KEYINPUT11), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n584_), .A2(new_n586_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n588_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  OAI211_X1 g390(.A(new_n591_), .B(new_n513_), .C1(new_n526_), .C2(new_n527_), .ZN(new_n592_));
  INV_X1    g391(.A(G230gat), .ZN(new_n593_));
  INV_X1    g392(.A(G233gat), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n592_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT12), .ZN(new_n598_));
  INV_X1    g397(.A(new_n591_), .ZN(new_n599_));
  AND3_X1   g398(.A1(new_n548_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n598_), .B1(new_n548_), .B2(new_n599_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n597_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n548_), .A2(new_n599_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(new_n592_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(new_n595_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n602_), .A2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n579_), .B(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT13), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n434_), .A2(new_n458_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n610_), .A2(G231gat), .A3(G233gat), .ZN(new_n611_));
  NAND2_X1  g410(.A1(G231gat), .A2(G233gat), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n434_), .A2(new_n458_), .A3(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(new_n591_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT77), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G127gat), .B(G155gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT16), .ZN(new_n619_));
  XOR2_X1   g418(.A(G183gat), .B(G211gat), .Z(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(KEYINPUT17), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n617_), .B(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT17), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n615_), .A2(new_n626_), .A3(new_n621_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n625_), .A2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n572_), .A2(new_n609_), .A3(new_n628_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n202_), .B1(new_n497_), .B2(new_n629_), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n572_), .A2(new_n628_), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n496_), .A2(KEYINPUT102), .A3(new_n609_), .A4(new_n631_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n630_), .A2(new_n342_), .A3(new_n431_), .A4(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT38), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT103), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n568_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n636_), .B1(new_n414_), .B2(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n485_), .A2(KEYINPUT103), .A3(new_n637_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n609_), .A2(new_n494_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n628_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n641_), .A2(new_n342_), .A3(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(G1gat), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n633_), .A2(new_n634_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n635_), .A2(new_n646_), .A3(new_n647_), .ZN(G1324gat));
  INV_X1    g447(.A(new_n409_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n349_), .A2(new_n407_), .A3(KEYINPUT27), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n630_), .A2(new_n422_), .A3(new_n651_), .A4(new_n632_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n641_), .A2(new_n651_), .A3(new_n644_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(KEYINPUT104), .B(KEYINPUT39), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n653_), .A2(G8gat), .A3(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n654_), .B1(new_n653_), .B2(G8gat), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n652_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT40), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n657_), .B(new_n658_), .ZN(G1325gat));
  AND2_X1   g458(.A1(new_n630_), .A2(new_n632_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n660_), .A2(new_n380_), .A3(new_n405_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n641_), .A2(new_n405_), .A3(new_n644_), .ZN(new_n662_));
  AOI21_X1  g461(.A(KEYINPUT41), .B1(new_n662_), .B2(G15gat), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n662_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n661_), .B1(new_n663_), .B2(new_n664_), .ZN(G1326gat));
  INV_X1    g464(.A(G22gat), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n660_), .A2(new_n666_), .A3(new_n378_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n641_), .A2(new_n378_), .A3(new_n644_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(G22gat), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n669_), .A2(KEYINPUT42), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n669_), .A2(KEYINPUT42), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n667_), .B1(new_n670_), .B2(new_n671_), .ZN(G1327gat));
  NOR2_X1   g471(.A1(new_n628_), .A2(new_n637_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(new_n609_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n674_), .B1(new_n482_), .B2(new_n495_), .ZN(new_n675_));
  AOI21_X1  g474(.A(G29gat), .B1(new_n675_), .B2(new_n342_), .ZN(new_n676_));
  OAI21_X1  g475(.A(KEYINPUT43), .B1(new_n414_), .B2(new_n572_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT43), .ZN(new_n678_));
  INV_X1    g477(.A(new_n572_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n485_), .A2(new_n678_), .A3(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n677_), .A2(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(KEYINPUT105), .B1(new_n642_), .B2(new_n628_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT105), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n643_), .A2(new_n683_), .A3(new_n494_), .A4(new_n609_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(KEYINPUT44), .B1(new_n681_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687_));
  INV_X1    g486(.A(new_n685_), .ZN(new_n688_));
  AOI211_X1 g487(.A(new_n687_), .B(new_n688_), .C1(new_n677_), .C2(new_n680_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n686_), .A2(new_n689_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n343_), .A2(new_n441_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n676_), .B1(new_n690_), .B2(new_n691_), .ZN(G1328gat));
  INV_X1    g491(.A(KEYINPUT46), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(KEYINPUT107), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n693_), .A2(KEYINPUT107), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n439_), .B1(new_n690_), .B2(new_n651_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n651_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(KEYINPUT106), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT106), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n651_), .A2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n698_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n702_), .A2(G36gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(KEYINPUT45), .B1(new_n675_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n675_), .A2(KEYINPUT45), .A3(new_n703_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n694_), .B(new_n695_), .C1(new_n696_), .C2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n681_), .A2(new_n685_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(new_n687_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n681_), .A2(KEYINPUT44), .A3(new_n685_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(G36gat), .B1(new_n712_), .B2(new_n697_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n705_), .A2(new_n706_), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n713_), .A2(new_n714_), .A3(KEYINPUT107), .A4(new_n693_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n708_), .A2(new_n715_), .ZN(G1329gat));
  INV_X1    g515(.A(new_n675_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n405_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n405_), .A2(G43gat), .ZN(new_n720_));
  OAI22_X1  g519(.A1(G43gat), .A2(new_n719_), .B1(new_n712_), .B2(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n721_), .B(new_n723_), .ZN(G1330gat));
  OAI21_X1  g523(.A(G50gat), .B1(new_n712_), .B2(new_n377_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n377_), .A2(G50gat), .ZN(new_n726_));
  XOR2_X1   g525(.A(new_n726_), .B(KEYINPUT109), .Z(new_n727_));
  OAI21_X1  g526(.A(new_n725_), .B1(new_n717_), .B2(new_n727_), .ZN(G1331gat));
  NOR2_X1   g527(.A1(new_n414_), .A2(new_n494_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n609_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n729_), .A2(new_n730_), .A3(new_n631_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(G57gat), .B1(new_n732_), .B2(new_n342_), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n643_), .A2(new_n494_), .A3(new_n609_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n735_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n343_), .A2(KEYINPUT110), .ZN(new_n737_));
  MUX2_X1   g536(.A(KEYINPUT110), .B(new_n737_), .S(G57gat), .Z(new_n738_));
  AOI21_X1  g537(.A(new_n733_), .B1(new_n736_), .B2(new_n738_), .ZN(G1332gat));
  OR3_X1    g538(.A1(new_n731_), .A2(G64gat), .A3(new_n702_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n736_), .A2(new_n701_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(G64gat), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n742_), .A2(KEYINPUT48), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n742_), .A2(KEYINPUT48), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n740_), .B1(new_n743_), .B2(new_n744_), .ZN(G1333gat));
  NAND3_X1  g544(.A1(new_n732_), .A2(new_n382_), .A3(new_n405_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n736_), .A2(new_n405_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(G71gat), .ZN(new_n748_));
  OR2_X1    g547(.A1(new_n748_), .A2(KEYINPUT112), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(KEYINPUT112), .ZN(new_n750_));
  XOR2_X1   g549(.A(KEYINPUT111), .B(KEYINPUT49), .Z(new_n751_));
  AND3_X1   g550(.A1(new_n749_), .A2(new_n750_), .A3(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n746_), .B1(new_n752_), .B2(new_n753_), .ZN(G1334gat));
  NOR2_X1   g553(.A1(new_n377_), .A2(G78gat), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT113), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n732_), .A2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT50), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n736_), .A2(new_n378_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n758_), .B1(new_n759_), .B2(G78gat), .ZN(new_n760_));
  AOI211_X1 g559(.A(KEYINPUT50), .B(new_n582_), .C1(new_n736_), .C2(new_n378_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n757_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT114), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n762_), .B(new_n763_), .ZN(G1335gat));
  NOR3_X1   g563(.A1(new_n628_), .A2(new_n609_), .A3(new_n637_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n729_), .A2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(G85gat), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n767_), .A2(new_n768_), .A3(new_n342_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n643_), .A2(new_n730_), .A3(new_n481_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT116), .ZN(new_n771_));
  OR2_X1    g570(.A1(new_n681_), .A2(KEYINPUT115), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n681_), .A2(KEYINPUT115), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n771_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n774_), .A2(new_n342_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n769_), .B1(new_n775_), .B2(new_n768_), .ZN(G1336gat));
  AOI21_X1  g575(.A(G92gat), .B1(new_n767_), .B2(new_n651_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n701_), .A2(new_n510_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n777_), .B1(new_n774_), .B2(new_n778_), .ZN(G1337gat));
  INV_X1    g578(.A(KEYINPUT51), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n767_), .A2(new_n405_), .A3(new_n502_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n774_), .A2(new_n405_), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n780_), .B(new_n781_), .C1(new_n782_), .C2(new_n521_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n521_), .B1(new_n774_), .B2(new_n405_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n781_), .ZN(new_n785_));
  OAI21_X1  g584(.A(KEYINPUT51), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n783_), .A2(new_n786_), .ZN(G1338gat));
  NAND3_X1  g586(.A1(new_n767_), .A2(new_n503_), .A3(new_n378_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n681_), .ZN(new_n789_));
  OR2_X1    g588(.A1(new_n771_), .A2(new_n377_), .ZN(new_n790_));
  OAI21_X1  g589(.A(G106gat), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n791_), .A2(KEYINPUT52), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n791_), .A2(KEYINPUT52), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n788_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(KEYINPUT53), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n796_), .B(new_n788_), .C1(new_n792_), .C2(new_n793_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n797_), .ZN(G1339gat));
  INV_X1    g597(.A(KEYINPUT54), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n631_), .A2(new_n799_), .A3(new_n481_), .A4(new_n609_), .ZN(new_n800_));
  OAI21_X1  g599(.A(KEYINPUT54), .B1(new_n629_), .B2(new_n494_), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n592_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n595_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n602_), .A2(new_n805_), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n597_), .B(KEYINPUT55), .C1(new_n600_), .C2(new_n601_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n804_), .A2(new_n806_), .A3(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n578_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT118), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT117), .B1(new_n811_), .B2(KEYINPUT56), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n810_), .A2(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n602_), .A2(new_n605_), .A3(new_n578_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n494_), .A2(new_n814_), .A3(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n808_), .A2(new_n817_), .A3(new_n809_), .ZN(new_n818_));
  AOI21_X1  g617(.A(KEYINPUT56), .B1(new_n818_), .B2(new_n811_), .ZN(new_n819_));
  OAI21_X1  g618(.A(KEYINPUT119), .B1(new_n816_), .B2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n811_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT56), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n815_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n481_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT119), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n823_), .A2(new_n825_), .A3(new_n826_), .A4(new_n814_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n465_), .B1(new_n469_), .B2(new_n474_), .ZN(new_n828_));
  NOR3_X1   g627(.A1(new_n461_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n418_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n417_), .B1(new_n479_), .B2(new_n466_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  OR2_X1    g631(.A1(new_n832_), .A2(new_n607_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n820_), .A2(new_n827_), .A3(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n637_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(KEYINPUT120), .A2(KEYINPUT57), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT121), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n824_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n808_), .A2(new_n822_), .A3(new_n809_), .ZN(new_n840_));
  AND2_X1   g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n810_), .A2(KEYINPUT56), .ZN(new_n842_));
  AOI21_X1  g641(.A(KEYINPUT58), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n838_), .B1(new_n572_), .B2(new_n843_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n842_), .A2(KEYINPUT58), .A3(new_n840_), .A4(new_n839_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT122), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n845_), .B(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT58), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n839_), .A2(new_n840_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n822_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n848_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n851_), .B(KEYINPUT121), .C1(new_n570_), .C2(new_n571_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n844_), .A2(new_n847_), .A3(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n836_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n834_), .A2(new_n637_), .A3(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n837_), .A2(new_n853_), .A3(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n802_), .B1(new_n856_), .B2(new_n643_), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n651_), .A2(new_n411_), .A3(new_n343_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n857_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(G113gat), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(new_n861_), .A3(new_n494_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT59), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n863_), .B1(new_n857_), .B2(new_n859_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n855_), .A2(new_n853_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n628_), .B1(new_n865_), .B2(new_n837_), .ZN(new_n866_));
  OAI211_X1 g665(.A(KEYINPUT59), .B(new_n858_), .C1(new_n866_), .C2(new_n802_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n481_), .B1(new_n864_), .B2(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n862_), .B1(new_n868_), .B2(new_n861_), .ZN(G1340gat));
  INV_X1    g668(.A(KEYINPUT123), .ZN(new_n870_));
  INV_X1    g669(.A(G120gat), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n864_), .A2(new_n867_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n871_), .B1(new_n872_), .B2(new_n730_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n860_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n871_), .B1(new_n609_), .B2(KEYINPUT60), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n875_), .B1(KEYINPUT60), .B2(new_n871_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n874_), .A2(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n870_), .B1(new_n873_), .B2(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n609_), .B1(new_n864_), .B2(new_n867_), .ZN(new_n879_));
  OAI221_X1 g678(.A(KEYINPUT123), .B1(new_n874_), .B2(new_n876_), .C1(new_n879_), .C2(new_n871_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n878_), .A2(new_n880_), .ZN(G1341gat));
  INV_X1    g680(.A(G127gat), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n882_), .B1(new_n872_), .B2(new_n628_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n628_), .A2(new_n882_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n874_), .A2(new_n884_), .ZN(new_n885_));
  OAI21_X1  g684(.A(KEYINPUT124), .B1(new_n883_), .B2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT124), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n643_), .B1(new_n864_), .B2(new_n867_), .ZN(new_n888_));
  OAI221_X1 g687(.A(new_n887_), .B1(new_n874_), .B2(new_n884_), .C1(new_n888_), .C2(new_n882_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n886_), .A2(new_n889_), .ZN(G1342gat));
  AOI21_X1  g689(.A(G134gat), .B1(new_n860_), .B2(new_n638_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT125), .ZN(new_n892_));
  OR2_X1    g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n891_), .A2(new_n892_), .ZN(new_n894_));
  AND2_X1   g693(.A1(new_n679_), .A2(G134gat), .ZN(new_n895_));
  AOI22_X1  g694(.A1(new_n893_), .A2(new_n894_), .B1(new_n872_), .B2(new_n895_), .ZN(G1343gat));
  NOR4_X1   g695(.A1(new_n857_), .A2(new_n412_), .A3(new_n343_), .A4(new_n701_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n494_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g698(.A1(new_n897_), .A2(new_n730_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g700(.A1(new_n897_), .A2(new_n628_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(KEYINPUT61), .B(G155gat), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n902_), .B(new_n903_), .ZN(G1346gat));
  INV_X1    g703(.A(G162gat), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n897_), .A2(new_n905_), .A3(new_n638_), .ZN(new_n906_));
  AND2_X1   g705(.A1(new_n897_), .A2(new_n679_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n907_), .B2(new_n905_), .ZN(G1347gat));
  INV_X1    g707(.A(KEYINPUT62), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n701_), .A2(new_n343_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n910_), .A2(new_n411_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n857_), .A2(new_n912_), .A3(new_n481_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(KEYINPUT126), .ZN(new_n914_));
  INV_X1    g713(.A(new_n914_), .ZN(new_n915_));
  OAI21_X1  g714(.A(G169gat), .B1(new_n913_), .B2(KEYINPUT126), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n909_), .B1(new_n915_), .B2(new_n916_), .ZN(new_n917_));
  OR2_X1    g716(.A1(new_n913_), .A2(KEYINPUT126), .ZN(new_n918_));
  NAND4_X1  g717(.A1(new_n918_), .A2(KEYINPUT62), .A3(new_n914_), .A4(G169gat), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n913_), .A2(new_n230_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n917_), .A2(new_n919_), .A3(new_n920_), .ZN(G1348gat));
  NOR2_X1   g720(.A1(new_n857_), .A2(new_n912_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(new_n730_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n923_), .A2(new_n254_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n924_), .B1(new_n231_), .B2(new_n923_), .ZN(G1349gat));
  NAND2_X1  g724(.A1(new_n922_), .A2(new_n628_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n926_), .A2(new_n248_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n927_), .B1(new_n235_), .B2(new_n926_), .ZN(G1350gat));
  INV_X1    g727(.A(new_n922_), .ZN(new_n929_));
  OAI21_X1  g728(.A(G190gat), .B1(new_n929_), .B2(new_n572_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n922_), .A2(new_n249_), .A3(new_n638_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(G1351gat));
  NOR3_X1   g731(.A1(new_n857_), .A2(new_n412_), .A3(new_n910_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(new_n494_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n934_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g734(.A1(new_n857_), .A2(new_n412_), .ZN(new_n936_));
  INV_X1    g735(.A(new_n910_), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n936_), .A2(new_n730_), .A3(new_n937_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n938_), .A2(new_n216_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n933_), .A2(new_n209_), .A3(new_n730_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n939_), .A2(new_n940_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n941_), .A2(KEYINPUT127), .ZN(new_n942_));
  INV_X1    g741(.A(KEYINPUT127), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n939_), .A2(new_n940_), .A3(new_n943_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n942_), .A2(new_n944_), .ZN(G1353gat));
  NAND2_X1  g744(.A1(new_n933_), .A2(new_n628_), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n946_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n947_));
  XOR2_X1   g746(.A(KEYINPUT63), .B(G211gat), .Z(new_n948_));
  OAI21_X1  g747(.A(new_n947_), .B1(new_n946_), .B2(new_n948_), .ZN(G1354gat));
  INV_X1    g748(.A(G218gat), .ZN(new_n950_));
  NAND3_X1  g749(.A1(new_n933_), .A2(new_n950_), .A3(new_n638_), .ZN(new_n951_));
  AND2_X1   g750(.A1(new_n933_), .A2(new_n679_), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n951_), .B1(new_n952_), .B2(new_n950_), .ZN(G1355gat));
endmodule


