//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 1 1 1 1 1 1 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n786_, new_n787_, new_n788_, new_n790_, new_n791_,
    new_n792_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n903_, new_n904_, new_n905_,
    new_n907_, new_n908_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n919_, new_n920_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n942_, new_n943_, new_n945_, new_n946_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n953_, new_n954_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n968_, new_n969_, new_n970_,
    new_n971_, new_n972_, new_n973_;
  XNOR2_X1  g000(.A(G211gat), .B(G218gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT95), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT21), .ZN(new_n205_));
  INV_X1    g004(.A(G197gat), .ZN(new_n206_));
  OR2_X1    g005(.A1(KEYINPUT94), .A2(G204gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(KEYINPUT94), .A2(G204gat), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n206_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(G197gat), .A2(G204gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n205_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n207_), .A2(new_n206_), .A3(new_n208_), .ZN(new_n212_));
  INV_X1    g011(.A(G204gat), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n212_), .B(KEYINPUT21), .C1(new_n206_), .C2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n204_), .A2(new_n211_), .A3(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n202_), .B(KEYINPUT95), .ZN(new_n216_));
  NOR3_X1   g015(.A1(new_n209_), .A2(new_n205_), .A3(new_n210_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n215_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(G183gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT85), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT85), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(G183gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n221_), .A2(new_n223_), .A3(KEYINPUT25), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT86), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT85), .B(G183gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n227_), .A2(KEYINPUT86), .A3(KEYINPUT25), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT25), .ZN(new_n229_));
  AND2_X1   g028(.A1(new_n229_), .A2(KEYINPUT87), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n229_), .A2(KEYINPUT87), .ZN(new_n231_));
  OAI21_X1  g030(.A(G183gat), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT26), .B(G190gat), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n226_), .A2(new_n228_), .A3(new_n232_), .A4(new_n233_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(G169gat), .A2(G176gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(KEYINPUT88), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT88), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n237_), .B1(G169gat), .B2(G176gat), .ZN(new_n238_));
  AOI21_X1  g037(.A(KEYINPUT24), .B1(new_n236_), .B2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G183gat), .A2(G190gat), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT23), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n239_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n236_), .A2(new_n238_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT24), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n246_), .B1(G169gat), .B2(G176gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n234_), .A2(new_n243_), .A3(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT90), .ZN(new_n250_));
  INV_X1    g049(.A(G169gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT22), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT22), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(G169gat), .ZN(new_n254_));
  INV_X1    g053(.A(G176gat), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n252_), .A2(new_n254_), .A3(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT89), .ZN(new_n257_));
  INV_X1    g056(.A(G190gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n227_), .A2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n240_), .B(KEYINPUT23), .ZN(new_n260_));
  AOI22_X1  g059(.A1(new_n259_), .A2(new_n260_), .B1(G169gat), .B2(G176gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n257_), .A2(new_n261_), .ZN(new_n262_));
  AND3_X1   g061(.A1(new_n249_), .A2(new_n250_), .A3(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n250_), .B1(new_n249_), .B2(new_n262_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n219_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G226gat), .A2(G233gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT19), .ZN(new_n267_));
  OAI211_X1 g066(.A(KEYINPUT99), .B(new_n260_), .C1(new_n245_), .C2(KEYINPUT24), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT99), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n269_), .B1(new_n239_), .B2(new_n242_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n268_), .A2(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(KEYINPUT25), .B(G183gat), .ZN(new_n272_));
  AOI22_X1  g071(.A1(new_n245_), .A2(new_n247_), .B1(new_n233_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n252_), .A2(new_n254_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT100), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(new_n255_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n220_), .A2(new_n258_), .ZN(new_n277_));
  AOI22_X1  g076(.A1(new_n260_), .A2(new_n277_), .B1(G169gat), .B2(G176gat), .ZN(new_n278_));
  AOI22_X1  g077(.A1(new_n271_), .A2(new_n273_), .B1(new_n276_), .B2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n219_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n267_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n265_), .A2(KEYINPUT20), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT101), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NOR3_X1   g083(.A1(new_n263_), .A2(new_n264_), .A3(new_n219_), .ZN(new_n285_));
  OAI21_X1  g084(.A(KEYINPUT20), .B1(new_n279_), .B2(new_n280_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n267_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n265_), .A2(new_n281_), .A3(KEYINPUT101), .A4(KEYINPUT20), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n284_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  XOR2_X1   g088(.A(G8gat), .B(G36gat), .Z(new_n290_));
  XNOR2_X1  g089(.A(G64gat), .B(G92gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT102), .B(KEYINPUT18), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n289_), .A2(new_n295_), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n284_), .A2(new_n287_), .A3(new_n294_), .A4(new_n288_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT27), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT96), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n219_), .A2(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n215_), .A2(new_n218_), .A3(KEYINPUT96), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n301_), .A2(new_n279_), .A3(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n265_), .A2(KEYINPUT20), .A3(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(new_n267_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n279_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(new_n219_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n264_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n249_), .A2(new_n250_), .A3(new_n262_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  OAI211_X1 g109(.A(new_n307_), .B(KEYINPUT20), .C1(new_n310_), .C2(new_n219_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n305_), .B1(new_n267_), .B2(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n299_), .B1(new_n312_), .B2(new_n295_), .ZN(new_n313_));
  AOI22_X1  g112(.A1(new_n298_), .A2(new_n299_), .B1(new_n313_), .B2(new_n297_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT3), .ZN(new_n315_));
  INV_X1    g114(.A(G141gat), .ZN(new_n316_));
  INV_X1    g115(.A(G148gat), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n315_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G141gat), .A2(G148gat), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT2), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n322_));
  OAI21_X1  g121(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n318_), .A2(new_n321_), .A3(new_n322_), .A4(new_n323_), .ZN(new_n324_));
  OR2_X1    g123(.A1(G155gat), .A2(G162gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G155gat), .A2(G162gat), .ZN(new_n326_));
  AND2_X1   g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n324_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(KEYINPUT1), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT1), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n330_), .A2(G155gat), .A3(G162gat), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n329_), .A2(new_n331_), .A3(new_n325_), .ZN(new_n332_));
  XOR2_X1   g131(.A(G141gat), .B(G148gat), .Z(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n328_), .A2(new_n334_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n335_), .A2(KEYINPUT29), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT28), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G22gat), .B(G50gat), .ZN(new_n338_));
  AND2_X1   g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n337_), .A2(new_n338_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(G228gat), .ZN(new_n342_));
  INV_X1    g141(.A(G233gat), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n335_), .A2(KEYINPUT29), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n219_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n347_));
  AOI22_X1  g146(.A1(new_n301_), .A2(new_n302_), .B1(KEYINPUT29), .B2(new_n335_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n347_), .B1(new_n348_), .B2(new_n345_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G78gat), .B(G106gat), .ZN(new_n350_));
  XOR2_X1   g149(.A(new_n350_), .B(KEYINPUT97), .Z(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n349_), .A2(new_n352_), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n351_), .B(new_n347_), .C1(new_n348_), .C2(new_n345_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n341_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n341_), .A2(new_n354_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n350_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n301_), .A2(new_n302_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(new_n346_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(new_n344_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n357_), .B1(new_n360_), .B2(new_n347_), .ZN(new_n361_));
  OAI21_X1  g160(.A(KEYINPUT98), .B1(new_n356_), .B2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n349_), .A2(new_n350_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT98), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n363_), .A2(new_n364_), .A3(new_n341_), .A4(new_n354_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n355_), .B1(new_n362_), .B2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G71gat), .B(G99gat), .ZN(new_n367_));
  INV_X1    g166(.A(G43gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n310_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n369_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n308_), .A2(new_n309_), .A3(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n370_), .A2(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G127gat), .B(G134gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G113gat), .B(G120gat), .ZN(new_n375_));
  AND2_X1   g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n374_), .A2(new_n375_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n373_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n378_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n370_), .A2(new_n380_), .A3(new_n372_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n379_), .A2(new_n381_), .ZN(new_n382_));
  XOR2_X1   g181(.A(KEYINPUT92), .B(G15gat), .Z(new_n383_));
  NAND2_X1  g182(.A1(G227gat), .A2(G233gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT91), .B(KEYINPUT30), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT93), .B(KEYINPUT31), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n382_), .A2(new_n390_), .ZN(new_n391_));
  OAI22_X1  g190(.A1(new_n335_), .A2(KEYINPUT103), .B1(new_n376_), .B2(new_n377_), .ZN(new_n392_));
  AOI22_X1  g191(.A1(new_n324_), .A2(new_n327_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT103), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n378_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n392_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(KEYINPUT4), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G225gat), .A2(G233gat), .ZN(new_n398_));
  XOR2_X1   g197(.A(new_n398_), .B(KEYINPUT104), .Z(new_n399_));
  OR3_X1    g198(.A1(new_n380_), .A2(KEYINPUT4), .A3(new_n393_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n397_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G1gat), .B(G29gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(G85gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT0), .B(G57gat), .ZN(new_n404_));
  XOR2_X1   g203(.A(new_n403_), .B(new_n404_), .Z(new_n405_));
  INV_X1    g204(.A(new_n399_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n396_), .A2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n401_), .A2(new_n405_), .A3(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n405_), .B1(new_n401_), .B2(new_n407_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n379_), .A2(new_n381_), .A3(new_n389_), .ZN(new_n412_));
  AND3_X1   g211(.A1(new_n391_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n413_));
  AND3_X1   g212(.A1(new_n314_), .A2(new_n366_), .A3(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n411_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n362_), .A2(new_n365_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n355_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n415_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n314_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT105), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT33), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n408_), .A2(new_n420_), .A3(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n396_), .A2(new_n399_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n405_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT106), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n423_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n397_), .A2(new_n406_), .A3(new_n400_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n406_), .B1(new_n392_), .B2(new_n395_), .ZN(new_n428_));
  OAI21_X1  g227(.A(KEYINPUT106), .B1(new_n428_), .B2(new_n405_), .ZN(new_n429_));
  AND3_X1   g228(.A1(new_n426_), .A2(new_n427_), .A3(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n408_), .A2(new_n420_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n430_), .B1(new_n431_), .B2(KEYINPUT33), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n296_), .A2(new_n297_), .A3(new_n422_), .A4(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n294_), .A2(KEYINPUT32), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n312_), .A2(new_n435_), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n284_), .A2(new_n287_), .A3(new_n434_), .A4(new_n288_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n436_), .A2(new_n415_), .A3(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n433_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(new_n366_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n419_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n391_), .A2(new_n412_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n414_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  XOR2_X1   g242(.A(KEYINPUT70), .B(G71gat), .Z(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(G78gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(KEYINPUT70), .B(G71gat), .ZN(new_n446_));
  INV_X1    g245(.A(G78gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G57gat), .B(G64gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT11), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n449_), .A2(KEYINPUT11), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n445_), .B(new_n448_), .C1(new_n451_), .C2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n448_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n446_), .A2(new_n447_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n450_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT71), .ZN(new_n457_));
  AND3_X1   g256(.A1(new_n453_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n457_), .B1(new_n453_), .B2(new_n456_), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT12), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  XOR2_X1   g259(.A(G85gat), .B(G92gat), .Z(new_n461_));
  XOR2_X1   g260(.A(KEYINPUT66), .B(G92gat), .Z(new_n462_));
  INV_X1    g261(.A(G85gat), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n463_), .A2(KEYINPUT9), .ZN(new_n464_));
  AOI22_X1  g263(.A1(KEYINPUT9), .A2(new_n461_), .B1(new_n462_), .B2(new_n464_), .ZN(new_n465_));
  AND3_X1   g264(.A1(KEYINPUT67), .A2(G99gat), .A3(G106gat), .ZN(new_n466_));
  AOI21_X1  g265(.A(KEYINPUT67), .B1(G99gat), .B2(G106gat), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT6), .ZN(new_n468_));
  NOR3_X1   g267(.A1(new_n466_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G99gat), .A2(G106gat), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT67), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(KEYINPUT67), .A2(G99gat), .A3(G106gat), .ZN(new_n473_));
  AOI21_X1  g272(.A(KEYINPUT6), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n469_), .A2(new_n474_), .ZN(new_n475_));
  XOR2_X1   g274(.A(KEYINPUT10), .B(G99gat), .Z(new_n476_));
  INV_X1    g275(.A(G106gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n465_), .A2(new_n475_), .A3(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT8), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT68), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n481_), .A2(KEYINPUT6), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n468_), .A2(KEYINPUT68), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n472_), .B(new_n473_), .C1(new_n482_), .C2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT7), .ZN(new_n485_));
  INV_X1    g284(.A(G99gat), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n485_), .A2(new_n486_), .A3(new_n477_), .ZN(new_n487_));
  OAI21_X1  g286(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n488_));
  AND2_X1   g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n468_), .A2(KEYINPUT68), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n481_), .A2(KEYINPUT6), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n490_), .B(new_n491_), .C1(new_n466_), .C2(new_n467_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n484_), .A2(new_n489_), .A3(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n480_), .B1(new_n493_), .B2(new_n461_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n461_), .A2(new_n480_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n495_), .B1(new_n475_), .B2(new_n489_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n479_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n460_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n453_), .A2(new_n456_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n466_), .A2(new_n467_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(KEYINPUT6), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n468_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n502_), .A2(new_n489_), .A3(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n495_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n461_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n487_), .A2(new_n488_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n490_), .A2(new_n491_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n508_), .B1(new_n501_), .B2(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n507_), .B1(new_n510_), .B2(new_n492_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n506_), .B1(new_n511_), .B2(new_n480_), .ZN(new_n512_));
  AOI21_X1  g311(.A(KEYINPUT69), .B1(new_n512_), .B2(new_n479_), .ZN(new_n513_));
  OAI211_X1 g312(.A(KEYINPUT69), .B(new_n479_), .C1(new_n494_), .C2(new_n496_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n500_), .B1(new_n513_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT12), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n499_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT69), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n497_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n500_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n520_), .A2(new_n521_), .A3(new_n514_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G230gat), .A2(G233gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n523_), .B(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n522_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n516_), .A2(new_n522_), .ZN(new_n528_));
  AOI22_X1  g327(.A1(new_n518_), .A2(new_n527_), .B1(new_n528_), .B2(new_n525_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT73), .ZN(new_n530_));
  XOR2_X1   g329(.A(G120gat), .B(G148gat), .Z(new_n531_));
  XNOR2_X1  g330(.A(G176gat), .B(G204gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n533_), .B(new_n534_), .Z(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n529_), .A2(new_n530_), .A3(new_n536_), .ZN(new_n537_));
  AND3_X1   g336(.A1(new_n520_), .A2(new_n521_), .A3(new_n514_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n521_), .B1(new_n520_), .B2(new_n514_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n525_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n459_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n453_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n543_), .A2(KEYINPUT12), .A3(new_n497_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n544_), .B1(new_n539_), .B2(KEYINPUT12), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n522_), .A2(new_n526_), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n540_), .B(new_n536_), .C1(new_n545_), .C2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(KEYINPUT73), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n537_), .A2(new_n548_), .ZN(new_n549_));
  OR2_X1    g348(.A1(new_n529_), .A2(new_n536_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT13), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n549_), .A2(KEYINPUT13), .A3(new_n550_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT15), .ZN(new_n556_));
  INV_X1    g355(.A(G36gat), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(G29gat), .ZN(new_n558_));
  INV_X1    g357(.A(G29gat), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(G36gat), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT74), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n558_), .A2(new_n560_), .A3(KEYINPUT74), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G43gat), .B(G50gat), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n563_), .A2(new_n564_), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n565_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n556_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n568_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n570_), .A2(KEYINPUT15), .A3(new_n566_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G15gat), .B(G22gat), .ZN(new_n573_));
  INV_X1    g372(.A(G1gat), .ZN(new_n574_));
  INV_X1    g373(.A(G8gat), .ZN(new_n575_));
  OAI21_X1  g374(.A(KEYINPUT14), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n573_), .A2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G1gat), .B(G8gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n572_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n579_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n567_), .A2(new_n568_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(G229gat), .A2(G233gat), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n580_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n579_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n583_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n584_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n585_), .A2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G113gat), .B(G141gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G169gat), .B(G197gat), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n591_), .B(new_n592_), .Z(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n590_), .B1(KEYINPUT83), .B2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(KEYINPUT83), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n596_), .B1(new_n585_), .B2(new_n589_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  OR2_X1    g397(.A1(new_n598_), .A2(KEYINPUT84), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(KEYINPUT84), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NOR3_X1   g401(.A1(new_n443_), .A2(new_n555_), .A3(new_n602_), .ZN(new_n603_));
  XOR2_X1   g402(.A(G127gat), .B(G155gat), .Z(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT16), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G183gat), .B(G211gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT17), .ZN(new_n608_));
  AND2_X1   g407(.A1(G231gat), .A2(G233gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n579_), .B(new_n609_), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n610_), .A2(new_n521_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n521_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n608_), .A2(new_n611_), .A3(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT82), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT17), .ZN(new_n615_));
  AOI211_X1 g414(.A(new_n615_), .B(new_n607_), .C1(new_n543_), .C2(new_n610_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n616_), .B1(new_n543_), .B2(new_n610_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n614_), .A2(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n520_), .A2(new_n582_), .A3(new_n514_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(KEYINPUT77), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT77), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n520_), .A2(new_n621_), .A3(new_n582_), .A4(new_n514_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT76), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT75), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n572_), .A2(new_n625_), .A3(new_n497_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n625_), .B1(new_n572_), .B2(new_n497_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n624_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n628_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n630_), .A2(KEYINPUT76), .A3(new_n626_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n623_), .A2(new_n629_), .A3(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(G232gat), .A2(G233gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT34), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT35), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n632_), .A2(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(G190gat), .B(G218gat), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT78), .ZN(new_n639_));
  XNOR2_X1  g438(.A(G134gat), .B(G162gat), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n639_), .B(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n642_), .A2(KEYINPUT36), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n634_), .A2(KEYINPUT35), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n644_), .B1(KEYINPUT79), .B2(new_n635_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n645_), .B1(KEYINPUT79), .B2(new_n635_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n646_), .B1(new_n630_), .B2(new_n626_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n623_), .A2(KEYINPUT80), .A3(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(KEYINPUT80), .B1(new_n623_), .B2(new_n647_), .ZN(new_n650_));
  OAI211_X1 g449(.A(new_n637_), .B(new_n643_), .C1(new_n649_), .C2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n623_), .A2(new_n647_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT80), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  AOI22_X1  g453(.A1(new_n654_), .A2(new_n648_), .B1(new_n636_), .B2(new_n632_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n641_), .B(KEYINPUT36), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n656_), .B(KEYINPUT81), .Z(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n651_), .B1(new_n655_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT37), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  OAI211_X1 g460(.A(new_n651_), .B(KEYINPUT37), .C1(new_n655_), .C2(new_n658_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  AND3_X1   g463(.A1(new_n603_), .A2(new_n618_), .A3(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n665_), .A2(new_n574_), .A3(new_n415_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT38), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n314_), .A2(new_n366_), .A3(new_n413_), .ZN(new_n668_));
  AOI22_X1  g467(.A1(new_n418_), .A2(new_n314_), .B1(new_n439_), .B2(new_n366_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n442_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n668_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n671_), .A2(new_n618_), .A3(new_n659_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n598_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n553_), .A2(new_n673_), .A3(new_n554_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(KEYINPUT107), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT107), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n553_), .A2(new_n676_), .A3(new_n673_), .A4(new_n554_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n672_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(G1gat), .B1(new_n680_), .B2(new_n411_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n667_), .A2(new_n681_), .ZN(G1324gat));
  INV_X1    g481(.A(new_n314_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n665_), .A2(new_n575_), .A3(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT39), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n679_), .A2(new_n683_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n685_), .B1(new_n686_), .B2(G8gat), .ZN(new_n687_));
  AOI211_X1 g486(.A(KEYINPUT39), .B(new_n575_), .C1(new_n679_), .C2(new_n683_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n684_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n691_), .ZN(new_n692_));
  OAI211_X1 g491(.A(new_n684_), .B(new_n690_), .C1(new_n687_), .C2(new_n688_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1325gat));
  INV_X1    g493(.A(G15gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n695_), .B1(new_n679_), .B2(new_n670_), .ZN(new_n696_));
  XOR2_X1   g495(.A(KEYINPUT109), .B(KEYINPUT41), .Z(new_n697_));
  OR2_X1    g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n665_), .A2(new_n695_), .A3(new_n670_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n696_), .A2(new_n697_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n698_), .A2(new_n699_), .A3(new_n700_), .ZN(G1326gat));
  INV_X1    g500(.A(G22gat), .ZN(new_n702_));
  INV_X1    g501(.A(new_n366_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n665_), .A2(new_n702_), .A3(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT42), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n679_), .A2(new_n703_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n705_), .B1(new_n706_), .B2(G22gat), .ZN(new_n707_));
  AOI211_X1 g506(.A(KEYINPUT42), .B(new_n702_), .C1(new_n679_), .C2(new_n703_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n704_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT110), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  OAI211_X1 g510(.A(KEYINPUT110), .B(new_n704_), .C1(new_n707_), .C2(new_n708_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(G1327gat));
  INV_X1    g512(.A(new_n618_), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n675_), .A2(new_n677_), .A3(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT43), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n670_), .B1(new_n419_), .B2(new_n440_), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n716_), .B(new_n663_), .C1(new_n717_), .C2(new_n414_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n716_), .B1(new_n671_), .B2(new_n663_), .ZN(new_n720_));
  OAI211_X1 g519(.A(KEYINPUT44), .B(new_n715_), .C1(new_n719_), .C2(new_n720_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n675_), .A2(new_n677_), .A3(new_n714_), .ZN(new_n722_));
  OAI21_X1  g521(.A(KEYINPUT43), .B1(new_n443_), .B2(new_n664_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n722_), .B1(new_n723_), .B2(new_n718_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(KEYINPUT111), .B(KEYINPUT44), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n721_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n726_));
  OR3_X1    g525(.A1(new_n726_), .A2(new_n559_), .A3(new_n411_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n659_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(new_n714_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n603_), .A2(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n559_), .B1(new_n731_), .B2(new_n411_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n727_), .A2(new_n732_), .ZN(G1328gat));
  OAI211_X1 g532(.A(new_n721_), .B(new_n683_), .C1(new_n724_), .C2(new_n725_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(G36gat), .ZN(new_n735_));
  NAND4_X1  g534(.A1(new_n603_), .A2(new_n557_), .A3(new_n683_), .A4(new_n730_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT45), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT46), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n735_), .A2(new_n737_), .A3(KEYINPUT46), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(G1329gat));
  OAI21_X1  g541(.A(new_n368_), .B1(new_n731_), .B2(new_n442_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n670_), .A2(G43gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n743_), .B1(new_n726_), .B2(new_n744_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g545(.A1(new_n703_), .A2(G50gat), .ZN(new_n747_));
  OR2_X1    g546(.A1(new_n726_), .A2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(G50gat), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n749_), .B1(new_n731_), .B2(new_n366_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n748_), .A2(new_n750_), .ZN(G1331gat));
  NAND3_X1  g550(.A1(new_n671_), .A2(new_n598_), .A3(new_n555_), .ZN(new_n752_));
  NOR3_X1   g551(.A1(new_n752_), .A2(new_n714_), .A3(new_n663_), .ZN(new_n753_));
  INV_X1    g552(.A(G57gat), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n753_), .A2(new_n754_), .A3(new_n415_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n443_), .A2(new_n728_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n601_), .A2(new_n714_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n555_), .A2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(G57gat), .B1(new_n759_), .B2(new_n411_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n755_), .A2(new_n760_), .ZN(G1332gat));
  OAI21_X1  g560(.A(G64gat), .B1(new_n759_), .B2(new_n314_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT48), .ZN(new_n763_));
  INV_X1    g562(.A(G64gat), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n753_), .A2(new_n764_), .A3(new_n683_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n763_), .A2(new_n765_), .ZN(G1333gat));
  OAI21_X1  g565(.A(G71gat), .B1(new_n759_), .B2(new_n442_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT49), .ZN(new_n768_));
  INV_X1    g567(.A(G71gat), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n753_), .A2(new_n769_), .A3(new_n670_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(G1334gat));
  NAND3_X1  g570(.A1(new_n753_), .A2(new_n447_), .A3(new_n703_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n759_), .A2(new_n366_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n773_), .A2(new_n447_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n774_), .A2(new_n775_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n772_), .B1(new_n776_), .B2(new_n777_), .ZN(G1335gat));
  INV_X1    g577(.A(new_n555_), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n779_), .A2(new_n673_), .A3(new_n618_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n780_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n781_));
  OAI21_X1  g580(.A(G85gat), .B1(new_n781_), .B2(new_n411_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n752_), .A2(new_n729_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n783_), .A2(new_n463_), .A3(new_n415_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(G1336gat));
  AOI21_X1  g584(.A(G92gat), .B1(new_n783_), .B2(new_n683_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n781_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n683_), .A2(new_n462_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n786_), .B1(new_n787_), .B2(new_n788_), .ZN(G1337gat));
  NAND3_X1  g588(.A1(new_n783_), .A2(new_n476_), .A3(new_n670_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n781_), .A2(new_n442_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n790_), .B1(new_n791_), .B2(new_n486_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n792_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g592(.A1(new_n783_), .A2(new_n477_), .A3(new_n703_), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n703_), .B(new_n780_), .C1(new_n719_), .C2(new_n720_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n795_), .A2(new_n796_), .A3(G106gat), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n796_), .B1(new_n795_), .B2(G106gat), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n794_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT53), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n801_), .B(new_n794_), .C1(new_n797_), .C2(new_n798_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n802_), .ZN(G1339gat));
  NAND3_X1  g602(.A1(new_n580_), .A2(new_n583_), .A3(new_n588_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n587_), .A2(new_n584_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n593_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n594_), .B1(new_n585_), .B2(new_n589_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n808_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n809_));
  AOI21_X1  g608(.A(KEYINPUT114), .B1(new_n549_), .B2(new_n673_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT114), .ZN(new_n811_));
  AOI211_X1 g610(.A(new_n811_), .B(new_n598_), .C1(new_n537_), .C2(new_n548_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n810_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT56), .ZN(new_n814_));
  OAI21_X1  g613(.A(KEYINPUT55), .B1(new_n545_), .B2(new_n546_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n516_), .A2(new_n517_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n527_), .A2(new_n816_), .A3(new_n817_), .A4(new_n544_), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n522_), .B(new_n544_), .C1(new_n539_), .C2(KEYINPUT12), .ZN(new_n819_));
  AOI22_X1  g618(.A1(new_n815_), .A2(new_n818_), .B1(new_n525_), .B2(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n814_), .B1(new_n820_), .B2(new_n536_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT115), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n536_), .A2(new_n814_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n822_), .B1(new_n820_), .B2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n819_), .A2(new_n525_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n817_), .B1(new_n518_), .B2(new_n527_), .ZN(new_n827_));
  NOR3_X1   g626(.A1(new_n545_), .A2(KEYINPUT55), .A3(new_n546_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n826_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n829_), .A2(KEYINPUT115), .A3(new_n823_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n821_), .A2(new_n825_), .A3(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n809_), .B1(new_n813_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT57), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n728_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n808_), .B1(new_n537_), .B2(new_n548_), .ZN(new_n836_));
  AOI21_X1  g635(.A(KEYINPUT56), .B1(new_n829_), .B2(new_n535_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n820_), .A2(new_n824_), .ZN(new_n838_));
  OAI211_X1 g637(.A(KEYINPUT58), .B(new_n836_), .C1(new_n837_), .C2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n662_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n637_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n657_), .ZN(new_n842_));
  AOI21_X1  g641(.A(KEYINPUT37), .B1(new_n842_), .B2(new_n651_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n839_), .B1(new_n840_), .B2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n838_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n821_), .ZN(new_n846_));
  AOI21_X1  g645(.A(KEYINPUT58), .B1(new_n846_), .B2(new_n836_), .ZN(new_n847_));
  OAI22_X1  g646(.A1(new_n832_), .A2(new_n835_), .B1(new_n844_), .B2(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n530_), .B1(new_n529_), .B2(new_n536_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n547_), .A2(KEYINPUT73), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n673_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n811_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n549_), .A2(KEYINPUT114), .A3(new_n673_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n831_), .A2(new_n852_), .A3(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n809_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(KEYINPUT57), .B1(new_n856_), .B2(new_n659_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n714_), .B1(new_n848_), .B2(new_n857_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n664_), .A2(new_n779_), .A3(new_n757_), .A4(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n757_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n859_), .B1(new_n862_), .B2(new_n663_), .ZN(new_n863_));
  AND2_X1   g662(.A1(new_n861_), .A2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n858_), .A2(new_n864_), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n683_), .A2(new_n411_), .A3(new_n442_), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n865_), .A2(new_n673_), .A3(new_n366_), .A4(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(G113gat), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(KEYINPUT116), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT116), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n867_), .A2(new_n871_), .A3(new_n868_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n847_), .ZN(new_n873_));
  OAI22_X1  g672(.A1(new_n849_), .A2(new_n850_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n874_), .B1(new_n845_), .B2(new_n821_), .ZN(new_n875_));
  AOI22_X1  g674(.A1(new_n875_), .A2(KEYINPUT58), .B1(new_n661_), .B2(new_n662_), .ZN(new_n876_));
  AOI22_X1  g675(.A1(new_n873_), .A2(new_n876_), .B1(new_n856_), .B2(new_n834_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n833_), .B1(new_n832_), .B2(new_n728_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n618_), .B1(new_n877_), .B2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n861_), .A2(new_n863_), .ZN(new_n880_));
  OAI211_X1 g679(.A(new_n366_), .B(new_n866_), .C1(new_n879_), .C2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT59), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n703_), .B1(new_n858_), .B2(new_n864_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n884_), .A2(KEYINPUT59), .A3(new_n866_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n885_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n602_), .A2(new_n868_), .ZN(new_n887_));
  AOI22_X1  g686(.A1(new_n870_), .A2(new_n872_), .B1(new_n886_), .B2(new_n887_), .ZN(G1340gat));
  INV_X1    g687(.A(new_n881_), .ZN(new_n889_));
  INV_X1    g688(.A(G120gat), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n890_), .B1(new_n779_), .B2(KEYINPUT60), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n889_), .B(new_n891_), .C1(KEYINPUT60), .C2(new_n890_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n779_), .B1(new_n883_), .B2(new_n885_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n893_), .B2(new_n890_), .ZN(G1341gat));
  AOI21_X1  g693(.A(G127gat), .B1(new_n889_), .B2(new_n618_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n618_), .A2(G127gat), .ZN(new_n896_));
  XOR2_X1   g695(.A(new_n896_), .B(KEYINPUT117), .Z(new_n897_));
  AOI21_X1  g696(.A(new_n895_), .B1(new_n886_), .B2(new_n897_), .ZN(G1342gat));
  AOI21_X1  g697(.A(G134gat), .B1(new_n889_), .B2(new_n728_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(KEYINPUT118), .B(G134gat), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n664_), .A2(new_n900_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n899_), .B1(new_n886_), .B2(new_n901_), .ZN(G1343gat));
  NOR4_X1   g701(.A1(new_n683_), .A2(new_n411_), .A3(new_n366_), .A4(new_n670_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n865_), .A2(new_n903_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n904_), .A2(new_n598_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(new_n316_), .ZN(G1344gat));
  NOR2_X1   g705(.A1(new_n904_), .A2(new_n779_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(KEYINPUT119), .B(G148gat), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n907_), .B(new_n908_), .ZN(G1345gat));
  OAI211_X1 g708(.A(new_n618_), .B(new_n903_), .C1(new_n879_), .C2(new_n880_), .ZN(new_n910_));
  XOR2_X1   g709(.A(KEYINPUT61), .B(G155gat), .Z(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(KEYINPUT120), .B(KEYINPUT121), .ZN(new_n913_));
  INV_X1    g712(.A(new_n911_), .ZN(new_n914_));
  NAND4_X1  g713(.A1(new_n865_), .A2(new_n618_), .A3(new_n903_), .A4(new_n914_), .ZN(new_n915_));
  AND3_X1   g714(.A1(new_n912_), .A2(new_n913_), .A3(new_n915_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n913_), .B1(new_n912_), .B2(new_n915_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n916_), .A2(new_n917_), .ZN(G1346gat));
  OAI21_X1  g717(.A(G162gat), .B1(new_n904_), .B2(new_n664_), .ZN(new_n919_));
  OR2_X1    g718(.A1(new_n659_), .A2(G162gat), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n919_), .B1(new_n904_), .B2(new_n920_), .ZN(G1347gat));
  NAND2_X1  g720(.A1(new_n683_), .A2(new_n413_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n922_), .ZN(new_n923_));
  NAND4_X1  g722(.A1(new_n865_), .A2(new_n673_), .A3(new_n366_), .A4(new_n923_), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT122), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n251_), .B1(new_n925_), .B2(KEYINPUT62), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n924_), .A2(new_n926_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT62), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n927_), .A2(KEYINPUT122), .A3(new_n928_), .ZN(new_n929_));
  NAND4_X1  g728(.A1(new_n884_), .A2(new_n673_), .A3(new_n275_), .A4(new_n923_), .ZN(new_n930_));
  OAI211_X1 g729(.A(new_n924_), .B(new_n926_), .C1(new_n925_), .C2(KEYINPUT62), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n929_), .A2(new_n930_), .A3(new_n931_), .ZN(G1348gat));
  NAND2_X1  g731(.A1(new_n865_), .A2(new_n366_), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT123), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n933_), .A2(new_n934_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n884_), .A2(KEYINPUT123), .ZN(new_n936_));
  NOR3_X1   g735(.A1(new_n779_), .A2(new_n255_), .A3(new_n922_), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n935_), .A2(new_n936_), .A3(new_n937_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n884_), .A2(new_n923_), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n255_), .B1(new_n939_), .B2(new_n779_), .ZN(new_n940_));
  AND2_X1   g739(.A1(new_n938_), .A2(new_n940_), .ZN(G1349gat));
  NOR3_X1   g740(.A1(new_n939_), .A2(new_n714_), .A3(new_n272_), .ZN(new_n942_));
  NAND4_X1  g741(.A1(new_n935_), .A2(new_n618_), .A3(new_n923_), .A4(new_n936_), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n942_), .B1(new_n943_), .B2(new_n227_), .ZN(G1350gat));
  OAI21_X1  g743(.A(G190gat), .B1(new_n939_), .B2(new_n664_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n728_), .A2(new_n233_), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n945_), .B1(new_n939_), .B2(new_n946_), .ZN(G1351gat));
  NAND3_X1  g746(.A1(new_n683_), .A2(new_n418_), .A3(new_n442_), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n948_), .B1(new_n858_), .B2(new_n864_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n949_), .A2(new_n673_), .ZN(new_n950_));
  XOR2_X1   g749(.A(KEYINPUT124), .B(G197gat), .Z(new_n951_));
  XNOR2_X1  g750(.A(new_n950_), .B(new_n951_), .ZN(G1352gat));
  NAND2_X1  g751(.A1(new_n949_), .A2(new_n555_), .ZN(new_n953_));
  AOI21_X1  g752(.A(new_n953_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n954_), .B1(new_n213_), .B2(new_n953_), .ZN(G1353gat));
  INV_X1    g754(.A(KEYINPUT125), .ZN(new_n956_));
  XNOR2_X1  g755(.A(KEYINPUT63), .B(G211gat), .ZN(new_n957_));
  NAND3_X1  g756(.A1(new_n949_), .A2(new_n618_), .A3(new_n957_), .ZN(new_n958_));
  INV_X1    g757(.A(new_n948_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n865_), .A2(new_n959_), .ZN(new_n960_));
  NOR2_X1   g759(.A1(new_n960_), .A2(new_n714_), .ZN(new_n961_));
  NOR2_X1   g760(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n962_));
  OAI211_X1 g761(.A(new_n956_), .B(new_n958_), .C1(new_n961_), .C2(new_n962_), .ZN(new_n963_));
  AND3_X1   g762(.A1(new_n949_), .A2(new_n618_), .A3(new_n957_), .ZN(new_n964_));
  AOI21_X1  g763(.A(new_n962_), .B1(new_n949_), .B2(new_n618_), .ZN(new_n965_));
  OAI21_X1  g764(.A(KEYINPUT125), .B1(new_n964_), .B2(new_n965_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n963_), .A2(new_n966_), .ZN(G1354gat));
  XNOR2_X1  g766(.A(KEYINPUT127), .B(G218gat), .ZN(new_n968_));
  NOR3_X1   g767(.A1(new_n960_), .A2(new_n664_), .A3(new_n968_), .ZN(new_n969_));
  OAI21_X1  g768(.A(KEYINPUT126), .B1(new_n960_), .B2(new_n659_), .ZN(new_n970_));
  INV_X1    g769(.A(KEYINPUT126), .ZN(new_n971_));
  NAND3_X1  g770(.A1(new_n949_), .A2(new_n971_), .A3(new_n728_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n970_), .A2(new_n972_), .ZN(new_n973_));
  AOI21_X1  g772(.A(new_n969_), .B1(new_n973_), .B2(new_n968_), .ZN(G1355gat));
endmodule


