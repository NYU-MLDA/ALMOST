//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 1 0 1 1 1 1 1 1 0 1 1 0 1 0 0 1 0 0 1 0 0 0 0 1 1 1 1 0 1 1 1 1 0 0 0 1 0 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n630_, new_n631_, new_n632_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n711_, new_n712_, new_n713_, new_n715_,
    new_n716_, new_n717_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n832_, new_n833_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n839_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n850_, new_n851_,
    new_n852_, new_n854_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n884_, new_n885_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_;
  NOR2_X1   g000(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G169gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G183gat), .ZN(new_n205_));
  INV_X1    g004(.A(G190gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT23), .B1(new_n205_), .B2(new_n206_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT23), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n209_), .A2(G183gat), .A3(G190gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n204_), .B1(new_n207_), .B2(new_n211_), .ZN(new_n212_));
  MUX2_X1   g011(.A(new_n210_), .B(new_n211_), .S(KEYINPUT79), .Z(new_n213_));
  OR3_X1    g012(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT95), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n215_), .B(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n218_), .B1(G169gat), .B2(G176gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT26), .B(G190gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(KEYINPUT94), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT25), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(G183gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n222_), .A2(G183gat), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n219_), .B1(new_n221_), .B2(new_n226_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n212_), .B1(new_n217_), .B2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G211gat), .B(G218gat), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n229_), .A2(KEYINPUT88), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(KEYINPUT88), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT89), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n230_), .A2(KEYINPUT89), .A3(new_n231_), .ZN(new_n235_));
  INV_X1    g034(.A(G197gat), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n236_), .A2(G204gat), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n236_), .A2(G204gat), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT87), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n237_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n240_), .B1(new_n239_), .B2(new_n238_), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n234_), .A2(new_n235_), .A3(KEYINPUT21), .A4(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT21), .B1(new_n238_), .B2(new_n237_), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n232_), .B(new_n243_), .C1(new_n241_), .C2(KEYINPUT21), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n228_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT20), .ZN(new_n248_));
  AND2_X1   g047(.A1(new_n213_), .A2(new_n207_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT26), .ZN(new_n250_));
  OAI21_X1  g049(.A(KEYINPUT78), .B1(new_n250_), .B2(G190gat), .ZN(new_n251_));
  OAI221_X1 g050(.A(new_n251_), .B1(new_n225_), .B2(KEYINPUT76), .C1(new_n224_), .C2(KEYINPUT77), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n220_), .A2(KEYINPUT78), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n225_), .A2(KEYINPUT76), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT77), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n254_), .B1(new_n223_), .B2(new_n255_), .ZN(new_n256_));
  NOR3_X1   g055(.A1(new_n252_), .A2(new_n253_), .A3(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n219_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n258_), .A2(new_n211_), .A3(new_n214_), .ZN(new_n259_));
  OAI22_X1  g058(.A1(new_n249_), .A2(new_n204_), .B1(new_n257_), .B2(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n248_), .B1(new_n260_), .B2(new_n245_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n247_), .A2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G226gat), .A2(G233gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n262_), .A2(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT20), .B1(new_n260_), .B2(new_n245_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT93), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT96), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n271_), .B1(new_n228_), .B2(new_n246_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n215_), .B(KEYINPUT95), .ZN(new_n273_));
  INV_X1    g072(.A(new_n227_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  OAI211_X1 g074(.A(KEYINPUT96), .B(new_n245_), .C1(new_n275_), .C2(new_n212_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n270_), .A2(new_n272_), .A3(new_n276_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n267_), .B1(new_n277_), .B2(new_n266_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G8gat), .B(G36gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT18), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G64gat), .B(G92gat), .ZN(new_n281_));
  XOR2_X1   g080(.A(new_n280_), .B(new_n281_), .Z(new_n282_));
  NAND3_X1  g081(.A1(new_n278_), .A2(KEYINPUT32), .A3(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n262_), .A2(new_n266_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n284_), .B1(new_n277_), .B2(new_n266_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n282_), .A2(KEYINPUT32), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G141gat), .A2(G148gat), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT81), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(G141gat), .A2(G148gat), .ZN(new_n291_));
  AND2_X1   g090(.A1(G155gat), .A2(G162gat), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n291_), .B1(new_n292_), .B2(KEYINPUT1), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G155gat), .B(G162gat), .ZN(new_n294_));
  OAI211_X1 g093(.A(new_n290_), .B(new_n293_), .C1(KEYINPUT1), .C2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT82), .ZN(new_n296_));
  OR2_X1    g095(.A1(new_n291_), .A2(KEYINPUT83), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n291_), .A2(KEYINPUT83), .ZN(new_n298_));
  NOR2_X1   g097(.A1(KEYINPUT84), .A2(KEYINPUT3), .ZN(new_n299_));
  AND2_X1   g098(.A1(KEYINPUT84), .A2(KEYINPUT3), .ZN(new_n300_));
  OAI211_X1 g099(.A(new_n297_), .B(new_n298_), .C1(new_n299_), .C2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT2), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n290_), .A2(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT85), .ZN(new_n305_));
  OR2_X1    g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n291_), .ZN(new_n307_));
  AOI22_X1  g106(.A1(new_n307_), .A2(KEYINPUT3), .B1(new_n304_), .B2(new_n305_), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n301_), .A2(new_n303_), .A3(new_n306_), .A4(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n294_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n296_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G127gat), .B(G134gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT80), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G113gat), .B(G120gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n313_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n317_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n312_), .A2(new_n319_), .ZN(new_n320_));
  AND2_X1   g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT97), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G225gat), .A2(G233gat), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n321_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT4), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n312_), .A2(new_n325_), .A3(new_n319_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n323_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n318_), .A2(new_n320_), .ZN(new_n328_));
  OAI211_X1 g127(.A(new_n326_), .B(new_n327_), .C1(new_n328_), .C2(new_n325_), .ZN(new_n329_));
  OAI21_X1  g128(.A(KEYINPUT97), .B1(new_n328_), .B2(new_n327_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n324_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G1gat), .B(G29gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(G85gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT0), .B(G57gat), .ZN(new_n334_));
  XOR2_X1   g133(.A(new_n333_), .B(new_n334_), .Z(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n331_), .A2(new_n336_), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n324_), .A2(new_n329_), .A3(new_n335_), .A4(new_n330_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n283_), .A2(new_n287_), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n282_), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n272_), .A2(new_n276_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n265_), .B1(new_n342_), .B2(new_n270_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n341_), .B1(new_n343_), .B2(new_n284_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT33), .ZN(new_n345_));
  OR2_X1    g144(.A1(new_n338_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n277_), .A2(new_n266_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n284_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n347_), .A2(new_n282_), .A3(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n335_), .B1(new_n321_), .B2(new_n327_), .ZN(new_n350_));
  OAI211_X1 g149(.A(new_n326_), .B(new_n323_), .C1(new_n328_), .C2(new_n325_), .ZN(new_n351_));
  AND3_X1   g150(.A1(new_n350_), .A2(KEYINPUT99), .A3(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(KEYINPUT99), .B1(new_n350_), .B2(new_n351_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n344_), .A2(new_n346_), .A3(new_n349_), .A4(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT98), .ZN(new_n356_));
  AND3_X1   g155(.A1(new_n338_), .A2(new_n356_), .A3(new_n345_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n356_), .B1(new_n338_), .B2(new_n345_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n340_), .B1(new_n355_), .B2(new_n359_), .ZN(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT28), .B1(new_n312_), .B2(KEYINPUT29), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NOR3_X1   g161(.A1(new_n312_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G22gat), .B(G50gat), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NOR3_X1   g164(.A1(new_n362_), .A2(new_n363_), .A3(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n363_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n364_), .B1(new_n367_), .B2(new_n361_), .ZN(new_n368_));
  OAI21_X1  g167(.A(KEYINPUT86), .B1(new_n366_), .B2(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n365_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n367_), .A2(new_n361_), .A3(new_n364_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT86), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n370_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT29), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n245_), .B1(new_n313_), .B2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G228gat), .A2(G233gat), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n376_), .B1(new_n245_), .B2(KEYINPUT90), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  OAI221_X1 g177(.A(new_n245_), .B1(KEYINPUT90), .B2(new_n376_), .C1(new_n313_), .C2(new_n374_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G78gat), .B(G106gat), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n381_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n383_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n369_), .B(new_n373_), .C1(new_n382_), .C2(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(KEYINPUT91), .B1(new_n380_), .B2(new_n381_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n384_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT91), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n378_), .A2(new_n379_), .A3(new_n388_), .A4(new_n383_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n366_), .A2(new_n368_), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n386_), .A2(new_n387_), .A3(new_n389_), .A4(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n385_), .A2(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G71gat), .B(G99gat), .ZN(new_n393_));
  INV_X1    g192(.A(G43gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n260_), .B(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(new_n319_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G227gat), .A2(G233gat), .ZN(new_n398_));
  INV_X1    g197(.A(G15gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT30), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT31), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n397_), .A2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n396_), .B(new_n317_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n402_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n403_), .A2(new_n406_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n392_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n407_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n392_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n407_), .A2(new_n385_), .A3(new_n391_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n339_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n344_), .A2(new_n349_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT27), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n414_), .B1(new_n285_), .B2(new_n282_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n278_), .A2(new_n341_), .ZN(new_n416_));
  AOI22_X1  g215(.A1(new_n413_), .A2(new_n414_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  AOI22_X1  g216(.A1(new_n360_), .A2(new_n408_), .B1(new_n412_), .B2(new_n417_), .ZN(new_n418_));
  XOR2_X1   g217(.A(G29gat), .B(G36gat), .Z(new_n419_));
  XOR2_X1   g218(.A(G43gat), .B(G50gat), .Z(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(KEYINPUT15), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G15gat), .B(G22gat), .ZN(new_n423_));
  INV_X1    g222(.A(G1gat), .ZN(new_n424_));
  INV_X1    g223(.A(G8gat), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT14), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n423_), .A2(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G1gat), .B(G8gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n427_), .B(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n422_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n429_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(new_n421_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G229gat), .A2(G233gat), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n430_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n421_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n429_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n432_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n433_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n439_), .A2(KEYINPUT75), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n439_), .A2(KEYINPUT75), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n434_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G113gat), .B(G141gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G169gat), .B(G197gat), .ZN(new_n444_));
  XOR2_X1   g243(.A(new_n443_), .B(new_n444_), .Z(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n442_), .A2(new_n446_), .ZN(new_n447_));
  OAI211_X1 g246(.A(new_n434_), .B(new_n445_), .C1(new_n440_), .C2(new_n441_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n418_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(G99gat), .A2(G106gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT6), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT6), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n454_), .A2(G99gat), .A3(G106gat), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT67), .ZN(new_n456_));
  AND3_X1   g255(.A1(new_n453_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n456_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT7), .ZN(new_n459_));
  INV_X1    g258(.A(G99gat), .ZN(new_n460_));
  INV_X1    g259(.A(G106gat), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n459_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NOR3_X1   g263(.A1(new_n457_), .A2(new_n458_), .A3(new_n464_), .ZN(new_n465_));
  XOR2_X1   g264(.A(G85gat), .B(G92gat), .Z(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  OAI21_X1  g266(.A(KEYINPUT8), .B1(new_n465_), .B2(new_n467_), .ZN(new_n468_));
  AND2_X1   g267(.A1(new_n462_), .A2(new_n463_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n453_), .A2(new_n455_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  OR2_X1    g270(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n472_));
  NAND2_X1  g271(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n471_), .A2(new_n466_), .A3(new_n472_), .A4(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT65), .ZN(new_n475_));
  OAI211_X1 g274(.A(G85gat), .B(G92gat), .C1(KEYINPUT64), .C2(KEYINPUT9), .ZN(new_n476_));
  OAI211_X1 g275(.A(KEYINPUT64), .B(KEYINPUT9), .C1(G85gat), .C2(G92gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND4_X1  g277(.A1(KEYINPUT64), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  OR2_X1    g280(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n482_), .A2(new_n461_), .A3(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(new_n470_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n475_), .B1(new_n481_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n485_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n487_), .A2(KEYINPUT65), .A3(new_n480_), .ZN(new_n488_));
  AOI22_X1  g287(.A1(new_n468_), .A2(new_n474_), .B1(new_n486_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(G71gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(KEYINPUT68), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT68), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(G71gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n491_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(G78gat), .ZN(new_n495_));
  INV_X1    g294(.A(G78gat), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n491_), .A2(new_n493_), .A3(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(G64gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(G57gat), .ZN(new_n499_));
  INV_X1    g298(.A(G57gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(G64gat), .ZN(new_n501_));
  AND3_X1   g300(.A1(new_n499_), .A2(new_n501_), .A3(KEYINPUT11), .ZN(new_n502_));
  AOI21_X1  g301(.A(KEYINPUT11), .B1(new_n499_), .B2(new_n501_), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n495_), .B(new_n497_), .C1(new_n502_), .C2(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n499_), .A2(new_n501_), .A3(KEYINPUT11), .ZN(new_n505_));
  INV_X1    g304(.A(new_n497_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n496_), .B1(new_n491_), .B2(new_n493_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n505_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  AND2_X1   g307(.A1(new_n504_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n489_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT8), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n470_), .A2(KEYINPUT67), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n453_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n512_), .A2(new_n513_), .A3(new_n469_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n511_), .B1(new_n514_), .B2(new_n466_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n466_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n516_), .B1(new_n470_), .B2(new_n469_), .ZN(new_n517_));
  AOI21_X1  g316(.A(KEYINPUT65), .B1(new_n487_), .B2(new_n480_), .ZN(new_n518_));
  AND4_X1   g317(.A1(KEYINPUT65), .A2(new_n480_), .A3(new_n470_), .A4(new_n484_), .ZN(new_n519_));
  OAI22_X1  g318(.A1(new_n515_), .A2(new_n517_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n509_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n510_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(G230gat), .ZN(new_n524_));
  INV_X1    g323(.A(G233gat), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n523_), .A2(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n526_), .B1(new_n489_), .B2(new_n509_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n458_), .A2(new_n464_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n467_), .B1(new_n529_), .B2(new_n513_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n474_), .B1(new_n530_), .B2(new_n511_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n486_), .A2(new_n488_), .ZN(new_n532_));
  AOI211_X1 g331(.A(KEYINPUT12), .B(new_n509_), .C1(new_n531_), .C2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT12), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n534_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n528_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G120gat), .B(G148gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT5), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G176gat), .B(G204gat), .ZN(new_n539_));
  XOR2_X1   g338(.A(new_n538_), .B(new_n539_), .Z(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n527_), .A2(new_n536_), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n541_), .B1(new_n527_), .B2(new_n536_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n545_), .A2(KEYINPUT13), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n545_), .A2(KEYINPUT13), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT69), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n549_), .A2(new_n550_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT74), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G127gat), .B(G155gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT16), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G183gat), .B(G211gat), .ZN(new_n558_));
  XOR2_X1   g357(.A(new_n557_), .B(new_n558_), .Z(new_n559_));
  NAND2_X1  g358(.A1(G231gat), .A2(G233gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n429_), .B(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(new_n521_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(KEYINPUT73), .B(KEYINPUT17), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n559_), .B1(new_n562_), .B2(new_n564_), .ZN(new_n565_));
  XOR2_X1   g364(.A(KEYINPUT72), .B(KEYINPUT17), .Z(new_n566_));
  NAND2_X1  g365(.A1(new_n562_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  NOR3_X1   g367(.A1(new_n562_), .A2(new_n559_), .A3(new_n564_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n555_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n569_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n571_), .A2(KEYINPUT74), .A3(new_n565_), .A4(new_n567_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT37), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n422_), .A2(new_n520_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G232gat), .A2(G233gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT71), .ZN(new_n577_));
  XOR2_X1   g376(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n579_), .A2(KEYINPUT35), .ZN(new_n580_));
  OAI211_X1 g379(.A(new_n575_), .B(new_n580_), .C1(new_n435_), .C2(new_n520_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(KEYINPUT35), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  OR2_X1    g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n581_), .A2(new_n583_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G190gat), .B(G218gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G134gat), .B(G162gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n588_), .A2(KEYINPUT36), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n584_), .A2(new_n585_), .A3(new_n589_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n584_), .A2(new_n585_), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n588_), .B(KEYINPUT36), .Z(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n574_), .B(new_n590_), .C1(new_n591_), .C2(new_n593_), .ZN(new_n594_));
  AND3_X1   g393(.A1(new_n584_), .A2(new_n585_), .A3(new_n589_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n593_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n596_));
  OAI21_X1  g395(.A(KEYINPUT37), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  AND2_X1   g396(.A1(new_n594_), .A2(new_n597_), .ZN(new_n598_));
  NOR3_X1   g397(.A1(new_n554_), .A2(new_n573_), .A3(new_n598_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n451_), .A2(new_n599_), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n339_), .B(KEYINPUT100), .Z(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n600_), .A2(new_n424_), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT38), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT101), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n590_), .B1(new_n591_), .B2(new_n593_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n418_), .A2(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n552_), .A2(new_n449_), .A3(new_n553_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n610_), .A2(new_n573_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n609_), .A2(new_n611_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n612_), .A2(new_n339_), .ZN(new_n613_));
  OAI221_X1 g412(.A(new_n606_), .B1(new_n604_), .B2(new_n603_), .C1(new_n424_), .C2(new_n613_), .ZN(G1324gat));
  INV_X1    g413(.A(new_n417_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n600_), .A2(new_n425_), .A3(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT102), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n609_), .A2(new_n617_), .A3(new_n615_), .A4(new_n611_), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n618_), .A2(G8gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(KEYINPUT103), .B(KEYINPUT39), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n609_), .A2(new_n615_), .A3(new_n611_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(KEYINPUT102), .ZN(new_n622_));
  AND3_X1   g421(.A1(new_n619_), .A2(new_n620_), .A3(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n620_), .B1(new_n619_), .B2(new_n622_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n616_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT40), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  OAI211_X1 g426(.A(KEYINPUT40), .B(new_n616_), .C1(new_n623_), .C2(new_n624_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(G1325gat));
  AOI21_X1  g428(.A(new_n399_), .B1(new_n612_), .B2(new_n407_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT41), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n600_), .A2(new_n399_), .A3(new_n407_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(G1326gat));
  INV_X1    g432(.A(G22gat), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n634_), .B1(new_n612_), .B2(new_n392_), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n635_), .B(KEYINPUT42), .Z(new_n636_));
  NAND2_X1  g435(.A1(new_n392_), .A2(new_n634_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT104), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n600_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n636_), .A2(new_n639_), .ZN(G1327gat));
  NAND2_X1  g439(.A1(new_n360_), .A2(new_n408_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n412_), .A2(new_n417_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n554_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n573_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n645_), .A2(new_n607_), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n643_), .A2(new_n449_), .A3(new_n644_), .A4(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n339_), .ZN(new_n648_));
  OR3_X1    g447(.A1(new_n647_), .A2(G29gat), .A3(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT106), .ZN(new_n650_));
  INV_X1    g449(.A(new_n610_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(KEYINPUT105), .A2(KEYINPUT43), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(KEYINPUT105), .A2(KEYINPUT43), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n655_), .B1(new_n643_), .B2(new_n598_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n594_), .A2(new_n597_), .ZN(new_n657_));
  AOI211_X1 g456(.A(new_n657_), .B(new_n653_), .C1(new_n641_), .C2(new_n642_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n651_), .B1(new_n656_), .B2(new_n658_), .ZN(new_n659_));
  OAI211_X1 g458(.A(new_n650_), .B(KEYINPUT44), .C1(new_n659_), .C2(new_n645_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT44), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n645_), .A2(new_n650_), .ZN(new_n662_));
  OAI22_X1  g461(.A1(new_n418_), .A2(new_n657_), .B1(new_n653_), .B2(new_n654_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n643_), .A2(new_n598_), .A3(new_n652_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n610_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  OAI211_X1 g464(.A(new_n661_), .B(new_n662_), .C1(new_n665_), .C2(KEYINPUT106), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n660_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT107), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n667_), .A2(new_n668_), .A3(new_n602_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(G29gat), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n668_), .B1(new_n667_), .B2(new_n602_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n649_), .B1(new_n670_), .B2(new_n671_), .ZN(G1328gat));
  NOR3_X1   g471(.A1(new_n647_), .A2(G36gat), .A3(new_n417_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT45), .Z(new_n674_));
  AOI21_X1  g473(.A(new_n417_), .B1(new_n660_), .B2(new_n666_), .ZN(new_n675_));
  INV_X1    g474(.A(G36gat), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n674_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT46), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n674_), .B(KEYINPUT46), .C1(new_n675_), .C2(new_n676_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(G1329gat));
  XNOR2_X1  g480(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n394_), .B1(new_n667_), .B2(new_n407_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n407_), .A2(new_n394_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n647_), .A2(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n683_), .B1(new_n684_), .B2(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n409_), .B1(new_n660_), .B2(new_n666_), .ZN(new_n688_));
  OAI221_X1 g487(.A(new_n682_), .B1(new_n647_), .B2(new_n685_), .C1(new_n688_), .C2(new_n394_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n689_), .ZN(G1330gat));
  INV_X1    g489(.A(new_n392_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n647_), .A2(new_n691_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n692_), .A2(G50gat), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n392_), .A2(G50gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n667_), .B2(new_n694_), .ZN(G1331gat));
  NAND3_X1  g494(.A1(new_n554_), .A2(new_n645_), .A3(new_n657_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT109), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n418_), .A2(new_n449_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n696_), .A2(new_n697_), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n698_), .A2(new_n699_), .A3(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(new_n602_), .ZN(new_n702_));
  AND3_X1   g501(.A1(new_n702_), .A2(KEYINPUT110), .A3(new_n500_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n573_), .A2(new_n449_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n609_), .A2(new_n554_), .A3(new_n704_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(KEYINPUT111), .B(G57gat), .ZN(new_n706_));
  NOR3_X1   g505(.A1(new_n705_), .A2(new_n648_), .A3(new_n706_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT112), .ZN(new_n708_));
  AOI21_X1  g507(.A(KEYINPUT110), .B1(new_n702_), .B2(new_n500_), .ZN(new_n709_));
  NOR3_X1   g508(.A1(new_n703_), .A2(new_n708_), .A3(new_n709_), .ZN(G1332gat));
  OAI21_X1  g509(.A(G64gat), .B1(new_n705_), .B2(new_n417_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT48), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n701_), .A2(new_n498_), .A3(new_n615_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1333gat));
  OAI21_X1  g513(.A(G71gat), .B1(new_n705_), .B2(new_n409_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT49), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n701_), .A2(new_n490_), .A3(new_n407_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(G1334gat));
  OAI21_X1  g517(.A(G78gat), .B1(new_n705_), .B2(new_n691_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT50), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n701_), .A2(new_n496_), .A3(new_n392_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1335gat));
  NAND3_X1  g521(.A1(new_n554_), .A2(new_n450_), .A3(new_n573_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n723_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n724_), .A2(new_n339_), .ZN(new_n725_));
  INV_X1    g524(.A(G85gat), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n699_), .A2(new_n554_), .A3(new_n646_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n602_), .A2(new_n726_), .ZN(new_n728_));
  OAI22_X1  g527(.A1(new_n725_), .A2(new_n726_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT113), .ZN(G1336gat));
  AND2_X1   g529(.A1(new_n724_), .A2(new_n615_), .ZN(new_n731_));
  INV_X1    g530(.A(G92gat), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n615_), .A2(new_n732_), .ZN(new_n733_));
  OAI22_X1  g532(.A1(new_n731_), .A2(new_n732_), .B1(new_n727_), .B2(new_n733_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT114), .Z(G1337gat));
  NAND2_X1  g534(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n407_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n736_), .B1(new_n727_), .B2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n724_), .A2(new_n407_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n739_), .B2(G99gat), .ZN(new_n740_));
  NOR2_X1   g539(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n740_), .B(new_n741_), .ZN(G1338gat));
  NOR3_X1   g541(.A1(new_n727_), .A2(G106gat), .A3(new_n691_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT116), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n461_), .B1(new_n724_), .B2(new_n392_), .ZN(new_n745_));
  OR2_X1    g544(.A1(new_n745_), .A2(KEYINPUT52), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(KEYINPUT52), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n744_), .A2(new_n746_), .A3(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(KEYINPUT53), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT53), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n744_), .A2(new_n746_), .A3(new_n750_), .A4(new_n747_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n749_), .A2(new_n751_), .ZN(G1339gat));
  XNOR2_X1  g551(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n704_), .A2(new_n548_), .A3(new_n547_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n754_), .B1(new_n755_), .B2(new_n598_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n549_), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n757_), .A2(new_n657_), .A3(new_n704_), .A4(new_n753_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n445_), .B1(new_n437_), .B2(new_n433_), .ZN(new_n760_));
  OR2_X1    g559(.A1(new_n760_), .A2(KEYINPUT119), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n437_), .A2(new_n433_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n762_), .A2(KEYINPUT119), .A3(new_n446_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n430_), .A2(new_n432_), .A3(new_n438_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n761_), .A2(new_n763_), .A3(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n448_), .A2(new_n765_), .A3(new_n542_), .ZN(new_n766_));
  OAI211_X1 g565(.A(new_n528_), .B(KEYINPUT55), .C1(new_n533_), .C2(new_n535_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT118), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(KEYINPUT12), .B1(new_n489_), .B2(new_n509_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n520_), .A2(new_n534_), .A3(new_n521_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n772_), .A2(KEYINPUT118), .A3(KEYINPUT55), .A4(new_n528_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT55), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n536_), .A2(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n510_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n526_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n769_), .A2(new_n773_), .A3(new_n775_), .A4(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(new_n540_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT56), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n778_), .A2(KEYINPUT56), .A3(new_n540_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n766_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n657_), .B1(new_n783_), .B2(KEYINPUT58), .ZN(new_n784_));
  XOR2_X1   g583(.A(KEYINPUT121), .B(KEYINPUT58), .Z(new_n785_));
  OAI21_X1  g584(.A(new_n785_), .B1(new_n783_), .B2(KEYINPUT120), .ZN(new_n786_));
  INV_X1    g585(.A(new_n766_), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n778_), .A2(KEYINPUT56), .A3(new_n540_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT56), .B1(new_n778_), .B2(new_n540_), .ZN(new_n789_));
  OAI211_X1 g588(.A(KEYINPUT120), .B(new_n787_), .C1(new_n788_), .C2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n784_), .B1(new_n786_), .B2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n449_), .A2(new_n542_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n793_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n765_), .A2(new_n448_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n545_), .A2(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n607_), .B1(new_n794_), .B2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT57), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n788_), .A2(new_n789_), .ZN(new_n800_));
  OAI22_X1  g599(.A1(new_n800_), .A2(new_n793_), .B1(new_n545_), .B2(new_n795_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n801_), .A2(KEYINPUT57), .A3(new_n607_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n792_), .A2(new_n799_), .A3(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n759_), .B1(new_n803_), .B2(new_n573_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n615_), .A2(new_n601_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n411_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(KEYINPUT59), .B1(new_n804_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT122), .ZN(new_n809_));
  OAI211_X1 g608(.A(KEYINPUT58), .B(new_n787_), .C1(new_n788_), .C2(new_n789_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n598_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n785_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n787_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT120), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n812_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n811_), .B1(new_n815_), .B2(new_n790_), .ZN(new_n816_));
  AOI21_X1  g615(.A(KEYINPUT57), .B1(new_n801_), .B2(new_n607_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n809_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n792_), .A2(KEYINPUT122), .A3(new_n799_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n818_), .A2(new_n819_), .A3(new_n802_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n759_), .B1(new_n820_), .B2(new_n573_), .ZN(new_n821_));
  OR2_X1    g620(.A1(new_n807_), .A2(KEYINPUT59), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n808_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT123), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n808_), .B(KEYINPUT123), .C1(new_n821_), .C2(new_n822_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n825_), .A2(new_n449_), .A3(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(G113gat), .ZN(new_n828_));
  OR2_X1    g627(.A1(new_n804_), .A2(new_n807_), .ZN(new_n829_));
  OR2_X1    g628(.A1(new_n450_), .A2(G113gat), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n828_), .B1(new_n829_), .B2(new_n830_), .ZN(G1340gat));
  OAI21_X1  g630(.A(G120gat), .B1(new_n823_), .B2(new_n644_), .ZN(new_n832_));
  INV_X1    g631(.A(G120gat), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n833_), .B1(new_n644_), .B2(KEYINPUT60), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n834_), .B1(KEYINPUT60), .B2(new_n833_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n832_), .B1(new_n829_), .B2(new_n835_), .ZN(G1341gat));
  NAND3_X1  g635(.A1(new_n825_), .A2(new_n645_), .A3(new_n826_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(G127gat), .ZN(new_n838_));
  OR2_X1    g637(.A1(new_n573_), .A2(G127gat), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n838_), .B1(new_n829_), .B2(new_n839_), .ZN(G1342gat));
  INV_X1    g639(.A(G134gat), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n657_), .A2(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n825_), .A2(new_n826_), .A3(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n841_), .B1(new_n829_), .B2(new_n607_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT124), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n843_), .A2(KEYINPUT124), .A3(new_n844_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(G1343gat));
  NOR2_X1   g648(.A1(new_n804_), .A2(new_n410_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n805_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n851_), .A2(new_n450_), .ZN(new_n852_));
  XOR2_X1   g651(.A(new_n852_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g652(.A1(new_n851_), .A2(new_n644_), .ZN(new_n854_));
  XOR2_X1   g653(.A(new_n854_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g654(.A1(new_n851_), .A2(new_n573_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(KEYINPUT61), .B(G155gat), .ZN(new_n857_));
  XOR2_X1   g656(.A(new_n856_), .B(new_n857_), .Z(G1346gat));
  OAI21_X1  g657(.A(G162gat), .B1(new_n851_), .B2(new_n657_), .ZN(new_n859_));
  OR2_X1    g658(.A1(new_n607_), .A2(G162gat), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n851_), .B2(new_n860_), .ZN(G1347gat));
  NOR2_X1   g660(.A1(new_n602_), .A2(new_n417_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n806_), .ZN(new_n863_));
  NOR3_X1   g662(.A1(new_n821_), .A2(new_n450_), .A3(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(G169gat), .ZN(new_n865_));
  OAI21_X1  g664(.A(KEYINPUT125), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  OR2_X1    g665(.A1(new_n866_), .A2(KEYINPUT62), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n865_), .A2(KEYINPUT22), .ZN(new_n868_));
  OR2_X1    g667(.A1(new_n865_), .A2(KEYINPUT22), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n864_), .A2(new_n868_), .A3(new_n869_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n864_), .A2(KEYINPUT125), .A3(new_n865_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n866_), .A2(KEYINPUT62), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n867_), .B(new_n870_), .C1(new_n871_), .C2(new_n872_), .ZN(G1348gat));
  NOR2_X1   g672(.A1(new_n821_), .A2(new_n863_), .ZN(new_n874_));
  AOI21_X1  g673(.A(G176gat), .B1(new_n874_), .B2(new_n554_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n804_), .A2(new_n392_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n862_), .A2(new_n407_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  AND3_X1   g677(.A1(new_n878_), .A2(G176gat), .A3(new_n554_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n875_), .B1(new_n876_), .B2(new_n879_), .ZN(G1349gat));
  NOR2_X1   g679(.A1(new_n573_), .A2(new_n226_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n876_), .A2(new_n645_), .A3(new_n878_), .ZN(new_n882_));
  AOI22_X1  g681(.A1(new_n874_), .A2(new_n881_), .B1(new_n882_), .B2(new_n205_), .ZN(G1350gat));
  NAND3_X1  g682(.A1(new_n874_), .A2(new_n221_), .A3(new_n608_), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n821_), .A2(new_n657_), .A3(new_n863_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n885_), .B2(new_n206_), .ZN(G1351gat));
  NAND3_X1  g685(.A1(new_n850_), .A2(new_n615_), .A3(new_n648_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n887_), .A2(new_n450_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(new_n236_), .ZN(G1352gat));
  NOR2_X1   g688(.A1(new_n887_), .A2(new_n644_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  XOR2_X1   g691(.A(KEYINPUT126), .B(G204gat), .Z(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n890_), .B2(new_n893_), .ZN(G1353gat));
  NOR2_X1   g693(.A1(new_n887_), .A2(new_n573_), .ZN(new_n895_));
  NOR3_X1   g694(.A1(new_n895_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n896_));
  XOR2_X1   g695(.A(KEYINPUT63), .B(G211gat), .Z(new_n897_));
  AOI21_X1  g696(.A(new_n896_), .B1(new_n895_), .B2(new_n897_), .ZN(G1354gat));
  INV_X1    g697(.A(G218gat), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n887_), .A2(new_n899_), .A3(new_n657_), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n887_), .A2(KEYINPUT127), .A3(new_n607_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n901_), .A2(G218gat), .ZN(new_n902_));
  OAI21_X1  g701(.A(KEYINPUT127), .B1(new_n887_), .B2(new_n607_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n900_), .B1(new_n902_), .B2(new_n903_), .ZN(G1355gat));
endmodule


