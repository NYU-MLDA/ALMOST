//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 0 0 0 1 1 0 1 0 0 0 1 1 1 0 1 0 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 0 1 1 0 1 1 0 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n713_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n774_, new_n775_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n817_, new_n818_, new_n819_, new_n821_,
    new_n822_, new_n823_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n922_, new_n923_,
    new_n925_, new_n927_, new_n928_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n949_, new_n950_, new_n951_, new_n953_,
    new_n954_, new_n956_, new_n957_, new_n958_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n966_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n975_, new_n976_,
    new_n977_, new_n978_, new_n979_, new_n980_, new_n981_;
  XNOR2_X1  g000(.A(G71gat), .B(G78gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G57gat), .B(G64gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT67), .ZN(new_n204_));
  AOI21_X1  g003(.A(new_n202_), .B1(new_n204_), .B2(KEYINPUT11), .ZN(new_n205_));
  AND2_X1   g004(.A1(new_n203_), .A2(KEYINPUT67), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n203_), .A2(KEYINPUT67), .ZN(new_n207_));
  OR3_X1    g006(.A1(new_n206_), .A2(new_n207_), .A3(KEYINPUT11), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n205_), .A2(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n204_), .A2(KEYINPUT11), .A3(new_n202_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT12), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT8), .ZN(new_n214_));
  OR2_X1    g013(.A1(KEYINPUT66), .A2(KEYINPUT6), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G99gat), .A2(G106gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(KEYINPUT66), .A2(KEYINPUT6), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  AND2_X1   g017(.A1(G99gat), .A2(G106gat), .ZN(new_n219_));
  AND2_X1   g018(.A1(KEYINPUT66), .A2(KEYINPUT6), .ZN(new_n220_));
  NOR2_X1   g019(.A1(KEYINPUT66), .A2(KEYINPUT6), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n219_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n223_));
  AND3_X1   g022(.A1(new_n218_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G99gat), .ZN(new_n225_));
  INV_X1    g024(.A(G106gat), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT7), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n225_), .B(new_n226_), .C1(new_n227_), .C2(KEYINPUT64), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT64), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n229_), .A2(KEYINPUT7), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT65), .B1(new_n228_), .B2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n227_), .A2(KEYINPUT64), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n229_), .A2(KEYINPUT7), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT65), .ZN(new_n234_));
  NOR2_X1   g033(.A1(G99gat), .A2(G106gat), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n232_), .A2(new_n233_), .A3(new_n234_), .A4(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n231_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n224_), .A2(new_n237_), .ZN(new_n238_));
  XOR2_X1   g037(.A(G85gat), .B(G92gat), .Z(new_n239_));
  AOI21_X1  g038(.A(new_n214_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n239_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n219_), .A2(KEYINPUT6), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT6), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n216_), .A2(new_n243_), .ZN(new_n244_));
  AND3_X1   g043(.A1(new_n242_), .A2(new_n244_), .A3(new_n223_), .ZN(new_n245_));
  AOI211_X1 g044(.A(KEYINPUT8), .B(new_n241_), .C1(new_n237_), .C2(new_n245_), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT70), .B1(new_n240_), .B2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n237_), .A2(new_n245_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n241_), .A2(KEYINPUT8), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT70), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n241_), .B1(new_n224_), .B2(new_n237_), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n250_), .B(new_n251_), .C1(new_n252_), .C2(new_n214_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n247_), .A2(new_n253_), .ZN(new_n254_));
  XOR2_X1   g053(.A(KEYINPUT10), .B(G99gat), .Z(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(new_n226_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n239_), .A2(KEYINPUT9), .ZN(new_n257_));
  AND2_X1   g056(.A1(new_n242_), .A2(new_n244_), .ZN(new_n258_));
  INV_X1    g057(.A(G85gat), .ZN(new_n259_));
  INV_X1    g058(.A(G92gat), .ZN(new_n260_));
  OR3_X1    g059(.A1(new_n259_), .A2(new_n260_), .A3(KEYINPUT9), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n256_), .A2(new_n257_), .A3(new_n258_), .A4(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(KEYINPUT71), .B1(new_n254_), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT71), .ZN(new_n264_));
  INV_X1    g063(.A(new_n262_), .ZN(new_n265_));
  AOI211_X1 g064(.A(new_n264_), .B(new_n265_), .C1(new_n247_), .C2(new_n253_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n213_), .B1(new_n263_), .B2(new_n266_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n240_), .A2(new_n246_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n268_), .A2(new_n265_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n212_), .B1(new_n269_), .B2(new_n211_), .ZN(new_n270_));
  AND2_X1   g069(.A1(G230gat), .A2(G233gat), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n271_), .B1(new_n269_), .B2(new_n211_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n267_), .A2(new_n270_), .A3(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT69), .B1(new_n269_), .B2(new_n211_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT68), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n269_), .A2(new_n275_), .A3(new_n211_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n211_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n262_), .B1(new_n240_), .B2(new_n246_), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT68), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT69), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n277_), .A2(new_n280_), .A3(new_n278_), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n274_), .A2(new_n276_), .A3(new_n279_), .A4(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(new_n271_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n273_), .A2(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(G120gat), .B(G148gat), .Z(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G176gat), .B(G204gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n284_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT73), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n273_), .A2(new_n283_), .A3(new_n289_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n291_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n284_), .A2(KEYINPUT73), .A3(new_n290_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT13), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n294_), .A2(KEYINPUT13), .A3(new_n295_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  XOR2_X1   g099(.A(G134gat), .B(G162gat), .Z(new_n301_));
  XNOR2_X1  g100(.A(G190gat), .B(G218gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT36), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  OR2_X1    g104(.A1(new_n303_), .A2(new_n304_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G29gat), .B(G36gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT75), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G43gat), .B(G50gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT15), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n311_), .B1(new_n263_), .B2(new_n266_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT76), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n269_), .A2(new_n310_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n312_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G232gat), .A2(G233gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT35), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  AND3_X1   g121(.A1(new_n314_), .A2(new_n316_), .A3(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n322_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n324_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n320_), .A2(new_n321_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n312_), .A2(new_n315_), .A3(new_n326_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n325_), .A2(new_n327_), .ZN(new_n328_));
  OAI211_X1 g127(.A(new_n305_), .B(new_n306_), .C1(new_n323_), .C2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n314_), .A2(new_n322_), .ZN(new_n330_));
  AND3_X1   g129(.A1(new_n312_), .A2(new_n315_), .A3(new_n326_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n325_), .A2(new_n316_), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n332_), .A2(new_n304_), .A3(new_n303_), .A4(new_n333_), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n329_), .A2(new_n334_), .A3(KEYINPUT77), .A4(KEYINPUT37), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n329_), .A2(new_n334_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT77), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT37), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(KEYINPUT77), .A2(KEYINPUT37), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n336_), .A2(new_n340_), .A3(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT81), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G231gat), .A2(G233gat), .ZN(new_n345_));
  XOR2_X1   g144(.A(new_n211_), .B(new_n345_), .Z(new_n346_));
  XOR2_X1   g145(.A(G15gat), .B(G22gat), .Z(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT78), .B(G1gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(G8gat), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n347_), .B1(new_n349_), .B2(KEYINPUT14), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT79), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G1gat), .B(G8gat), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n351_), .B(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n346_), .B(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G127gat), .B(G155gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(KEYINPUT16), .ZN(new_n357_));
  XOR2_X1   g156(.A(G183gat), .B(G211gat), .Z(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT17), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n355_), .A2(new_n361_), .ZN(new_n362_));
  OR2_X1    g161(.A1(new_n346_), .A2(new_n354_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n346_), .A2(new_n354_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT17), .ZN(new_n365_));
  OAI211_X1 g164(.A(new_n363_), .B(new_n364_), .C1(new_n365_), .C2(new_n359_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT80), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n362_), .A2(new_n366_), .A3(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n367_), .B1(new_n362_), .B2(new_n366_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n344_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n370_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n372_), .A2(KEYINPUT81), .A3(new_n368_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n371_), .A2(new_n373_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n300_), .A2(new_n335_), .A3(new_n343_), .A4(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G71gat), .B(G99gat), .ZN(new_n376_));
  INV_X1    g175(.A(G176gat), .ZN(new_n377_));
  INV_X1    g176(.A(G169gat), .ZN(new_n378_));
  OAI21_X1  g177(.A(KEYINPUT22), .B1(new_n378_), .B2(KEYINPUT89), .ZN(new_n379_));
  OR2_X1    g178(.A1(new_n378_), .A2(KEYINPUT22), .ZN(new_n380_));
  OAI211_X1 g179(.A(new_n377_), .B(new_n379_), .C1(new_n380_), .C2(KEYINPUT89), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G169gat), .A2(G176gat), .ZN(new_n382_));
  AND2_X1   g181(.A1(KEYINPUT84), .A2(G183gat), .ZN(new_n383_));
  NOR2_X1   g182(.A1(KEYINPUT84), .A2(G183gat), .ZN(new_n384_));
  NOR3_X1   g183(.A1(new_n383_), .A2(new_n384_), .A3(G190gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G183gat), .A2(G190gat), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT23), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n381_), .B(new_n382_), .C1(new_n385_), .C2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT24), .ZN(new_n393_));
  NOR2_X1   g192(.A1(G169gat), .A2(G176gat), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n390_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n394_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n396_), .A2(KEYINPUT24), .A3(new_n382_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n395_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT25), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(G183gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(KEYINPUT86), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT86), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n402_), .A2(new_n399_), .A3(G183gat), .ZN(new_n403_));
  INV_X1    g202(.A(G190gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(KEYINPUT26), .ZN(new_n405_));
  AND3_X1   g204(.A1(new_n401_), .A2(new_n403_), .A3(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT26), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(G190gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT87), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT85), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n383_), .A2(new_n384_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n410_), .B1(new_n411_), .B2(KEYINPUT25), .ZN(new_n412_));
  NOR4_X1   g211(.A1(new_n383_), .A2(new_n384_), .A3(KEYINPUT85), .A4(new_n399_), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n406_), .B(new_n409_), .C1(new_n412_), .C2(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n398_), .B1(new_n414_), .B2(KEYINPUT88), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n406_), .A2(new_n409_), .ZN(new_n416_));
  OR2_X1    g215(.A1(new_n412_), .A2(new_n413_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT88), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n416_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n392_), .B1(new_n415_), .B2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(KEYINPUT30), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n420_), .A2(KEYINPUT30), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n376_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G227gat), .A2(G233gat), .ZN(new_n425_));
  INV_X1    g224(.A(G15gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n425_), .B(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(G43gat), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n420_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT30), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n376_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n432_), .A2(new_n433_), .A3(new_n421_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n424_), .A2(new_n429_), .A3(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n429_), .B1(new_n424_), .B2(new_n434_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G127gat), .B(G134gat), .ZN(new_n438_));
  INV_X1    g237(.A(G120gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(G113gat), .ZN(new_n440_));
  INV_X1    g239(.A(G113gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(G120gat), .ZN(new_n442_));
  AND3_X1   g241(.A1(new_n440_), .A2(new_n442_), .A3(KEYINPUT91), .ZN(new_n443_));
  AOI21_X1  g242(.A(KEYINPUT91), .B1(new_n440_), .B2(new_n442_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n438_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT91), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n441_), .A2(G120gat), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n439_), .A2(G113gat), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n446_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n438_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n440_), .A2(new_n442_), .A3(KEYINPUT91), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n449_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n445_), .A2(new_n452_), .A3(KEYINPUT92), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT92), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n454_), .B(new_n438_), .C1(new_n443_), .C2(new_n444_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(KEYINPUT31), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT93), .B1(new_n457_), .B2(KEYINPUT90), .ZN(new_n458_));
  NOR3_X1   g257(.A1(new_n436_), .A2(new_n437_), .A3(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n458_), .B1(KEYINPUT93), .B2(new_n457_), .ZN(new_n460_));
  NOR3_X1   g259(.A1(new_n422_), .A2(new_n376_), .A3(new_n423_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n433_), .B1(new_n432_), .B2(new_n421_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n428_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n460_), .B1(new_n463_), .B2(new_n435_), .ZN(new_n464_));
  AND2_X1   g263(.A1(G155gat), .A2(G162gat), .ZN(new_n465_));
  NOR2_X1   g264(.A1(G155gat), .A2(G162gat), .ZN(new_n466_));
  NOR3_X1   g265(.A1(new_n465_), .A2(new_n466_), .A3(KEYINPUT1), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G155gat), .A2(G162gat), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT1), .ZN(new_n469_));
  OAI22_X1  g268(.A1(new_n468_), .A2(new_n469_), .B1(G141gat), .B2(G148gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G155gat), .B(G162gat), .ZN(new_n471_));
  OAI22_X1  g270(.A1(new_n467_), .A2(new_n470_), .B1(KEYINPUT2), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G141gat), .A2(G148gat), .ZN(new_n473_));
  XOR2_X1   g272(.A(new_n473_), .B(KEYINPUT94), .Z(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(G141gat), .ZN(new_n476_));
  INV_X1    g275(.A(G148gat), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n476_), .A2(new_n477_), .A3(KEYINPUT95), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT3), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT3), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n480_), .A2(new_n476_), .A3(new_n477_), .A4(KEYINPUT95), .ZN(new_n481_));
  NAND3_X1  g280(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT96), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT96), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n484_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n479_), .A2(new_n481_), .A3(new_n483_), .A4(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n471_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n475_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n456_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT104), .ZN(new_n491_));
  AOI22_X1  g290(.A1(new_n472_), .A2(new_n474_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n445_), .A2(new_n452_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n491_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n490_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G225gat), .A2(G233gat), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n456_), .A2(new_n491_), .A3(new_n489_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n495_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n490_), .A2(KEYINPUT4), .ZN(new_n499_));
  AND2_X1   g298(.A1(new_n445_), .A2(new_n452_), .ZN(new_n500_));
  OAI21_X1  g299(.A(KEYINPUT104), .B1(new_n489_), .B2(new_n500_), .ZN(new_n501_));
  AOI22_X1  g300(.A1(new_n453_), .A2(new_n455_), .B1(new_n475_), .B2(new_n488_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n497_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n499_), .B1(new_n503_), .B2(KEYINPUT4), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n498_), .B1(new_n504_), .B2(new_n496_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G1gat), .B(G29gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(G85gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(KEYINPUT0), .B(G57gat), .ZN(new_n508_));
  XOR2_X1   g307(.A(new_n507_), .B(new_n508_), .Z(new_n509_));
  NAND2_X1  g308(.A1(new_n505_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n496_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT4), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n512_), .B1(new_n495_), .B2(new_n497_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n511_), .B1(new_n513_), .B2(new_n499_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n509_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n514_), .A2(new_n515_), .A3(new_n498_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n510_), .A2(new_n516_), .ZN(new_n517_));
  NOR3_X1   g316(.A1(new_n459_), .A2(new_n464_), .A3(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G8gat), .B(G36gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT18), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G64gat), .B(G92gat), .ZN(new_n521_));
  XOR2_X1   g320(.A(new_n520_), .B(new_n521_), .Z(new_n522_));
  INV_X1    g321(.A(KEYINPUT101), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n408_), .A2(new_n405_), .ZN(new_n524_));
  INV_X1    g323(.A(G183gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(KEYINPUT25), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n400_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT100), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n400_), .A2(new_n526_), .A3(KEYINPUT100), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n524_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n397_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n523_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  AND3_X1   g332(.A1(new_n400_), .A2(new_n526_), .A3(KEYINPUT100), .ZN(new_n534_));
  AOI21_X1  g333(.A(KEYINPUT100), .B1(new_n400_), .B2(new_n526_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  OAI211_X1 g335(.A(KEYINPUT101), .B(new_n397_), .C1(new_n536_), .C2(new_n524_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n533_), .A2(new_n537_), .A3(new_n395_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT22), .B(G169gat), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(new_n377_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(G183gat), .A2(G190gat), .ZN(new_n541_));
  OAI211_X1 g340(.A(new_n540_), .B(new_n382_), .C1(new_n390_), .C2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT102), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G197gat), .B(G204gat), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT21), .ZN(new_n545_));
  OR2_X1    g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(new_n545_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G211gat), .B(G218gat), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n546_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n549_));
  OR3_X1    g348(.A1(new_n544_), .A2(new_n548_), .A3(new_n545_), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n538_), .A2(new_n543_), .A3(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G226gat), .A2(G233gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT19), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT20), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n552_), .B(new_n556_), .C1(new_n420_), .C2(new_n551_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n549_), .A2(new_n550_), .ZN(new_n558_));
  AOI211_X1 g357(.A(new_n558_), .B(new_n392_), .C1(new_n415_), .C2(new_n419_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n551_), .B1(new_n538_), .B2(new_n543_), .ZN(new_n560_));
  NOR3_X1   g359(.A1(new_n559_), .A2(new_n560_), .A3(new_n555_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n554_), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n522_), .B(new_n557_), .C1(new_n561_), .C2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT103), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n560_), .A2(new_n555_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n415_), .A2(new_n419_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n567_), .A2(new_n551_), .A3(new_n391_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n566_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(new_n554_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n570_), .A2(KEYINPUT103), .A3(new_n522_), .A4(new_n557_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n522_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n562_), .B1(new_n566_), .B2(new_n568_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n557_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n572_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n565_), .A2(new_n571_), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT27), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n538_), .A2(new_n551_), .A3(new_n542_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(KEYINPUT20), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n551_), .B1(new_n567_), .B2(new_n391_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n554_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n538_), .A2(new_n543_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(new_n558_), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n583_), .A2(new_n568_), .A3(KEYINPUT20), .A4(new_n562_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n581_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(new_n572_), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n563_), .A2(KEYINPUT27), .ZN(new_n587_));
  AOI22_X1  g386(.A1(new_n576_), .A2(new_n577_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(KEYINPUT28), .B1(new_n489_), .B2(KEYINPUT29), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT28), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT29), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n492_), .A2(new_n590_), .A3(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G22gat), .B(G50gat), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n589_), .A2(new_n592_), .A3(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n593_), .B1(new_n589_), .B2(new_n592_), .ZN(new_n596_));
  OAI21_X1  g395(.A(KEYINPUT99), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(G228gat), .A2(G233gat), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n489_), .A2(KEYINPUT29), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT97), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT98), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n600_), .A2(new_n601_), .A3(new_n602_), .A4(new_n558_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n492_), .A2(new_n591_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n558_), .A2(new_n602_), .ZN(new_n605_));
  OAI21_X1  g404(.A(KEYINPUT97), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n599_), .B1(new_n603_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n589_), .A2(new_n592_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n593_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT99), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n611_), .A2(new_n612_), .A3(new_n594_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n603_), .A2(new_n606_), .A3(new_n599_), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n597_), .A2(new_n608_), .A3(new_n613_), .A4(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n611_), .A2(new_n594_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n614_), .ZN(new_n617_));
  OAI211_X1 g416(.A(KEYINPUT99), .B(new_n616_), .C1(new_n617_), .C2(new_n607_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n615_), .A2(new_n618_), .ZN(new_n619_));
  XOR2_X1   g418(.A(G78gat), .B(G106gat), .Z(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n615_), .A2(new_n618_), .A3(new_n620_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  AND3_X1   g424(.A1(new_n518_), .A2(new_n588_), .A3(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n522_), .A2(KEYINPUT32), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n585_), .A2(new_n628_), .ZN(new_n629_));
  OAI211_X1 g428(.A(new_n557_), .B(new_n627_), .C1(new_n561_), .C2(new_n562_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n631_), .B1(new_n516_), .B2(new_n510_), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n513_), .A2(new_n511_), .A3(new_n499_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n503_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n515_), .B1(new_n634_), .B2(new_n496_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT33), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n515_), .B1(new_n514_), .B2(new_n498_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT105), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n637_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n510_), .A2(KEYINPUT105), .A3(KEYINPUT33), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n636_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n565_), .A2(new_n571_), .A3(new_n575_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n632_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n517_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n624_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n576_), .A2(new_n577_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n587_), .A2(new_n586_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  OAI22_X1  g448(.A1(new_n644_), .A2(new_n624_), .B1(new_n646_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n459_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n464_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n626_), .B1(new_n650_), .B2(new_n653_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n351_), .B(new_n352_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n310_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n354_), .A2(new_n310_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT82), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n657_), .A2(new_n658_), .A3(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n655_), .A2(KEYINPUT82), .A3(new_n656_), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n660_), .A2(G229gat), .A3(G233gat), .A4(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n311_), .A2(new_n655_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(G229gat), .A2(G233gat), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n663_), .A2(new_n658_), .A3(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n662_), .A2(new_n665_), .ZN(new_n666_));
  XOR2_X1   g465(.A(G113gat), .B(G141gat), .Z(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT83), .ZN(new_n668_));
  XNOR2_X1  g467(.A(G169gat), .B(G197gat), .ZN(new_n669_));
  XOR2_X1   g468(.A(new_n668_), .B(new_n669_), .Z(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n666_), .A2(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n662_), .A2(new_n665_), .A3(new_n670_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n375_), .A2(new_n654_), .A3(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n517_), .B(KEYINPUT106), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n677_), .A2(new_n348_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n678_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT38), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n654_), .B1(new_n334_), .B2(new_n329_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n369_), .A2(new_n370_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n294_), .A2(KEYINPUT13), .A3(new_n295_), .ZN(new_n684_));
  AOI21_X1  g483(.A(KEYINPUT13), .B1(new_n294_), .B2(new_n295_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n674_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT107), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  OAI211_X1 g487(.A(KEYINPUT107), .B(new_n674_), .C1(new_n684_), .C2(new_n685_), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n681_), .A2(new_n683_), .A3(new_n688_), .A4(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(G1gat), .B1(new_n690_), .B2(new_n645_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n680_), .A2(new_n691_), .ZN(G1324gat));
  INV_X1    g491(.A(G8gat), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n676_), .A2(new_n693_), .A3(new_n649_), .ZN(new_n694_));
  OAI21_X1  g493(.A(G8gat), .B1(new_n690_), .B2(new_n588_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n695_), .A2(KEYINPUT39), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT39), .ZN(new_n697_));
  OAI211_X1 g496(.A(new_n697_), .B(G8gat), .C1(new_n690_), .C2(new_n588_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n694_), .B1(new_n696_), .B2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT40), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n700_), .B(new_n701_), .ZN(G1325gat));
  OAI21_X1  g501(.A(G15gat), .B1(new_n690_), .B2(new_n653_), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n703_), .A2(KEYINPUT41), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(KEYINPUT41), .ZN(new_n705_));
  INV_X1    g504(.A(new_n653_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n676_), .A2(new_n426_), .A3(new_n706_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT108), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n704_), .A2(new_n705_), .A3(new_n708_), .ZN(G1326gat));
  OAI21_X1  g508(.A(G22gat), .B1(new_n690_), .B2(new_n625_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT42), .ZN(new_n711_));
  INV_X1    g510(.A(G22gat), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n676_), .A2(new_n712_), .A3(new_n624_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(G1327gat));
  NAND2_X1  g513(.A1(new_n640_), .A2(new_n641_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n636_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n715_), .A2(new_n643_), .A3(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n632_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n624_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n649_), .A2(new_n646_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n653_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n626_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n374_), .A2(new_n336_), .ZN(new_n724_));
  AND4_X1   g523(.A1(new_n723_), .A2(new_n674_), .A3(new_n300_), .A4(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(G29gat), .B1(new_n725_), .B2(new_n517_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n374_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n688_), .A2(new_n689_), .A3(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n343_), .A2(new_n335_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT43), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n723_), .B(new_n729_), .C1(KEYINPUT109), .C2(new_n730_), .ZN(new_n731_));
  AOI211_X1 g530(.A(new_n339_), .B(new_n341_), .C1(new_n329_), .C2(new_n334_), .ZN(new_n732_));
  AND4_X1   g531(.A1(KEYINPUT77), .A2(new_n329_), .A3(KEYINPUT37), .A4(new_n334_), .ZN(new_n733_));
  OAI21_X1  g532(.A(KEYINPUT109), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n732_), .A2(new_n733_), .ZN(new_n735_));
  OAI211_X1 g534(.A(new_n734_), .B(KEYINPUT43), .C1(new_n735_), .C2(new_n654_), .ZN(new_n736_));
  AOI211_X1 g535(.A(KEYINPUT44), .B(new_n728_), .C1(new_n731_), .C2(new_n736_), .ZN(new_n737_));
  XOR2_X1   g536(.A(KEYINPUT110), .B(KEYINPUT44), .Z(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n736_), .A2(new_n731_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n728_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n739_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n737_), .A2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n677_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n744_), .A2(G29gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n726_), .B1(new_n743_), .B2(new_n745_), .ZN(G1328gat));
  NOR2_X1   g545(.A1(new_n737_), .A2(new_n742_), .ZN(new_n747_));
  OAI21_X1  g546(.A(G36gat), .B1(new_n747_), .B2(new_n588_), .ZN(new_n748_));
  INV_X1    g547(.A(G36gat), .ZN(new_n749_));
  OR2_X1    g548(.A1(new_n588_), .A2(KEYINPUT111), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n588_), .A2(KEYINPUT111), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n725_), .A2(new_n749_), .A3(new_n752_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(KEYINPUT112), .B(KEYINPUT45), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n753_), .B(new_n754_), .Z(new_n755_));
  NAND2_X1  g554(.A1(new_n748_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT46), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n748_), .A2(KEYINPUT46), .A3(new_n755_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(G1329gat));
  INV_X1    g559(.A(G43gat), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n653_), .A2(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n762_), .B1(new_n737_), .B2(new_n742_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT113), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  OAI211_X1 g564(.A(KEYINPUT113), .B(new_n762_), .C1(new_n737_), .C2(new_n742_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n725_), .A2(new_n706_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(new_n761_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n765_), .A2(new_n766_), .A3(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT47), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT47), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n765_), .A2(new_n771_), .A3(new_n766_), .A4(new_n768_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(G1330gat));
  AOI21_X1  g572(.A(G50gat), .B1(new_n725_), .B2(new_n624_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n624_), .A2(G50gat), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n743_), .B2(new_n775_), .ZN(G1331gat));
  NOR2_X1   g575(.A1(new_n300_), .A2(new_n674_), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n681_), .A2(new_n374_), .A3(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n778_), .A2(G57gat), .A3(new_n517_), .ZN(new_n779_));
  OR2_X1    g578(.A1(new_n779_), .A2(KEYINPUT114), .ZN(new_n780_));
  INV_X1    g579(.A(G57gat), .ZN(new_n781_));
  NOR3_X1   g580(.A1(new_n654_), .A2(new_n674_), .A3(new_n300_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n729_), .A2(new_n727_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n781_), .B1(new_n784_), .B2(new_n677_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n779_), .A2(KEYINPUT114), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n780_), .A2(new_n785_), .A3(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT115), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n787_), .B(new_n788_), .ZN(G1332gat));
  INV_X1    g588(.A(G64gat), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n790_), .B1(new_n778_), .B2(new_n752_), .ZN(new_n791_));
  XOR2_X1   g590(.A(new_n791_), .B(KEYINPUT48), .Z(new_n792_));
  INV_X1    g591(.A(new_n784_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n793_), .A2(new_n790_), .A3(new_n752_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(G1333gat));
  INV_X1    g594(.A(KEYINPUT49), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n778_), .A2(new_n706_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n796_), .B1(new_n797_), .B2(G71gat), .ZN(new_n798_));
  INV_X1    g597(.A(G71gat), .ZN(new_n799_));
  AOI211_X1 g598(.A(KEYINPUT49), .B(new_n799_), .C1(new_n778_), .C2(new_n706_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n706_), .A2(new_n799_), .ZN(new_n801_));
  OAI22_X1  g600(.A1(new_n798_), .A2(new_n800_), .B1(new_n784_), .B2(new_n801_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(KEYINPUT116), .ZN(G1334gat));
  INV_X1    g602(.A(G78gat), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(new_n778_), .B2(new_n624_), .ZN(new_n805_));
  XOR2_X1   g604(.A(new_n805_), .B(KEYINPUT50), .Z(new_n806_));
  NAND3_X1  g605(.A1(new_n793_), .A2(new_n804_), .A3(new_n624_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(G1335gat));
  NAND2_X1  g607(.A1(new_n777_), .A2(new_n727_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n809_), .B1(new_n736_), .B2(new_n731_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(G85gat), .B1(new_n811_), .B2(new_n645_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n782_), .A2(new_n724_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n814_), .A2(new_n259_), .A3(new_n744_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n812_), .A2(new_n815_), .ZN(G1336gat));
  INV_X1    g615(.A(new_n752_), .ZN(new_n817_));
  OAI21_X1  g616(.A(G92gat), .B1(new_n811_), .B2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n814_), .A2(new_n260_), .A3(new_n649_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(G1337gat));
  NAND3_X1  g619(.A1(new_n814_), .A2(new_n255_), .A3(new_n706_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n811_), .A2(new_n653_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n821_), .B1(new_n822_), .B2(new_n225_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n823_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n810_), .A2(new_n624_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n825_), .B1(new_n826_), .B2(G106gat), .ZN(new_n827_));
  AOI211_X1 g626(.A(KEYINPUT52), .B(new_n226_), .C1(new_n810_), .C2(new_n624_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n624_), .A2(new_n226_), .ZN(new_n829_));
  OAI22_X1  g628(.A1(new_n827_), .A2(new_n828_), .B1(new_n813_), .B2(new_n829_), .ZN(new_n830_));
  XNOR2_X1  g629(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n830_), .B(new_n832_), .ZN(G1339gat));
  NAND2_X1  g632(.A1(new_n674_), .A2(new_n293_), .ZN(new_n834_));
  XOR2_X1   g633(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n835_));
  NAND2_X1  g634(.A1(new_n273_), .A2(KEYINPUT55), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT55), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n267_), .A2(new_n837_), .A3(new_n272_), .A4(new_n270_), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n267_), .A2(new_n270_), .A3(new_n279_), .A4(new_n276_), .ZN(new_n839_));
  AOI22_X1  g638(.A1(new_n836_), .A2(new_n838_), .B1(new_n271_), .B2(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n835_), .B1(new_n840_), .B2(new_n289_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n836_), .A2(new_n838_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n839_), .A2(new_n271_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT56), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n289_), .A2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n834_), .B1(new_n841_), .B2(new_n847_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n660_), .A2(new_n661_), .A3(new_n664_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n664_), .B1(new_n354_), .B2(new_n310_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n670_), .B1(new_n850_), .B2(new_n663_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n851_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n673_), .A2(new_n852_), .ZN(new_n853_));
  AND3_X1   g652(.A1(new_n294_), .A2(new_n295_), .A3(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n336_), .B1(new_n848_), .B2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT57), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  OAI211_X1 g656(.A(KEYINPUT57), .B(new_n336_), .C1(new_n848_), .C2(new_n854_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n844_), .A2(KEYINPUT119), .A3(new_n846_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT119), .ZN(new_n860_));
  INV_X1    g659(.A(new_n846_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(new_n840_), .B2(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n845_), .B1(new_n840_), .B2(new_n289_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n859_), .A2(new_n862_), .A3(new_n863_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n853_), .A2(new_n293_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n864_), .A2(KEYINPUT58), .A3(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n729_), .ZN(new_n867_));
  AOI21_X1  g666(.A(KEYINPUT58), .B1(new_n864_), .B2(new_n865_), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n857_), .B(new_n858_), .C1(new_n867_), .C2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(KEYINPUT120), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n864_), .A2(new_n865_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT58), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n873_), .A2(new_n729_), .A3(new_n866_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT120), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n874_), .A2(new_n875_), .A3(new_n857_), .A4(new_n858_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n870_), .A2(new_n682_), .A3(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT54), .ZN(new_n878_));
  NAND4_X1  g677(.A1(new_n783_), .A2(new_n878_), .A3(new_n675_), .A4(new_n300_), .ZN(new_n879_));
  OAI21_X1  g678(.A(KEYINPUT54), .B1(new_n375_), .B2(new_n674_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n877_), .A2(new_n881_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n649_), .A2(new_n624_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n883_), .A2(new_n706_), .A3(new_n744_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n882_), .A2(KEYINPUT121), .A3(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT121), .ZN(new_n887_));
  AND2_X1   g686(.A1(new_n879_), .A2(new_n880_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n683_), .B1(new_n869_), .B2(KEYINPUT120), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n888_), .B1(new_n889_), .B2(new_n876_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n887_), .B1(new_n890_), .B2(new_n884_), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n886_), .A2(new_n891_), .A3(new_n441_), .A4(new_n674_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n869_), .A2(new_n727_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(new_n881_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT59), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n894_), .A2(new_n895_), .A3(new_n885_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n884_), .B1(new_n877_), .B2(new_n881_), .ZN(new_n897_));
  OAI211_X1 g696(.A(new_n674_), .B(new_n896_), .C1(new_n897_), .C2(new_n895_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n892_), .B1(new_n899_), .B2(new_n441_), .ZN(G1340gat));
  XNOR2_X1  g699(.A(KEYINPUT122), .B(G120gat), .ZN(new_n901_));
  OR2_X1    g700(.A1(new_n901_), .A2(KEYINPUT60), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n300_), .B2(KEYINPUT60), .ZN(new_n903_));
  NAND4_X1  g702(.A1(new_n886_), .A2(new_n891_), .A3(new_n902_), .A4(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n300_), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n905_), .B(new_n896_), .C1(new_n897_), .C2(new_n895_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n906_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n904_), .B1(new_n907_), .B2(new_n901_), .ZN(G1341gat));
  INV_X1    g707(.A(G127gat), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n886_), .A2(new_n891_), .A3(new_n374_), .ZN(new_n910_));
  AOI211_X1 g709(.A(KEYINPUT59), .B(new_n884_), .C1(new_n893_), .C2(new_n881_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n882_), .A2(new_n885_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n911_), .B1(new_n912_), .B2(KEYINPUT59), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n682_), .A2(new_n909_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(KEYINPUT123), .ZN(new_n915_));
  AOI22_X1  g714(.A1(new_n909_), .A2(new_n910_), .B1(new_n913_), .B2(new_n915_), .ZN(G1342gat));
  OAI21_X1  g715(.A(new_n896_), .B1(new_n897_), .B2(new_n895_), .ZN(new_n917_));
  OAI21_X1  g716(.A(G134gat), .B1(new_n917_), .B2(new_n735_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n336_), .A2(G134gat), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n886_), .A2(new_n891_), .A3(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n918_), .A2(new_n920_), .ZN(G1343gat));
  NOR4_X1   g720(.A1(new_n752_), .A2(new_n706_), .A3(new_n625_), .A4(new_n677_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n882_), .A2(new_n674_), .A3(new_n922_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g723(.A1(new_n882_), .A2(new_n905_), .A3(new_n922_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g725(.A1(new_n882_), .A2(new_n374_), .A3(new_n922_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(KEYINPUT61), .B(G155gat), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n927_), .B(new_n928_), .ZN(G1346gat));
  NOR2_X1   g728(.A1(new_n336_), .A2(G162gat), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n882_), .A2(new_n922_), .A3(new_n930_), .ZN(new_n931_));
  AND3_X1   g730(.A1(new_n882_), .A2(new_n729_), .A3(new_n922_), .ZN(new_n932_));
  INV_X1    g731(.A(G162gat), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n931_), .B1(new_n932_), .B2(new_n933_), .ZN(G1347gat));
  NOR3_X1   g733(.A1(new_n817_), .A2(new_n653_), .A3(new_n744_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(new_n625_), .ZN(new_n936_));
  INV_X1    g735(.A(new_n936_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n894_), .A2(new_n937_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n938_), .A2(KEYINPUT124), .ZN(new_n939_));
  INV_X1    g738(.A(KEYINPUT124), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n894_), .A2(new_n940_), .A3(new_n937_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n939_), .A2(new_n941_), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n942_), .A2(new_n539_), .A3(new_n674_), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n894_), .A2(new_n674_), .A3(new_n937_), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT62), .ZN(new_n945_));
  AND3_X1   g744(.A1(new_n944_), .A2(new_n945_), .A3(G169gat), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n945_), .B1(new_n944_), .B2(G169gat), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n943_), .B1(new_n946_), .B2(new_n947_), .ZN(G1348gat));
  NAND2_X1  g747(.A1(new_n942_), .A2(new_n905_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n890_), .A2(new_n624_), .ZN(new_n950_));
  AND3_X1   g749(.A1(new_n935_), .A2(G176gat), .A3(new_n905_), .ZN(new_n951_));
  AOI22_X1  g750(.A1(new_n949_), .A2(new_n377_), .B1(new_n950_), .B2(new_n951_), .ZN(G1349gat));
  NAND3_X1  g751(.A1(new_n950_), .A2(new_n374_), .A3(new_n935_), .ZN(new_n953_));
  NOR3_X1   g752(.A1(new_n682_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n954_));
  AOI22_X1  g753(.A1(new_n953_), .A2(new_n411_), .B1(new_n942_), .B2(new_n954_), .ZN(G1350gat));
  NOR2_X1   g754(.A1(new_n336_), .A2(new_n524_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n942_), .A2(new_n956_), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n735_), .B1(new_n939_), .B2(new_n941_), .ZN(new_n958_));
  OAI21_X1  g757(.A(new_n957_), .B1(new_n404_), .B2(new_n958_), .ZN(G1351gat));
  NOR3_X1   g758(.A1(new_n817_), .A2(new_n706_), .A3(new_n646_), .ZN(new_n960_));
  INV_X1    g759(.A(new_n960_), .ZN(new_n961_));
  NOR2_X1   g760(.A1(new_n890_), .A2(new_n961_), .ZN(new_n962_));
  AND3_X1   g761(.A1(new_n962_), .A2(G197gat), .A3(new_n674_), .ZN(new_n963_));
  AOI21_X1  g762(.A(G197gat), .B1(new_n962_), .B2(new_n674_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n963_), .A2(new_n964_), .ZN(G1352gat));
  NAND3_X1  g764(.A1(new_n882_), .A2(new_n905_), .A3(new_n960_), .ZN(new_n966_));
  XNOR2_X1  g765(.A(new_n966_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g766(.A(KEYINPUT125), .ZN(new_n968_));
  NOR3_X1   g767(.A1(new_n968_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n969_));
  AOI211_X1 g768(.A(new_n969_), .B(new_n682_), .C1(KEYINPUT63), .C2(G211gat), .ZN(new_n970_));
  NAND3_X1  g769(.A1(new_n882_), .A2(new_n960_), .A3(new_n970_), .ZN(new_n971_));
  OAI21_X1  g770(.A(new_n968_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n972_));
  XNOR2_X1  g771(.A(new_n972_), .B(KEYINPUT126), .ZN(new_n973_));
  XNOR2_X1  g772(.A(new_n971_), .B(new_n973_), .ZN(G1354gat));
  NAND2_X1  g773(.A1(new_n882_), .A2(new_n960_), .ZN(new_n975_));
  INV_X1    g774(.A(G218gat), .ZN(new_n976_));
  NOR3_X1   g775(.A1(new_n975_), .A2(new_n976_), .A3(new_n735_), .ZN(new_n977_));
  NOR3_X1   g776(.A1(new_n890_), .A2(new_n336_), .A3(new_n961_), .ZN(new_n978_));
  AOI21_X1  g777(.A(G218gat), .B1(new_n978_), .B2(KEYINPUT127), .ZN(new_n979_));
  INV_X1    g778(.A(KEYINPUT127), .ZN(new_n980_));
  OAI21_X1  g779(.A(new_n980_), .B1(new_n975_), .B2(new_n336_), .ZN(new_n981_));
  AOI21_X1  g780(.A(new_n977_), .B1(new_n979_), .B2(new_n981_), .ZN(G1355gat));
endmodule


