//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 0 0 0 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 0 0 0 0 0 1 1 1 1 1 0 1 1 0 0 1 1 0 1 0 1 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n694_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n745_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n848_, new_n849_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n861_, new_n863_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n910_, new_n911_, new_n912_,
    new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n927_, new_n929_, new_n930_, new_n931_, new_n932_, new_n934_,
    new_n935_, new_n936_;
  XNOR2_X1  g000(.A(G22gat), .B(G50gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XOR2_X1   g002(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n204_));
  NOR2_X1   g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206_));
  AOI21_X1  g005(.A(new_n205_), .B1(KEYINPUT1), .B2(new_n206_), .ZN(new_n207_));
  OR2_X1    g006(.A1(new_n206_), .A2(KEYINPUT1), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210_));
  INV_X1    g009(.A(G141gat), .ZN(new_n211_));
  INV_X1    g010(.A(G148gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n209_), .A2(new_n210_), .A3(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT88), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT87), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT85), .ZN(new_n218_));
  AND2_X1   g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  OAI211_X1 g018(.A(KEYINPUT85), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT86), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT2), .ZN(new_n223_));
  AND3_X1   g022(.A1(new_n210_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n222_), .B1(new_n210_), .B2(new_n223_), .ZN(new_n225_));
  OAI22_X1  g024(.A1(new_n219_), .A2(new_n221_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n210_), .A2(new_n223_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT84), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT3), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT83), .B1(G141gat), .B2(G148gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(KEYINPUT84), .A2(KEYINPUT3), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n231_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  NOR3_X1   g033(.A1(KEYINPUT83), .A2(G141gat), .A3(G148gat), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n228_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n216_), .B1(new_n226_), .B2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n210_), .A2(new_n223_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT86), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n210_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n217_), .A2(new_n218_), .ZN(new_n241_));
  AOI22_X1  g040(.A1(new_n239_), .A2(new_n240_), .B1(new_n241_), .B2(new_n220_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n235_), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n243_), .A2(new_n232_), .A3(new_n231_), .A4(new_n233_), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n242_), .A2(KEYINPUT87), .A3(new_n244_), .A4(new_n228_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n237_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n206_), .ZN(new_n247_));
  OR2_X1    g046(.A1(new_n247_), .A2(new_n205_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n215_), .B1(new_n246_), .B2(new_n249_), .ZN(new_n250_));
  AOI211_X1 g049(.A(KEYINPUT88), .B(new_n248_), .C1(new_n237_), .C2(new_n245_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n214_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(KEYINPUT89), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT89), .ZN(new_n254_));
  OAI211_X1 g053(.A(new_n254_), .B(new_n214_), .C1(new_n250_), .C2(new_n251_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT29), .ZN(new_n257_));
  AOI21_X1  g056(.A(KEYINPUT90), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT90), .ZN(new_n259_));
  AOI211_X1 g058(.A(new_n259_), .B(KEYINPUT29), .C1(new_n253_), .C2(new_n255_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n204_), .B1(new_n258_), .B2(new_n260_), .ZN(new_n261_));
  NOR3_X1   g060(.A1(new_n226_), .A2(new_n236_), .A3(new_n216_), .ZN(new_n262_));
  AND3_X1   g061(.A1(new_n231_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n227_), .B1(new_n263_), .B2(new_n243_), .ZN(new_n264_));
  AOI21_X1  g063(.A(KEYINPUT87), .B1(new_n264_), .B2(new_n242_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n249_), .B1(new_n262_), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(KEYINPUT88), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n246_), .A2(new_n215_), .A3(new_n249_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n254_), .B1(new_n269_), .B2(new_n214_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n255_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n257_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(new_n259_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n256_), .A2(KEYINPUT90), .A3(new_n257_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n204_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n273_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n203_), .B1(new_n261_), .B2(new_n276_), .ZN(new_n277_));
  AND3_X1   g076(.A1(new_n261_), .A2(new_n276_), .A3(new_n203_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n253_), .A2(KEYINPUT29), .A3(new_n255_), .ZN(new_n279_));
  INV_X1    g078(.A(G204gat), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n280_), .A2(G197gat), .ZN(new_n281_));
  INV_X1    g080(.A(G197gat), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n282_), .A2(G204gat), .ZN(new_n283_));
  OAI21_X1  g082(.A(KEYINPUT21), .B1(new_n281_), .B2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G211gat), .B(G218gat), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n283_), .B1(KEYINPUT93), .B2(new_n281_), .ZN(new_n286_));
  OR2_X1    g085(.A1(new_n281_), .A2(KEYINPUT93), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n284_), .B(new_n285_), .C1(new_n288_), .C2(KEYINPUT21), .ZN(new_n289_));
  INV_X1    g088(.A(new_n285_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n288_), .A2(KEYINPUT21), .A3(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n289_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(G233gat), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT92), .ZN(new_n295_));
  OR2_X1    g094(.A1(new_n295_), .A2(G228gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(G228gat), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n294_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n293_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n279_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(G78gat), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n257_), .B1(new_n269_), .B2(new_n214_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n298_), .B1(new_n302_), .B2(new_n293_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n300_), .A2(new_n301_), .A3(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n301_), .B1(new_n300_), .B2(new_n303_), .ZN(new_n306_));
  INV_X1    g105(.A(G106gat), .ZN(new_n307_));
  NOR3_X1   g106(.A1(new_n305_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n300_), .A2(new_n303_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(G78gat), .ZN(new_n310_));
  AOI21_X1  g109(.A(G106gat), .B1(new_n310_), .B2(new_n304_), .ZN(new_n311_));
  OAI22_X1  g110(.A1(new_n277_), .A2(new_n278_), .B1(new_n308_), .B2(new_n311_), .ZN(new_n312_));
  NOR3_X1   g111(.A1(new_n258_), .A2(new_n260_), .A3(new_n204_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n275_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n202_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n307_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n310_), .A2(G106gat), .A3(new_n304_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n261_), .A2(new_n276_), .A3(new_n203_), .ZN(new_n318_));
  NAND4_X1  g117(.A1(new_n315_), .A2(new_n316_), .A3(new_n317_), .A4(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n312_), .A2(new_n319_), .ZN(new_n320_));
  XOR2_X1   g119(.A(G127gat), .B(G134gat), .Z(new_n321_));
  XNOR2_X1  g120(.A(G113gat), .B(G120gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n253_), .A2(new_n255_), .A3(new_n323_), .ZN(new_n324_));
  OR2_X1    g123(.A1(new_n252_), .A2(new_n323_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G225gat), .A2(G233gat), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n324_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n324_), .A2(KEYINPUT4), .A3(new_n325_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT4), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n253_), .A2(new_n330_), .A3(new_n255_), .A4(new_n323_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n326_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n328_), .B1(new_n329_), .B2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G1gat), .B(G29gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(G85gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT0), .B(G57gat), .ZN(new_n338_));
  XOR2_X1   g137(.A(new_n337_), .B(new_n338_), .Z(new_n339_));
  NOR2_X1   g138(.A1(new_n335_), .A2(new_n339_), .ZN(new_n340_));
  AND3_X1   g139(.A1(new_n324_), .A2(KEYINPUT4), .A3(new_n325_), .ZN(new_n341_));
  OAI211_X1 g140(.A(new_n327_), .B(new_n339_), .C1(new_n341_), .C2(new_n333_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n340_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G183gat), .A2(G190gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT23), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n347_), .B1(G183gat), .B2(G190gat), .ZN(new_n348_));
  NOR2_X1   g147(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(G169gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT25), .B(G183gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT26), .B(G190gat), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G169gat), .A2(G176gat), .ZN(new_n356_));
  AOI22_X1  g155(.A1(new_n352_), .A2(new_n353_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  OR3_X1    g156(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n357_), .A2(new_n358_), .A3(new_n347_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n351_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n292_), .A2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT96), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n347_), .A2(new_n358_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT94), .ZN(new_n364_));
  XOR2_X1   g163(.A(KEYINPUT22), .B(G169gat), .Z(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT95), .ZN(new_n366_));
  INV_X1    g165(.A(G176gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  AND2_X1   g167(.A1(new_n348_), .A2(new_n356_), .ZN(new_n369_));
  AOI22_X1  g168(.A1(new_n364_), .A2(new_n357_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(new_n293_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G226gat), .A2(G233gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT19), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n362_), .A2(new_n371_), .A3(KEYINPUT20), .A4(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n370_), .A2(new_n293_), .ZN(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT20), .B1(new_n292_), .B2(new_n360_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n373_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n375_), .A2(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G8gat), .B(G36gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT18), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G64gat), .B(G92gat), .ZN(new_n382_));
  XOR2_X1   g181(.A(new_n381_), .B(new_n382_), .Z(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n379_), .A2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n375_), .A2(new_n383_), .A3(new_n378_), .ZN(new_n386_));
  AND2_X1   g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  OR2_X1    g186(.A1(new_n387_), .A2(KEYINPUT27), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT98), .B(KEYINPUT20), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n389_), .B1(new_n370_), .B2(new_n293_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n374_), .B1(new_n362_), .B2(new_n390_), .ZN(new_n391_));
  NOR3_X1   g190(.A1(new_n376_), .A2(new_n373_), .A3(new_n377_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n384_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n393_), .A2(KEYINPUT27), .A3(new_n386_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n388_), .A2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G71gat), .B(G99gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(G43gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n360_), .B(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G227gat), .A2(G233gat), .ZN(new_n399_));
  INV_X1    g198(.A(G15gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT30), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n398_), .B(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT81), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(KEYINPUT82), .ZN(new_n405_));
  XOR2_X1   g204(.A(new_n323_), .B(KEYINPUT31), .Z(new_n406_));
  OAI21_X1  g205(.A(new_n406_), .B1(new_n403_), .B2(KEYINPUT81), .ZN(new_n407_));
  AND2_X1   g206(.A1(new_n405_), .A2(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n405_), .A2(new_n407_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NOR4_X1   g209(.A1(new_n320_), .A2(new_n345_), .A3(new_n395_), .A4(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n395_), .ZN(new_n412_));
  AND4_X1   g211(.A1(new_n317_), .A2(new_n315_), .A3(new_n316_), .A4(new_n318_), .ZN(new_n413_));
  AOI22_X1  g212(.A1(new_n315_), .A2(new_n318_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n344_), .B(new_n412_), .C1(new_n413_), .C2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT33), .ZN(new_n416_));
  AND2_X1   g215(.A1(new_n342_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n339_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n418_), .A2(new_n416_), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n327_), .B(new_n419_), .C1(new_n341_), .C2(new_n333_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n324_), .A2(new_n325_), .A3(new_n332_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n331_), .A2(new_n326_), .ZN(new_n422_));
  OAI211_X1 g221(.A(new_n418_), .B(new_n421_), .C1(new_n341_), .C2(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n420_), .A2(new_n423_), .A3(new_n387_), .ZN(new_n424_));
  OAI21_X1  g223(.A(KEYINPUT97), .B1(new_n417_), .B2(new_n424_), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n423_), .A2(new_n387_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n342_), .A2(new_n416_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT97), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n426_), .A2(new_n427_), .A3(new_n428_), .A4(new_n420_), .ZN(new_n429_));
  OAI211_X1 g228(.A(KEYINPUT32), .B(new_n383_), .C1(new_n391_), .C2(new_n392_), .ZN(new_n430_));
  OR2_X1    g229(.A1(new_n430_), .A2(KEYINPUT99), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n383_), .A2(KEYINPUT32), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n375_), .A2(new_n378_), .A3(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n430_), .A2(KEYINPUT99), .ZN(new_n434_));
  AND3_X1   g233(.A1(new_n431_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n435_), .B1(new_n340_), .B2(new_n343_), .ZN(new_n436_));
  AND3_X1   g235(.A1(new_n425_), .A2(new_n429_), .A3(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n415_), .B1(new_n437_), .B2(new_n320_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n411_), .B1(new_n438_), .B2(new_n410_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G1gat), .B(G8gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT74), .ZN(new_n441_));
  INV_X1    g240(.A(G22gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n400_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G15gat), .A2(G22gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(G1gat), .A2(G8gat), .ZN(new_n445_));
  AOI22_X1  g244(.A1(new_n443_), .A2(new_n444_), .B1(KEYINPUT14), .B2(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n441_), .B(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G29gat), .B(G36gat), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n449_), .A2(KEYINPUT71), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n449_), .A2(KEYINPUT71), .ZN(new_n451_));
  XOR2_X1   g250(.A(G43gat), .B(G50gat), .Z(new_n452_));
  OR3_X1    g251(.A1(new_n450_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n452_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n454_));
  AND2_X1   g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  XOR2_X1   g254(.A(KEYINPUT72), .B(KEYINPUT15), .Z(new_n456_));
  AND2_X1   g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n455_), .A2(new_n456_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n448_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT79), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n455_), .B(new_n456_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT79), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n461_), .A2(new_n462_), .A3(new_n448_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G229gat), .A2(G233gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n455_), .A2(KEYINPUT78), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n453_), .A2(new_n454_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT78), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n465_), .A2(new_n447_), .A3(new_n468_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n460_), .A2(new_n463_), .A3(new_n464_), .A4(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n465_), .A2(new_n468_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(new_n448_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(new_n469_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n464_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n470_), .A2(KEYINPUT80), .A3(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n476_), .B1(KEYINPUT80), .B2(new_n470_), .ZN(new_n477_));
  XOR2_X1   g276(.A(G113gat), .B(G141gat), .Z(new_n478_));
  XNOR2_X1  g277(.A(G169gat), .B(G197gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n477_), .B(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n439_), .A2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G190gat), .B(G218gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G134gat), .B(G162gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  XOR2_X1   g285(.A(new_n486_), .B(KEYINPUT36), .Z(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  XOR2_X1   g287(.A(G85gat), .B(G92gat), .Z(new_n489_));
  NAND2_X1  g288(.A1(G99gat), .A2(G106gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT6), .ZN(new_n491_));
  OAI21_X1  g290(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n492_));
  OR2_X1    g291(.A1(new_n492_), .A2(KEYINPUT64), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(KEYINPUT64), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n491_), .A2(new_n493_), .A3(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(G99gat), .ZN(new_n496_));
  AND3_X1   g295(.A1(new_n496_), .A2(new_n307_), .A3(KEYINPUT65), .ZN(new_n497_));
  AOI21_X1  g296(.A(KEYINPUT65), .B1(new_n496_), .B2(new_n307_), .ZN(new_n498_));
  NOR3_X1   g297(.A1(new_n497_), .A2(new_n498_), .A3(KEYINPUT7), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n489_), .B1(new_n495_), .B2(new_n499_), .ZN(new_n500_));
  OR2_X1    g299(.A1(new_n500_), .A2(KEYINPUT8), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(KEYINPUT8), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  XOR2_X1   g302(.A(KEYINPUT10), .B(G99gat), .Z(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(new_n307_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n489_), .A2(KEYINPUT9), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT9), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n507_), .A2(G85gat), .A3(G92gat), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n505_), .A2(new_n506_), .A3(new_n491_), .A4(new_n508_), .ZN(new_n509_));
  XOR2_X1   g308(.A(new_n509_), .B(KEYINPUT69), .Z(new_n510_));
  NAND2_X1  g309(.A1(new_n503_), .A2(new_n510_), .ZN(new_n511_));
  AND2_X1   g310(.A1(new_n461_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G232gat), .A2(G233gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT34), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT35), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n503_), .A2(new_n509_), .ZN(new_n518_));
  OAI22_X1  g317(.A1(new_n518_), .A2(new_n466_), .B1(KEYINPUT35), .B2(new_n514_), .ZN(new_n519_));
  OR3_X1    g318(.A1(new_n512_), .A2(new_n517_), .A3(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n517_), .B1(new_n512_), .B2(new_n519_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n488_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n486_), .A2(KEYINPUT36), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n520_), .A2(new_n521_), .A3(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n523_), .A2(KEYINPUT37), .A3(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  OR2_X1    g326(.A1(new_n522_), .A2(KEYINPUT73), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n522_), .A2(KEYINPUT73), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n528_), .A2(new_n529_), .A3(new_n525_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT37), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n527_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G57gat), .B(G64gat), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT67), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT11), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT68), .ZN(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT66), .B(G71gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(G78gat), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n537_), .A2(new_n538_), .A3(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n538_), .B1(new_n537_), .B2(new_n540_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n535_), .A2(new_n536_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NOR3_X1   g343(.A1(new_n541_), .A2(new_n542_), .A3(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n537_), .A2(new_n540_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT68), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n537_), .A2(new_n538_), .A3(new_n540_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n543_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n518_), .B1(new_n545_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT12), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n544_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n547_), .A2(new_n548_), .A3(new_n543_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n551_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  AOI22_X1  g353(.A1(new_n550_), .A2(new_n551_), .B1(new_n554_), .B2(new_n511_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n509_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n556_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n557_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G230gat), .A2(G233gat), .ZN(new_n559_));
  AOI21_X1  g358(.A(KEYINPUT70), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  AND3_X1   g359(.A1(new_n558_), .A2(KEYINPUT70), .A3(new_n559_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n555_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n550_), .A2(new_n558_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n563_), .A2(G230gat), .A3(G233gat), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G120gat), .B(G148gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT5), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G176gat), .B(G204gat), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n567_), .B(new_n568_), .Z(new_n569_));
  NAND2_X1  g368(.A1(new_n565_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n569_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n562_), .A2(new_n564_), .A3(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n574_), .A2(KEYINPUT13), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(KEYINPUT13), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G231gat), .A2(G233gat), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n447_), .B(new_n577_), .Z(new_n578_));
  NAND2_X1  g377(.A1(new_n552_), .A2(new_n553_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G127gat), .B(G155gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT16), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G183gat), .B(G211gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(KEYINPUT75), .B(KEYINPUT17), .Z(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT76), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n580_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT77), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n584_), .B(KEYINPUT17), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n580_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n590_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n532_), .A2(new_n575_), .A3(new_n576_), .A4(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n483_), .A2(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT100), .ZN(new_n598_));
  INV_X1    g397(.A(G1gat), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n598_), .A2(new_n599_), .A3(new_n345_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT38), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n320_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n410_), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n603_), .A2(new_n344_), .A3(new_n412_), .A4(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n425_), .A2(new_n429_), .A3(new_n436_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n395_), .B1(new_n312_), .B2(new_n319_), .ZN(new_n607_));
  AOI22_X1  g406(.A1(new_n603_), .A2(new_n606_), .B1(new_n607_), .B2(new_n344_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n605_), .B1(new_n608_), .B2(new_n604_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n575_), .A2(new_n576_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NOR3_X1   g410(.A1(new_n611_), .A2(new_n482_), .A3(new_n593_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n609_), .A2(new_n530_), .A3(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(G1gat), .B1(new_n613_), .B2(new_n344_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n600_), .A2(new_n601_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n602_), .A2(new_n614_), .A3(new_n615_), .ZN(G1324gat));
  INV_X1    g415(.A(G8gat), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n598_), .A2(new_n617_), .A3(new_n395_), .ZN(new_n618_));
  OAI21_X1  g417(.A(G8gat), .B1(new_n613_), .B2(new_n412_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT39), .ZN(new_n620_));
  XNOR2_X1  g419(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n618_), .A2(new_n620_), .A3(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n621_), .B1(new_n618_), .B2(new_n620_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n623_), .A2(new_n624_), .ZN(G1325gat));
  OAI21_X1  g424(.A(G15gat), .B1(new_n613_), .B2(new_n410_), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n626_), .B(KEYINPUT41), .Z(new_n627_));
  INV_X1    g426(.A(new_n597_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n628_), .A2(new_n400_), .A3(new_n604_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n627_), .A2(new_n629_), .ZN(G1326gat));
  INV_X1    g429(.A(KEYINPUT102), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n320_), .B(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(G22gat), .B1(new_n613_), .B2(new_n633_), .ZN(new_n634_));
  XOR2_X1   g433(.A(KEYINPUT103), .B(KEYINPUT42), .Z(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n628_), .A2(new_n442_), .A3(new_n632_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(G1327gat));
  NOR2_X1   g437(.A1(new_n594_), .A2(new_n530_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n611_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n483_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(G29gat), .B1(new_n643_), .B2(new_n345_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n610_), .A2(new_n481_), .A3(new_n593_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT43), .ZN(new_n647_));
  INV_X1    g446(.A(new_n532_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n603_), .A2(new_n606_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n604_), .B1(new_n649_), .B2(new_n415_), .ZN(new_n650_));
  OAI211_X1 g449(.A(new_n647_), .B(new_n648_), .C1(new_n650_), .C2(new_n411_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n647_), .B1(new_n609_), .B2(new_n648_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n646_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT105), .ZN(new_n655_));
  XNOR2_X1  g454(.A(KEYINPUT104), .B(KEYINPUT44), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n654_), .A2(new_n655_), .A3(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(KEYINPUT43), .B1(new_n439_), .B2(new_n532_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n645_), .B1(new_n659_), .B2(new_n651_), .ZN(new_n660_));
  OAI21_X1  g459(.A(KEYINPUT105), .B1(new_n660_), .B2(new_n656_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n658_), .A2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n659_), .A2(new_n651_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n663_), .A2(KEYINPUT44), .A3(new_n646_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n345_), .A2(G29gat), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n644_), .B1(new_n666_), .B2(new_n667_), .ZN(G1328gat));
  INV_X1    g467(.A(KEYINPUT46), .ZN(new_n669_));
  INV_X1    g468(.A(G36gat), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n671_));
  AOI211_X1 g470(.A(new_n671_), .B(new_n645_), .C1(new_n659_), .C2(new_n651_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n672_), .A2(new_n412_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n670_), .B1(new_n662_), .B2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n395_), .A2(new_n670_), .ZN(new_n675_));
  OR3_X1    g474(.A1(new_n642_), .A2(KEYINPUT45), .A3(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(KEYINPUT45), .B1(new_n642_), .B2(new_n675_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n669_), .B1(new_n674_), .B2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n664_), .A2(new_n395_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n681_), .B1(new_n661_), .B2(new_n658_), .ZN(new_n682_));
  OAI211_X1 g481(.A(KEYINPUT46), .B(new_n678_), .C1(new_n682_), .C2(new_n670_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n680_), .A2(new_n683_), .ZN(G1329gat));
  NAND2_X1  g483(.A1(new_n604_), .A2(G43gat), .ZN(new_n685_));
  AOI211_X1 g484(.A(new_n672_), .B(new_n685_), .C1(new_n658_), .C2(new_n661_), .ZN(new_n686_));
  INV_X1    g485(.A(G43gat), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n687_), .B1(new_n642_), .B2(new_n410_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(KEYINPUT47), .B1(new_n686_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT47), .ZN(new_n691_));
  OAI211_X1 g490(.A(new_n691_), .B(new_n688_), .C1(new_n665_), .C2(new_n685_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n690_), .A2(new_n692_), .ZN(G1330gat));
  OAI21_X1  g492(.A(G50gat), .B1(new_n665_), .B2(new_n603_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n633_), .A2(G50gat), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT106), .Z(new_n696_));
  OAI21_X1  g495(.A(new_n694_), .B1(new_n642_), .B2(new_n696_), .ZN(G1331gat));
  NOR3_X1   g496(.A1(new_n610_), .A2(new_n481_), .A3(new_n593_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n609_), .A2(new_n530_), .A3(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(KEYINPUT108), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT108), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n609_), .A2(new_n701_), .A3(new_n530_), .A4(new_n698_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n700_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(G57gat), .B1(new_n704_), .B2(new_n344_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT107), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n706_), .B1(new_n439_), .B2(new_n481_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n609_), .A2(KEYINPUT107), .A3(new_n482_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NOR3_X1   g508(.A1(new_n610_), .A2(new_n593_), .A3(new_n648_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(G57gat), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n711_), .A2(new_n712_), .A3(new_n345_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n705_), .A2(new_n713_), .ZN(G1332gat));
  INV_X1    g513(.A(G64gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n703_), .B2(new_n395_), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT48), .Z(new_n717_));
  NAND3_X1  g516(.A1(new_n711_), .A2(new_n715_), .A3(new_n395_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1333gat));
  INV_X1    g518(.A(G71gat), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n711_), .A2(new_n720_), .A3(new_n604_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n703_), .B2(new_n604_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(KEYINPUT109), .B(KEYINPUT49), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n722_), .A2(new_n723_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n721_), .B1(new_n724_), .B2(new_n725_), .ZN(G1334gat));
  NAND3_X1  g525(.A1(new_n711_), .A2(new_n301_), .A3(new_n632_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n700_), .A2(new_n632_), .A3(new_n702_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT50), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n728_), .A2(new_n729_), .A3(G78gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n728_), .B2(G78gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n727_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT110), .ZN(G1335gat));
  NOR2_X1   g532(.A1(new_n610_), .A2(new_n640_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n709_), .A2(KEYINPUT111), .A3(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(KEYINPUT111), .B1(new_n709_), .B2(new_n734_), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(G85gat), .B1(new_n738_), .B2(new_n345_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n611_), .A2(new_n482_), .A3(new_n593_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(new_n659_), .B2(new_n651_), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n741_), .B(KEYINPUT112), .Z(new_n742_));
  AND2_X1   g541(.A1(new_n345_), .A2(G85gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n739_), .B1(new_n742_), .B2(new_n743_), .ZN(G1336gat));
  AOI21_X1  g543(.A(G92gat), .B1(new_n738_), .B2(new_n395_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n395_), .A2(G92gat), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT113), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n745_), .B1(new_n742_), .B2(new_n747_), .ZN(G1337gat));
  INV_X1    g547(.A(new_n741_), .ZN(new_n749_));
  OAI21_X1  g548(.A(G99gat), .B1(new_n749_), .B2(new_n410_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n736_), .A2(new_n737_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n604_), .A2(new_n504_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n750_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(KEYINPUT51), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT51), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n755_), .B(new_n750_), .C1(new_n751_), .C2(new_n752_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n756_), .ZN(G1338gat));
  OAI211_X1 g556(.A(new_n307_), .B(new_n320_), .C1(new_n736_), .C2(new_n737_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT52), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n741_), .A2(new_n320_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n760_), .B2(G106gat), .ZN(new_n761_));
  AOI211_X1 g560(.A(KEYINPUT52), .B(new_n307_), .C1(new_n741_), .C2(new_n320_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n758_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT53), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT53), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n758_), .B(new_n765_), .C1(new_n761_), .C2(new_n762_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(G1339gat));
  NOR3_X1   g566(.A1(new_n344_), .A2(new_n395_), .A3(new_n410_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n555_), .A2(new_n558_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n769_), .A2(G230gat), .A3(G233gat), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT114), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n558_), .A2(new_n559_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT70), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n558_), .A2(KEYINPUT70), .A3(new_n559_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n771_), .B1(new_n776_), .B2(new_n555_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT55), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n770_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  AOI211_X1 g578(.A(new_n771_), .B(KEYINPUT55), .C1(new_n776_), .C2(new_n555_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n569_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT56), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n460_), .A2(new_n463_), .A3(new_n474_), .A4(new_n469_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n480_), .B1(new_n473_), .B2(new_n464_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n785_), .B1(new_n477_), .B2(new_n480_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT56), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n787_), .B(new_n569_), .C1(new_n779_), .C2(new_n780_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n782_), .A2(new_n572_), .A3(new_n786_), .A4(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT58), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n532_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  OR2_X1    g590(.A1(new_n791_), .A2(KEYINPUT116), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n789_), .A2(new_n790_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n793_), .B1(new_n791_), .B2(KEYINPUT116), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n782_), .A2(new_n481_), .A3(new_n572_), .A4(new_n788_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n786_), .A2(new_n573_), .A3(KEYINPUT115), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(KEYINPUT115), .B1(new_n786_), .B2(new_n573_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n796_), .A2(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT57), .B1(new_n801_), .B2(new_n530_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT57), .ZN(new_n803_));
  INV_X1    g602(.A(new_n530_), .ZN(new_n804_));
  AOI211_X1 g603(.A(new_n803_), .B(new_n804_), .C1(new_n796_), .C2(new_n800_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n802_), .A2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n594_), .B1(new_n795_), .B2(new_n806_), .ZN(new_n807_));
  OR3_X1    g606(.A1(new_n595_), .A2(KEYINPUT54), .A3(new_n481_), .ZN(new_n808_));
  OAI21_X1  g607(.A(KEYINPUT54), .B1(new_n595_), .B2(new_n481_), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n603_), .B(new_n768_), .C1(new_n807_), .C2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(G113gat), .B1(new_n812_), .B2(new_n481_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT59), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n811_), .A2(new_n814_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n791_), .A2(KEYINPUT116), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT116), .ZN(new_n817_));
  AOI211_X1 g616(.A(new_n817_), .B(new_n532_), .C1(new_n789_), .C2(new_n790_), .ZN(new_n818_));
  NOR3_X1   g617(.A1(new_n816_), .A2(new_n818_), .A3(new_n793_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n801_), .A2(new_n530_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n803_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n801_), .A2(KEYINPUT57), .A3(new_n530_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n593_), .B1(new_n819_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n810_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n826_), .A2(KEYINPUT59), .A3(new_n603_), .A4(new_n768_), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n815_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n481_), .A2(G113gat), .ZN(new_n830_));
  XOR2_X1   g629(.A(new_n830_), .B(KEYINPUT117), .Z(new_n831_));
  AOI21_X1  g630(.A(new_n813_), .B1(new_n829_), .B2(new_n831_), .ZN(G1340gat));
  OAI21_X1  g631(.A(G120gat), .B1(new_n828_), .B2(new_n610_), .ZN(new_n833_));
  INV_X1    g632(.A(G120gat), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n834_), .B1(new_n610_), .B2(KEYINPUT60), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n835_), .B1(KEYINPUT60), .B2(new_n834_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n833_), .B1(new_n811_), .B2(new_n836_), .ZN(G1341gat));
  INV_X1    g636(.A(G127gat), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n838_), .B1(new_n811_), .B2(new_n593_), .ZN(new_n839_));
  NOR3_X1   g638(.A1(new_n593_), .A2(KEYINPUT118), .A3(new_n838_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n840_), .B1(KEYINPUT118), .B2(new_n838_), .ZN(new_n841_));
  OAI211_X1 g640(.A(KEYINPUT119), .B(new_n839_), .C1(new_n828_), .C2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT119), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n841_), .B1(new_n815_), .B2(new_n827_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n839_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n843_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n842_), .A2(new_n846_), .ZN(G1342gat));
  OAI21_X1  g646(.A(G134gat), .B1(new_n828_), .B2(new_n532_), .ZN(new_n848_));
  OR3_X1    g647(.A1(new_n811_), .A2(G134gat), .A3(new_n530_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(G1343gat));
  NAND2_X1  g649(.A1(new_n789_), .A2(new_n790_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n851_), .A2(KEYINPUT116), .A3(new_n648_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n793_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n821_), .B(new_n822_), .C1(new_n854_), .C2(new_n816_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n810_), .B1(new_n855_), .B2(new_n593_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n856_), .A2(new_n604_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n857_), .A2(new_n345_), .A3(new_n607_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n858_), .A2(new_n482_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(new_n211_), .ZN(G1344gat));
  NOR2_X1   g659(.A1(new_n858_), .A2(new_n610_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(new_n212_), .ZN(G1345gat));
  NOR2_X1   g661(.A1(new_n858_), .A2(new_n593_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(KEYINPUT61), .B(G155gat), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n863_), .B(new_n865_), .ZN(G1346gat));
  OAI21_X1  g665(.A(G162gat), .B1(new_n858_), .B2(new_n532_), .ZN(new_n867_));
  OR2_X1    g666(.A1(new_n530_), .A2(G162gat), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n867_), .B1(new_n858_), .B2(new_n868_), .ZN(G1347gat));
  NOR2_X1   g668(.A1(new_n345_), .A2(new_n412_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n604_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n632_), .A2(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n826_), .A2(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(G169gat), .B1(new_n873_), .B2(new_n482_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT120), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  OAI211_X1 g675(.A(KEYINPUT120), .B(G169gat), .C1(new_n873_), .C2(new_n482_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n876_), .A2(KEYINPUT62), .A3(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT62), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n874_), .A2(new_n875_), .A3(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT121), .ZN(new_n881_));
  INV_X1    g680(.A(new_n872_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n881_), .B1(new_n856_), .B2(new_n882_), .ZN(new_n883_));
  OAI211_X1 g682(.A(KEYINPUT121), .B(new_n872_), .C1(new_n807_), .C2(new_n810_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n481_), .A2(new_n366_), .ZN(new_n886_));
  XOR2_X1   g685(.A(new_n886_), .B(KEYINPUT122), .Z(new_n887_));
  NAND2_X1  g686(.A1(new_n885_), .A2(new_n887_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n878_), .A2(new_n880_), .A3(new_n888_), .ZN(G1348gat));
  INV_X1    g688(.A(new_n871_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n826_), .A2(new_n603_), .A3(new_n890_), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n891_), .A2(new_n367_), .A3(new_n610_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n885_), .A2(new_n611_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT123), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n893_), .A2(new_n894_), .A3(new_n367_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n610_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n896_));
  OAI21_X1  g695(.A(KEYINPUT123), .B1(new_n896_), .B2(G176gat), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n892_), .B1(new_n895_), .B2(new_n897_), .ZN(G1349gat));
  INV_X1    g697(.A(G183gat), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n899_), .B1(new_n891_), .B2(new_n593_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n352_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n594_), .A2(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n903_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n904_));
  OAI21_X1  g703(.A(KEYINPUT124), .B1(new_n901_), .B2(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n904_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT124), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n906_), .A2(new_n907_), .A3(new_n900_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n905_), .A2(new_n908_), .ZN(G1350gat));
  NAND3_X1  g708(.A1(new_n885_), .A2(new_n353_), .A3(new_n804_), .ZN(new_n910_));
  AOI21_X1  g709(.A(KEYINPUT121), .B1(new_n826_), .B2(new_n872_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n884_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n648_), .B1(new_n911_), .B2(new_n912_), .ZN(new_n913_));
  AOI21_X1  g712(.A(KEYINPUT125), .B1(new_n913_), .B2(G190gat), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n532_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT125), .ZN(new_n916_));
  INV_X1    g715(.A(G190gat), .ZN(new_n917_));
  NOR3_X1   g716(.A1(new_n915_), .A2(new_n916_), .A3(new_n917_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n910_), .B1(new_n914_), .B2(new_n918_), .ZN(G1351gat));
  AND2_X1   g718(.A1(new_n870_), .A2(new_n320_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n857_), .A2(new_n920_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n921_), .ZN(new_n922_));
  OAI211_X1 g721(.A(new_n922_), .B(new_n481_), .C1(KEYINPUT126), .C2(G197gat), .ZN(new_n923_));
  XNOR2_X1  g722(.A(KEYINPUT126), .B(G197gat), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n924_), .B1(new_n921_), .B2(new_n482_), .ZN(new_n925_));
  AND2_X1   g724(.A1(new_n923_), .A2(new_n925_), .ZN(G1352gat));
  NOR2_X1   g725(.A1(new_n921_), .A2(new_n610_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(new_n280_), .ZN(G1353gat));
  XOR2_X1   g727(.A(KEYINPUT63), .B(G211gat), .Z(new_n929_));
  NAND3_X1  g728(.A1(new_n922_), .A2(new_n594_), .A3(new_n929_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n931_), .B1(new_n921_), .B2(new_n593_), .ZN(new_n932_));
  AND2_X1   g731(.A1(new_n930_), .A2(new_n932_), .ZN(G1354gat));
  AOI21_X1  g732(.A(G218gat), .B1(new_n922_), .B2(new_n804_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n648_), .A2(G218gat), .ZN(new_n935_));
  XOR2_X1   g734(.A(new_n935_), .B(KEYINPUT127), .Z(new_n936_));
  AOI21_X1  g735(.A(new_n934_), .B1(new_n922_), .B2(new_n936_), .ZN(G1355gat));
endmodule


