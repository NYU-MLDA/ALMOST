//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 0 1 1 0 0 0 1 0 0 1 1 1 0 1 0 1 0 1 0 0 0 1 0 0 1 0 1 1 0 0 0 0 0 0 1 1 1 1 0 0 0 0 1 0 0 0 0 1 1 0 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n667_, new_n668_, new_n669_, new_n670_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n727_, new_n728_, new_n729_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n736_, new_n737_, new_n738_, new_n739_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n861_, new_n862_,
    new_n863_, new_n865_, new_n866_, new_n867_, new_n868_, new_n870_,
    new_n871_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n922_, new_n923_, new_n925_,
    new_n926_, new_n927_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n936_, new_n937_, new_n938_, new_n939_;
  NAND2_X1  g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202_));
  INV_X1    g001(.A(G169gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT22), .ZN(new_n204_));
  AOI21_X1  g003(.A(G176gat), .B1(new_n204_), .B2(KEYINPUT83), .ZN(new_n205_));
  OAI21_X1  g004(.A(new_n205_), .B1(KEYINPUT83), .B2(new_n204_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT84), .ZN(new_n207_));
  OR2_X1    g006(.A1(new_n207_), .A2(KEYINPUT22), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(KEYINPUT22), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n203_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n202_), .B1(new_n206_), .B2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT85), .ZN(new_n212_));
  OR2_X1    g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT23), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n214_), .B(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(G183gat), .A2(G190gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n218_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n213_), .A2(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221_));
  XOR2_X1   g020(.A(new_n221_), .B(KEYINPUT82), .Z(new_n222_));
  NAND3_X1  g021(.A1(new_n222_), .A2(KEYINPUT24), .A3(new_n202_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT25), .B(G183gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT26), .B(G190gat), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n216_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n223_), .B(new_n226_), .C1(KEYINPUT24), .C2(new_n222_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n220_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(G204gat), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT91), .B1(new_n229_), .B2(G197gat), .ZN(new_n230_));
  INV_X1    g029(.A(G197gat), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n230_), .B1(new_n231_), .B2(G204gat), .ZN(new_n232_));
  NOR3_X1   g031(.A1(new_n229_), .A2(KEYINPUT91), .A3(G197gat), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT21), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G211gat), .B(G218gat), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT92), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n236_), .B1(G197gat), .B2(new_n229_), .ZN(new_n237_));
  NOR3_X1   g036(.A1(new_n231_), .A2(KEYINPUT92), .A3(G204gat), .ZN(new_n238_));
  OAI22_X1  g037(.A1(new_n237_), .A2(new_n238_), .B1(G197gat), .B2(new_n229_), .ZN(new_n239_));
  OAI211_X1 g038(.A(new_n234_), .B(new_n235_), .C1(new_n239_), .C2(KEYINPUT21), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT21), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT93), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n241_), .B1(new_n235_), .B2(new_n242_), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n243_), .B(new_n239_), .C1(new_n242_), .C2(new_n235_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n240_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n228_), .A2(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(KEYINPUT19), .A2(G226gat), .A3(G233gat), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(KEYINPUT19), .B1(G226gat), .B2(G233gat), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n218_), .B1(G169gat), .B2(G176gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT22), .B(G169gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT97), .ZN(new_n254_));
  INV_X1    g053(.A(G176gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n252_), .A2(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT96), .B(KEYINPUT24), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n258_), .B1(G169gat), .B2(G176gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n222_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n258_), .A2(new_n221_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n260_), .A2(new_n226_), .A3(new_n261_), .ZN(new_n262_));
  AND2_X1   g061(.A1(new_n257_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n245_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n246_), .A2(KEYINPUT20), .A3(new_n251_), .A4(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT20), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n257_), .A2(new_n262_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n267_), .B1(new_n268_), .B2(new_n245_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n220_), .A2(new_n264_), .A3(new_n227_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n250_), .B(KEYINPUT95), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G8gat), .B(G36gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT18), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G64gat), .B(G92gat), .ZN(new_n276_));
  XOR2_X1   g075(.A(new_n275_), .B(new_n276_), .Z(new_n277_));
  NAND3_X1  g076(.A1(new_n266_), .A2(new_n273_), .A3(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n272_), .ZN(new_n279_));
  AND3_X1   g078(.A1(new_n269_), .A2(new_n270_), .A3(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n264_), .B1(new_n263_), .B2(KEYINPUT103), .ZN(new_n281_));
  AND3_X1   g080(.A1(new_n257_), .A2(KEYINPUT103), .A3(new_n262_), .ZN(new_n282_));
  OAI211_X1 g081(.A(new_n246_), .B(KEYINPUT20), .C1(new_n281_), .C2(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n280_), .B1(new_n283_), .B2(new_n250_), .ZN(new_n284_));
  OAI211_X1 g083(.A(KEYINPUT27), .B(new_n278_), .C1(new_n284_), .C2(new_n277_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT27), .ZN(new_n286_));
  OAI211_X1 g085(.A(KEYINPUT20), .B(new_n251_), .C1(new_n268_), .C2(new_n245_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n287_), .B1(new_n245_), .B2(new_n228_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n279_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n277_), .ZN(new_n290_));
  NOR3_X1   g089(.A1(new_n288_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n277_), .B1(new_n266_), .B2(new_n273_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n286_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(G155gat), .A2(G162gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT89), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G155gat), .A2(G162gat), .ZN(new_n296_));
  AND2_X1   g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G141gat), .A2(G148gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT2), .ZN(new_n299_));
  OR2_X1    g098(.A1(G141gat), .A2(G148gat), .ZN(new_n300_));
  OR2_X1    g099(.A1(new_n300_), .A2(KEYINPUT3), .ZN(new_n301_));
  OAI21_X1  g100(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n302_));
  OR2_X1    g101(.A1(new_n302_), .A2(KEYINPUT90), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(KEYINPUT90), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n299_), .A2(new_n301_), .A3(new_n303_), .A4(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n297_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n296_), .A2(KEYINPUT1), .ZN(new_n307_));
  OR2_X1    g106(.A1(new_n296_), .A2(KEYINPUT1), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n295_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n300_), .A2(new_n298_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n306_), .A2(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n264_), .B1(new_n312_), .B2(KEYINPUT29), .ZN(new_n313_));
  AOI22_X1  g112(.A1(new_n297_), .A2(new_n305_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT29), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  AND2_X1   g115(.A1(new_n316_), .A2(KEYINPUT28), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n316_), .A2(KEYINPUT28), .ZN(new_n318_));
  OR3_X1    g117(.A1(new_n313_), .A2(new_n317_), .A3(new_n318_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n313_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G78gat), .B(G106gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT94), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G228gat), .A2(G233gat), .ZN(new_n324_));
  XOR2_X1   g123(.A(new_n323_), .B(new_n324_), .Z(new_n325_));
  XOR2_X1   g124(.A(G22gat), .B(G50gat), .Z(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n321_), .A2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n319_), .A2(new_n320_), .A3(new_n327_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n285_), .A2(new_n293_), .A3(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT105), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G71gat), .B(G99gat), .ZN(new_n334_));
  XOR2_X1   g133(.A(new_n334_), .B(G43gat), .Z(new_n335_));
  NAND2_X1  g134(.A1(new_n228_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G227gat), .A2(G233gat), .ZN(new_n337_));
  INV_X1    g136(.A(G15gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT30), .ZN(new_n340_));
  INV_X1    g139(.A(new_n335_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n220_), .A2(new_n227_), .A3(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n336_), .A2(new_n340_), .A3(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n340_), .B1(new_n336_), .B2(new_n342_), .ZN(new_n345_));
  OAI21_X1  g144(.A(KEYINPUT87), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G127gat), .B(G134gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT86), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G113gat), .B(G120gat), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  OR2_X1    g150(.A1(new_n347_), .A2(KEYINPUT86), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n347_), .A2(KEYINPUT86), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n352_), .A2(new_n353_), .A3(new_n349_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n351_), .A2(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT31), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n346_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n345_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT87), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n358_), .A2(new_n359_), .A3(new_n343_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n357_), .B(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G225gat), .A2(G233gat), .ZN(new_n362_));
  AND2_X1   g161(.A1(new_n351_), .A2(new_n354_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n363_), .A2(KEYINPUT4), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n362_), .B1(new_n364_), .B2(new_n312_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n363_), .A2(KEYINPUT98), .A3(new_n314_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT98), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n355_), .B1(new_n312_), .B2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n366_), .A2(new_n368_), .A3(KEYINPUT4), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n365_), .A2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n366_), .A2(new_n368_), .A3(new_n362_), .ZN(new_n371_));
  XOR2_X1   g170(.A(G1gat), .B(G29gat), .Z(new_n372_));
  XNOR2_X1  g171(.A(G57gat), .B(G85gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n372_), .B(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n370_), .A2(new_n371_), .A3(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n377_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT105), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n285_), .A2(new_n293_), .A3(new_n331_), .A4(new_n382_), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n333_), .A2(new_n361_), .A3(new_n381_), .A4(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT106), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n290_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n387_));
  AND2_X1   g186(.A1(new_n366_), .A2(new_n368_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n362_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n389_), .B1(new_n364_), .B2(new_n312_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(new_n369_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n390_), .A2(new_n392_), .A3(new_n376_), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n387_), .A2(new_n278_), .A3(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT100), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT33), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n395_), .B1(new_n378_), .B2(new_n396_), .ZN(new_n397_));
  AOI22_X1  g196(.A1(new_n362_), .A2(new_n388_), .B1(new_n365_), .B2(new_n369_), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n398_), .A2(KEYINPUT100), .A3(KEYINPUT33), .A4(new_n377_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT101), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n398_), .A2(new_n401_), .A3(new_n377_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n378_), .A2(KEYINPUT101), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n402_), .A2(new_n403_), .A3(new_n396_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n394_), .A2(new_n400_), .A3(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(KEYINPUT102), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT102), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n394_), .A2(new_n400_), .A3(new_n404_), .A4(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n277_), .A2(KEYINPUT32), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n284_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n266_), .A2(new_n273_), .A3(new_n409_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n411_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n410_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n406_), .A2(new_n408_), .A3(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(new_n331_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT104), .ZN(new_n417_));
  INV_X1    g216(.A(new_n331_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n413_), .B1(new_n405_), .B2(KEYINPUT102), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n418_), .B1(new_n419_), .B2(new_n408_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT104), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n285_), .A2(new_n293_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n424_), .A2(new_n418_), .A3(new_n381_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n417_), .A2(new_n422_), .A3(new_n425_), .ZN(new_n426_));
  XOR2_X1   g225(.A(new_n361_), .B(KEYINPUT88), .Z(new_n427_));
  AOI21_X1  g226(.A(new_n386_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G1gat), .B(G8gat), .ZN(new_n429_));
  XOR2_X1   g228(.A(new_n429_), .B(KEYINPUT79), .Z(new_n430_));
  XNOR2_X1  g229(.A(G15gat), .B(G22gat), .ZN(new_n431_));
  INV_X1    g230(.A(G1gat), .ZN(new_n432_));
  INV_X1    g231(.A(G8gat), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT14), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n431_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n430_), .A2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n429_), .B(KEYINPUT79), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(new_n435_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(G36gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(G29gat), .ZN(new_n443_));
  INV_X1    g242(.A(G29gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(G36gat), .ZN(new_n445_));
  AOI21_X1  g244(.A(KEYINPUT72), .B1(new_n443_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n443_), .A2(new_n445_), .A3(KEYINPUT72), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G43gat), .B(G50gat), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n447_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n449_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n448_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n451_), .B1(new_n452_), .B2(new_n446_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n450_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT15), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n450_), .A2(new_n453_), .A3(KEYINPUT15), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n441_), .A2(new_n458_), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n450_), .A2(new_n453_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n440_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G229gat), .A2(G233gat), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n459_), .A2(new_n461_), .A3(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT81), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n437_), .A2(new_n454_), .A3(new_n439_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n461_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n462_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n464_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  AOI211_X1 g267(.A(KEYINPUT81), .B(new_n462_), .C1(new_n461_), .C2(new_n465_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n463_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  XOR2_X1   g269(.A(G113gat), .B(G141gat), .Z(new_n471_));
  XNOR2_X1  g270(.A(G169gat), .B(G197gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  XOR2_X1   g272(.A(new_n470_), .B(new_n473_), .Z(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n428_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(G99gat), .ZN(new_n477_));
  INV_X1    g276(.A(G106gat), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n477_), .A2(new_n478_), .A3(KEYINPUT65), .A4(KEYINPUT7), .ZN(new_n479_));
  NAND2_X1  g278(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n480_), .B1(G99gat), .B2(G106gat), .ZN(new_n481_));
  NOR2_X1   g280(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n479_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT6), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT64), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT64), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT6), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n485_), .A2(new_n487_), .A3(G99gat), .A4(G106gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G99gat), .A2(G106gat), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n486_), .A2(KEYINPUT6), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n484_), .A2(KEYINPUT64), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n489_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n483_), .A2(new_n488_), .A3(new_n492_), .ZN(new_n493_));
  AND2_X1   g292(.A1(G85gat), .A2(G92gat), .ZN(new_n494_));
  NOR2_X1   g293(.A1(G85gat), .A2(G92gat), .ZN(new_n495_));
  OAI21_X1  g294(.A(KEYINPUT67), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(G85gat), .ZN(new_n497_));
  INV_X1    g296(.A(G92gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT67), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G85gat), .A2(G92gat), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n499_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  AND2_X1   g301(.A1(new_n496_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n493_), .A2(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n496_), .A2(new_n502_), .A3(KEYINPUT66), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT8), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n504_), .A2(new_n507_), .ZN(new_n508_));
  AND2_X1   g307(.A1(new_n492_), .A2(new_n488_), .ZN(new_n509_));
  OR2_X1    g308(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n510_), .A2(new_n478_), .A3(new_n511_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n501_), .A2(KEYINPUT9), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n494_), .A2(new_n495_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n513_), .B1(new_n514_), .B2(KEYINPUT9), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n509_), .A2(new_n512_), .A3(new_n515_), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n493_), .B(new_n503_), .C1(KEYINPUT66), .C2(KEYINPUT8), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n508_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT68), .ZN(new_n519_));
  INV_X1    g318(.A(G64gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(G57gat), .ZN(new_n521_));
  INV_X1    g320(.A(G57gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(G64gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT11), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G71gat), .B(G78gat), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n519_), .B1(new_n526_), .B2(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(KEYINPUT11), .B1(new_n521_), .B2(new_n523_), .ZN(new_n530_));
  NOR3_X1   g329(.A1(new_n530_), .A2(KEYINPUT68), .A3(new_n527_), .ZN(new_n531_));
  OAI22_X1  g330(.A1(new_n529_), .A2(new_n531_), .B1(new_n525_), .B2(new_n524_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n526_), .A2(new_n519_), .A3(new_n528_), .ZN(new_n533_));
  OAI21_X1  g332(.A(KEYINPUT68), .B1(new_n530_), .B2(new_n527_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n524_), .A2(new_n525_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n533_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n532_), .A2(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(KEYINPUT12), .B1(new_n518_), .B2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n518_), .A2(new_n537_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G230gat), .A2(G233gat), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT70), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n515_), .A2(new_n512_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n492_), .A2(new_n488_), .ZN(new_n544_));
  OAI21_X1  g343(.A(KEYINPUT69), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT69), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n509_), .A2(new_n546_), .A3(new_n512_), .A4(new_n515_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n508_), .A2(new_n517_), .A3(new_n545_), .A4(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT12), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n549_), .B1(new_n532_), .B2(new_n536_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n542_), .B1(new_n548_), .B2(new_n550_), .ZN(new_n551_));
  AND3_X1   g350(.A1(new_n548_), .A2(new_n550_), .A3(new_n542_), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n540_), .B(new_n541_), .C1(new_n551_), .C2(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n518_), .B(new_n537_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n541_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n553_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G120gat), .B(G148gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT5), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G176gat), .B(G204gat), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n559_), .B(new_n560_), .Z(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n557_), .B(new_n562_), .ZN(new_n563_));
  XOR2_X1   g362(.A(new_n563_), .B(KEYINPUT13), .Z(new_n564_));
  NAND2_X1  g363(.A1(new_n548_), .A2(new_n458_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G232gat), .A2(G233gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT34), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(KEYINPUT35), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT71), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  OR2_X1    g369(.A1(new_n567_), .A2(KEYINPUT35), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n508_), .A2(new_n460_), .A3(new_n516_), .A4(new_n517_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n565_), .A2(new_n570_), .A3(new_n571_), .A4(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT75), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n572_), .A2(new_n571_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n569_), .B1(new_n548_), .B2(new_n458_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n577_), .A2(new_n578_), .A3(KEYINPUT75), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n575_), .A2(new_n579_), .ZN(new_n580_));
  XOR2_X1   g379(.A(G190gat), .B(G218gat), .Z(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT74), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G134gat), .B(G162gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n584_), .A2(KEYINPUT36), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT73), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n565_), .A2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n548_), .A2(new_n458_), .A3(KEYINPUT73), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n587_), .A2(new_n588_), .A3(new_n577_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(new_n569_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n580_), .A2(new_n585_), .A3(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT76), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n580_), .A2(new_n590_), .A3(KEYINPUT76), .A4(new_n585_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT37), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT77), .ZN(new_n597_));
  AND3_X1   g396(.A1(new_n577_), .A2(new_n578_), .A3(KEYINPUT75), .ZN(new_n598_));
  AOI21_X1  g397(.A(KEYINPUT75), .B1(new_n577_), .B2(new_n578_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n576_), .B1(new_n586_), .B2(new_n565_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n570_), .B1(new_n601_), .B2(new_n588_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n597_), .B1(new_n600_), .B2(new_n602_), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n584_), .B(KEYINPUT36), .Z(new_n604_));
  NAND3_X1  g403(.A1(new_n580_), .A2(KEYINPUT77), .A3(new_n590_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n603_), .A2(new_n604_), .A3(new_n605_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n595_), .A2(new_n596_), .A3(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n580_), .A2(new_n590_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(new_n604_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n596_), .B1(new_n595_), .B2(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(KEYINPUT78), .B1(new_n607_), .B2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(G231gat), .A2(G233gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n537_), .B(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(new_n441_), .ZN(new_n614_));
  XOR2_X1   g413(.A(G127gat), .B(G155gat), .Z(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT16), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G183gat), .B(G211gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT17), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n614_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT80), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n618_), .A2(new_n619_), .ZN(new_n624_));
  NOR3_X1   g423(.A1(new_n614_), .A2(new_n620_), .A3(new_n624_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n595_), .A2(new_n606_), .A3(new_n596_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT78), .ZN(new_n628_));
  AOI22_X1  g427(.A1(new_n593_), .A2(new_n594_), .B1(new_n608_), .B2(new_n604_), .ZN(new_n629_));
  OAI211_X1 g428(.A(new_n627_), .B(new_n628_), .C1(new_n596_), .C2(new_n629_), .ZN(new_n630_));
  AND4_X1   g429(.A1(new_n564_), .A2(new_n611_), .A3(new_n626_), .A4(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n476_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT107), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n381_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n634_), .A2(new_n432_), .A3(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT38), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n425_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n639_));
  AOI211_X1 g438(.A(KEYINPUT104), .B(new_n418_), .C1(new_n419_), .C2(new_n408_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n427_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n384_), .B(KEYINPUT106), .ZN(new_n642_));
  AOI22_X1  g441(.A1(new_n641_), .A2(new_n642_), .B1(new_n595_), .B2(new_n606_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n564_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n626_), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n644_), .A2(new_n645_), .A3(new_n475_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n643_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  OAI21_X1  g447(.A(G1gat), .B1(new_n648_), .B2(new_n381_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n636_), .A2(new_n637_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n638_), .A2(new_n649_), .A3(new_n650_), .ZN(G1324gat));
  NOR2_X1   g450(.A1(new_n424_), .A2(G8gat), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n634_), .A2(new_n652_), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n643_), .A2(KEYINPUT108), .A3(new_n423_), .A4(new_n646_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n654_), .A2(G8gat), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT39), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n643_), .A2(new_n423_), .A3(new_n646_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT108), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  AND3_X1   g458(.A1(new_n655_), .A2(new_n656_), .A3(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n656_), .B1(new_n655_), .B2(new_n659_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n653_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT40), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  OAI211_X1 g463(.A(new_n653_), .B(KEYINPUT40), .C1(new_n660_), .C2(new_n661_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1325gat));
  INV_X1    g465(.A(new_n427_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n338_), .B1(new_n647_), .B2(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT41), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n634_), .A2(new_n338_), .A3(new_n667_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(G1326gat));
  INV_X1    g470(.A(G22gat), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n331_), .B(KEYINPUT109), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n672_), .B1(new_n647_), .B2(new_n673_), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n674_), .B(KEYINPUT42), .Z(new_n675_));
  NAND3_X1  g474(.A1(new_n634_), .A2(new_n672_), .A3(new_n673_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1327gat));
  NAND2_X1  g476(.A1(new_n595_), .A2(new_n606_), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n626_), .A2(new_n678_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n644_), .A2(new_n679_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n476_), .A2(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n681_), .A2(new_n444_), .A3(new_n635_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n611_), .A2(new_n630_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(KEYINPUT43), .B1(new_n428_), .B2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n641_), .A2(new_n642_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n686_), .A2(new_n687_), .A3(new_n683_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n685_), .A2(new_n688_), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n644_), .A2(new_n475_), .A3(new_n626_), .ZN(new_n690_));
  AOI21_X1  g489(.A(KEYINPUT44), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n689_), .A2(KEYINPUT44), .A3(new_n690_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n692_), .A2(new_n635_), .A3(new_n693_), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n694_), .A2(KEYINPUT110), .A3(G29gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(KEYINPUT110), .B1(new_n694_), .B2(G29gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n682_), .B1(new_n695_), .B2(new_n696_), .ZN(G1328gat));
  NAND4_X1  g496(.A1(new_n476_), .A2(new_n442_), .A3(new_n423_), .A4(new_n680_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT45), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n700_));
  INV_X1    g499(.A(new_n690_), .ZN(new_n701_));
  AOI211_X1 g500(.A(new_n700_), .B(new_n701_), .C1(new_n685_), .C2(new_n688_), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n691_), .A2(new_n702_), .A3(new_n424_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n699_), .B1(new_n703_), .B2(new_n442_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT46), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  OAI211_X1 g505(.A(KEYINPUT46), .B(new_n699_), .C1(new_n703_), .C2(new_n442_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(G1329gat));
  AOI21_X1  g507(.A(G43gat), .B1(new_n681_), .B2(new_n667_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n691_), .A2(new_n702_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n361_), .A2(G43gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n709_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT47), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n712_), .B(new_n713_), .ZN(G1330gat));
  INV_X1    g513(.A(G50gat), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n673_), .A2(new_n715_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT111), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n681_), .A2(new_n717_), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n691_), .A2(new_n702_), .A3(new_n331_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n718_), .B1(new_n719_), .B2(new_n715_), .ZN(G1331gat));
  AND4_X1   g519(.A1(new_n475_), .A2(new_n643_), .A3(new_n644_), .A4(new_n626_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n522_), .B1(new_n721_), .B2(new_n635_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n683_), .A2(new_n645_), .ZN(new_n723_));
  AND4_X1   g522(.A1(new_n686_), .A2(new_n475_), .A3(new_n644_), .A4(new_n723_), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n724_), .A2(new_n522_), .A3(new_n635_), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n722_), .A2(new_n725_), .ZN(G1332gat));
  AOI21_X1  g525(.A(new_n520_), .B1(new_n721_), .B2(new_n423_), .ZN(new_n727_));
  XOR2_X1   g526(.A(new_n727_), .B(KEYINPUT48), .Z(new_n728_));
  NAND3_X1  g527(.A1(new_n724_), .A2(new_n520_), .A3(new_n423_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(G1333gat));
  INV_X1    g529(.A(G71gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n731_), .B1(new_n721_), .B2(new_n667_), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT49), .Z(new_n733_));
  NAND3_X1  g532(.A1(new_n724_), .A2(new_n731_), .A3(new_n667_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(G1334gat));
  INV_X1    g534(.A(G78gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n736_), .B1(new_n721_), .B2(new_n673_), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n737_), .B(KEYINPUT50), .Z(new_n738_));
  NAND3_X1  g537(.A1(new_n724_), .A2(new_n736_), .A3(new_n673_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(G1335gat));
  NOR4_X1   g539(.A1(new_n428_), .A2(new_n474_), .A3(new_n564_), .A4(new_n679_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n741_), .A2(new_n497_), .A3(new_n635_), .ZN(new_n742_));
  NOR3_X1   g541(.A1(new_n564_), .A2(new_n474_), .A3(new_n626_), .ZN(new_n743_));
  NOR3_X1   g542(.A1(new_n428_), .A2(KEYINPUT43), .A3(new_n684_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n687_), .B1(new_n686_), .B2(new_n683_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n743_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(KEYINPUT112), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT112), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n689_), .A2(new_n748_), .A3(new_n743_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n381_), .B1(new_n747_), .B2(new_n749_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n742_), .B1(new_n750_), .B2(new_n497_), .ZN(G1336gat));
  NAND3_X1  g550(.A1(new_n741_), .A2(new_n498_), .A3(new_n423_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n424_), .B1(new_n747_), .B2(new_n749_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n752_), .B1(new_n753_), .B2(new_n498_), .ZN(G1337gat));
  NAND4_X1  g553(.A1(new_n741_), .A2(new_n361_), .A3(new_n510_), .A4(new_n511_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n427_), .B1(new_n747_), .B2(new_n749_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n755_), .B1(new_n756_), .B2(new_n477_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(KEYINPUT51), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n759_), .B(new_n755_), .C1(new_n756_), .C2(new_n477_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(G1338gat));
  NAND3_X1  g560(.A1(new_n741_), .A2(new_n478_), .A3(new_n418_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n689_), .A2(new_n418_), .A3(new_n743_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT113), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n478_), .B1(new_n764_), .B2(KEYINPUT52), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n764_), .A2(KEYINPUT52), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n763_), .A2(new_n765_), .A3(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n763_), .B2(new_n765_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n762_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT53), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT53), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n771_), .B(new_n762_), .C1(new_n767_), .C2(new_n768_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(G1339gat));
  NAND2_X1  g572(.A1(new_n631_), .A2(new_n475_), .ZN(new_n774_));
  OAI21_X1  g573(.A(KEYINPUT114), .B1(new_n774_), .B2(KEYINPUT54), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT54), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n776_), .B1(new_n631_), .B2(new_n475_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n611_), .A2(new_n564_), .A3(new_n626_), .A4(new_n630_), .ZN(new_n779_));
  NOR4_X1   g578(.A1(new_n779_), .A2(KEYINPUT114), .A3(KEYINPUT54), .A4(new_n474_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n775_), .A2(new_n778_), .A3(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n473_), .B1(new_n466_), .B2(new_n462_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n459_), .A2(new_n461_), .A3(new_n467_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT116), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n463_), .B(new_n473_), .C1(new_n468_), .C2(new_n469_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT116), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n783_), .A2(new_n784_), .A3(new_n788_), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n786_), .A2(new_n787_), .A3(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n553_), .A2(new_n556_), .A3(new_n562_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT118), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n790_), .A2(new_n791_), .A3(KEYINPUT118), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT55), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n553_), .A2(new_n797_), .A3(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n552_), .A2(new_n551_), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n538_), .A2(new_n539_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n555_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n548_), .A2(new_n550_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(KEYINPUT70), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n548_), .A2(new_n550_), .A3(new_n542_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n807_), .A2(KEYINPUT55), .A3(new_n541_), .A4(new_n540_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n803_), .A2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n797_), .B1(new_n553_), .B2(new_n798_), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n800_), .A2(new_n809_), .A3(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT56), .ZN(new_n812_));
  NOR3_X1   g611(.A1(new_n811_), .A2(new_n812_), .A3(new_n562_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n553_), .A2(new_n798_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT115), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n815_), .A2(new_n799_), .A3(new_n808_), .A4(new_n803_), .ZN(new_n816_));
  AOI21_X1  g615(.A(KEYINPUT56), .B1(new_n816_), .B2(new_n561_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n796_), .B1(new_n813_), .B2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT58), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n796_), .B(KEYINPUT58), .C1(new_n813_), .C2(new_n817_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n683_), .A2(new_n820_), .A3(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n474_), .A2(new_n791_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n812_), .B1(new_n811_), .B2(new_n562_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n816_), .A2(KEYINPUT56), .A3(new_n561_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n823_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n790_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n563_), .A2(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n678_), .B1(new_n826_), .B2(new_n828_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(KEYINPUT117), .B(KEYINPUT57), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  OAI211_X1 g630(.A(KEYINPUT57), .B(new_n678_), .C1(new_n826_), .C2(new_n828_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n822_), .A2(new_n831_), .A3(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n645_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n782_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT59), .ZN(new_n836_));
  AND4_X1   g635(.A1(new_n635_), .A2(new_n333_), .A3(new_n361_), .A4(new_n383_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n835_), .A2(new_n836_), .A3(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT119), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n626_), .B1(new_n833_), .B2(new_n839_), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n822_), .A2(new_n831_), .A3(KEYINPUT119), .A4(new_n832_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n782_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n843_), .A2(new_n837_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n838_), .B1(new_n844_), .B2(new_n836_), .ZN(new_n845_));
  OAI21_X1  g644(.A(G113gat), .B1(new_n845_), .B2(new_n475_), .ZN(new_n846_));
  INV_X1    g645(.A(G113gat), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n844_), .A2(new_n847_), .A3(new_n474_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n848_), .ZN(G1340gat));
  NOR2_X1   g648(.A1(new_n564_), .A2(KEYINPUT60), .ZN(new_n850_));
  MUX2_X1   g649(.A(new_n850_), .B(KEYINPUT60), .S(G120gat), .Z(new_n851_));
  NAND2_X1  g650(.A1(new_n844_), .A2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT120), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n852_), .B(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(G120gat), .B1(new_n845_), .B2(new_n564_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(G1341gat));
  OAI21_X1  g655(.A(G127gat), .B1(new_n845_), .B2(new_n645_), .ZN(new_n857_));
  INV_X1    g656(.A(G127gat), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n844_), .A2(new_n858_), .A3(new_n626_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n859_), .ZN(G1342gat));
  OAI21_X1  g659(.A(G134gat), .B1(new_n845_), .B2(new_n684_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n678_), .A2(G134gat), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n844_), .A2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n863_), .ZN(G1343gat));
  NOR3_X1   g663(.A1(new_n423_), .A2(new_n331_), .A3(new_n381_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n843_), .A2(new_n427_), .A3(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n474_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(G141gat), .ZN(G1344gat));
  NOR2_X1   g668(.A1(new_n866_), .A2(new_n564_), .ZN(new_n870_));
  XOR2_X1   g669(.A(KEYINPUT121), .B(G148gat), .Z(new_n871_));
  XNOR2_X1  g670(.A(new_n870_), .B(new_n871_), .ZN(G1345gat));
  NAND4_X1  g671(.A1(new_n843_), .A2(new_n427_), .A3(new_n626_), .A4(new_n865_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n873_), .A2(KEYINPUT122), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n873_), .A2(KEYINPUT122), .ZN(new_n875_));
  XNOR2_X1  g674(.A(KEYINPUT61), .B(G155gat), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  OR3_X1    g676(.A1(new_n874_), .A2(new_n875_), .A3(new_n877_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1346gat));
  OAI21_X1  g679(.A(G162gat), .B1(new_n866_), .B2(new_n684_), .ZN(new_n881_));
  OR2_X1    g680(.A1(new_n678_), .A2(G162gat), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n881_), .B1(new_n866_), .B2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT123), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n881_), .B(KEYINPUT123), .C1(new_n866_), .C2(new_n882_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(G1347gat));
  INV_X1    g686(.A(KEYINPUT62), .ZN(new_n888_));
  INV_X1    g687(.A(new_n673_), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n427_), .A2(new_n635_), .A3(new_n424_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n835_), .A2(new_n889_), .A3(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n474_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n888_), .B1(new_n893_), .B2(G169gat), .ZN(new_n894_));
  AOI211_X1 g693(.A(KEYINPUT62), .B(new_n203_), .C1(new_n892_), .C2(new_n474_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n474_), .A2(new_n254_), .ZN(new_n896_));
  XOR2_X1   g695(.A(new_n896_), .B(KEYINPUT124), .Z(new_n897_));
  OAI22_X1  g696(.A1(new_n894_), .A2(new_n895_), .B1(new_n891_), .B2(new_n897_), .ZN(G1348gat));
  AOI21_X1  g697(.A(G176gat), .B1(new_n892_), .B2(new_n644_), .ZN(new_n899_));
  AND3_X1   g698(.A1(new_n890_), .A2(G176gat), .A3(new_n644_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n777_), .A2(new_n780_), .ZN(new_n901_));
  AOI22_X1  g700(.A1(new_n775_), .A2(new_n901_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n902_));
  OAI21_X1  g701(.A(KEYINPUT125), .B1(new_n902_), .B2(new_n418_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT125), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n843_), .A2(new_n905_), .A3(new_n331_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n906_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n900_), .B1(new_n904_), .B2(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT126), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  OAI211_X1 g709(.A(KEYINPUT126), .B(new_n900_), .C1(new_n904_), .C2(new_n907_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n899_), .B1(new_n910_), .B2(new_n911_), .ZN(G1349gat));
  NAND2_X1  g711(.A1(new_n890_), .A2(new_n626_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n913_), .A2(new_n224_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n835_), .A2(new_n889_), .A3(new_n914_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n913_), .B1(new_n903_), .B2(new_n906_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n915_), .B1(new_n916_), .B2(G183gat), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT127), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(new_n919_));
  OAI211_X1 g718(.A(new_n915_), .B(KEYINPUT127), .C1(new_n916_), .C2(G183gat), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n920_), .ZN(G1350gat));
  OAI21_X1  g720(.A(G190gat), .B1(new_n891_), .B2(new_n684_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n595_), .A2(new_n606_), .A3(new_n225_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n922_), .B1(new_n891_), .B2(new_n923_), .ZN(G1351gat));
  NAND3_X1  g723(.A1(new_n423_), .A2(new_n418_), .A3(new_n381_), .ZN(new_n925_));
  NOR3_X1   g724(.A1(new_n902_), .A2(new_n667_), .A3(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(new_n474_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g727(.A1(new_n926_), .A2(new_n644_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g729(.A1(new_n926_), .A2(new_n626_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n932_));
  AND2_X1   g731(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n933_));
  NOR3_X1   g732(.A1(new_n931_), .A2(new_n932_), .A3(new_n933_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n934_), .B1(new_n931_), .B2(new_n932_), .ZN(G1354gat));
  NAND2_X1  g734(.A1(new_n926_), .A2(new_n683_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n936_), .A2(G218gat), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n678_), .A2(G218gat), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n926_), .A2(new_n938_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n937_), .A2(new_n939_), .ZN(G1355gat));
endmodule


