//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 1 0 1 0 1 1 1 1 1 0 1 0 1 0 0 1 0 1 1 1 1 1 0 1 0 0 0 0 0 1 1 0 0 1 0 1 0 0 1 1 1 0 1 1 0 0 0 1 0 0 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n628_, new_n629_, new_n630_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n673_, new_n674_, new_n675_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n686_, new_n687_, new_n688_, new_n689_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n714_, new_n715_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n856_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n893_, new_n894_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n906_, new_n907_;
  INV_X1    g000(.A(KEYINPUT96), .ZN(new_n202_));
  XOR2_X1   g001(.A(G8gat), .B(G36gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(G92gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT18), .B(G64gat), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  INV_X1    g005(.A(G169gat), .ZN(new_n207_));
  INV_X1    g006(.A(G176gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  XOR2_X1   g008(.A(KEYINPUT22), .B(G169gat), .Z(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n209_), .B1(new_n211_), .B2(new_n208_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT86), .B(KEYINPUT23), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT87), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G183gat), .A2(G190gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n217_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT23), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n216_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n221_), .B1(new_n219_), .B2(new_n214_), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n218_), .B(new_n222_), .C1(G183gat), .C2(G190gat), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT94), .ZN(new_n224_));
  OR2_X1    g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n223_), .A2(new_n224_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n213_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  XOR2_X1   g026(.A(G197gat), .B(G204gat), .Z(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT21), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G211gat), .B(G218gat), .ZN(new_n230_));
  OR2_X1    g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n228_), .A2(KEYINPUT21), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n229_), .A2(new_n230_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n231_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(G183gat), .ZN(new_n235_));
  OR2_X1    g034(.A1(new_n235_), .A2(KEYINPUT25), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(KEYINPUT25), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(KEYINPUT26), .B(G190gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT24), .B1(new_n207_), .B2(new_n208_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(G169gat), .A2(G176gat), .ZN(new_n242_));
  MUX2_X1   g041(.A(new_n241_), .B(KEYINPUT24), .S(new_n242_), .Z(new_n243_));
  NAND2_X1  g042(.A1(new_n240_), .A2(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n219_), .A2(new_n220_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n245_), .B1(new_n219_), .B2(new_n214_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  NOR3_X1   g046(.A1(new_n227_), .A2(new_n234_), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n249_), .A2(KEYINPUT95), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(G183gat), .A2(G190gat), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n212_), .B1(new_n246_), .B2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n243_), .A2(new_n218_), .A3(new_n222_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n236_), .B(KEYINPUT83), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT26), .ZN(new_n256_));
  OR3_X1    g055(.A1(new_n256_), .A2(KEYINPUT84), .A3(G190gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(G190gat), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT85), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT84), .B1(new_n256_), .B2(G190gat), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n257_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n237_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n263_));
  NOR3_X1   g062(.A1(new_n255_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n253_), .B1(new_n254_), .B2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(new_n234_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G226gat), .A2(G233gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT19), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT20), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n266_), .A2(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n271_), .B1(new_n249_), .B2(KEYINPUT95), .ZN(new_n272_));
  AND2_X1   g071(.A1(new_n251_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n268_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n234_), .B1(new_n227_), .B2(new_n247_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n265_), .A2(new_n234_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n276_), .A2(new_n269_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n274_), .B1(new_n275_), .B2(new_n277_), .ZN(new_n278_));
  OAI211_X1 g077(.A(new_n202_), .B(new_n206_), .C1(new_n273_), .C2(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n278_), .B1(new_n251_), .B2(new_n272_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n206_), .ZN(new_n281_));
  OAI21_X1  g080(.A(KEYINPUT96), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n280_), .A2(new_n281_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n279_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT27), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n269_), .B1(new_n265_), .B2(new_n234_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n274_), .B1(new_n249_), .B2(new_n286_), .ZN(new_n287_));
  AND3_X1   g086(.A1(new_n275_), .A2(new_n274_), .A3(new_n277_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n206_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  AND2_X1   g088(.A1(new_n289_), .A2(KEYINPUT27), .ZN(new_n290_));
  AOI22_X1  g089(.A1(new_n284_), .A2(new_n285_), .B1(new_n283_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT92), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G141gat), .A2(G148gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT2), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT89), .ZN(new_n295_));
  OR4_X1    g094(.A1(new_n295_), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n296_));
  OR2_X1    g095(.A1(G141gat), .A2(G148gat), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT3), .B1(new_n297_), .B2(new_n295_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n294_), .A2(new_n296_), .A3(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G155gat), .A2(G162gat), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT88), .B1(G155gat), .B2(G162gat), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NOR3_X1   g101(.A1(KEYINPUT88), .A2(G155gat), .A3(G162gat), .ZN(new_n303_));
  OAI211_X1 g102(.A(new_n299_), .B(new_n300_), .C1(new_n302_), .C2(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n302_), .A2(new_n303_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n300_), .B(KEYINPUT1), .ZN(new_n306_));
  OAI211_X1 g105(.A(new_n297_), .B(new_n293_), .C1(new_n305_), .C2(new_n306_), .ZN(new_n307_));
  AND2_X1   g106(.A1(new_n304_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT29), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n292_), .B(new_n234_), .C1(new_n308_), .C2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(G233gat), .ZN(new_n311_));
  OR2_X1    g110(.A1(KEYINPUT91), .A2(G228gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(KEYINPUT91), .A2(G228gat), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n311_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n310_), .B(new_n314_), .ZN(new_n315_));
  XOR2_X1   g114(.A(G78gat), .B(G106gat), .Z(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n315_), .B(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(KEYINPUT93), .B1(new_n315_), .B2(new_n317_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n308_), .A2(new_n309_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT90), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G22gat), .B(G50gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT28), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n321_), .B(new_n323_), .ZN(new_n324_));
  OR3_X1    g123(.A1(new_n318_), .A2(new_n319_), .A3(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n318_), .B1(new_n324_), .B2(new_n319_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(KEYINPUT100), .B1(new_n291_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n291_), .A2(KEYINPUT100), .A3(new_n327_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G127gat), .B(G134gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G113gat), .B(G120gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  XOR2_X1   g133(.A(new_n308_), .B(new_n334_), .Z(new_n335_));
  NAND2_X1  g134(.A1(G225gat), .A2(G233gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT97), .ZN(new_n337_));
  OR2_X1    g136(.A1(new_n335_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n335_), .A2(KEYINPUT4), .ZN(new_n339_));
  OR3_X1    g138(.A1(new_n308_), .A2(KEYINPUT4), .A3(new_n334_), .ZN(new_n340_));
  AND2_X1   g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n337_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n338_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT98), .B(KEYINPUT0), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G1gat), .B(G29gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G57gat), .B(G85gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  OR2_X1    g147(.A1(new_n343_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n343_), .A2(new_n348_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G71gat), .B(G99gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(G43gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n265_), .B(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G227gat), .A2(G233gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n334_), .B(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT30), .B(G15gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT31), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n356_), .B(new_n358_), .ZN(new_n359_));
  OR2_X1    g158(.A1(new_n354_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n354_), .A2(new_n359_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n351_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n281_), .A2(KEYINPUT32), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n280_), .A2(new_n364_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n287_), .A2(new_n288_), .ZN(new_n366_));
  OAI211_X1 g165(.A(new_n351_), .B(new_n365_), .C1(new_n364_), .C2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n341_), .A2(new_n342_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n348_), .B1(new_n335_), .B2(new_n337_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(KEYINPUT99), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n350_), .A2(KEYINPUT33), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT33), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n343_), .A2(new_n373_), .A3(new_n348_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n372_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n371_), .A2(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n367_), .B1(new_n376_), .B2(new_n284_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(new_n327_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n327_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n351_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n291_), .A2(new_n379_), .A3(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n378_), .A2(new_n381_), .ZN(new_n382_));
  AOI22_X1  g181(.A1(new_n331_), .A2(new_n363_), .B1(new_n382_), .B2(new_n362_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT13), .ZN(new_n384_));
  XOR2_X1   g183(.A(G176gat), .B(G204gat), .Z(new_n385_));
  XNOR2_X1  g184(.A(G120gat), .B(G148gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT75), .B(KEYINPUT5), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G71gat), .B(G78gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G57gat), .B(G64gat), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n390_), .B1(KEYINPUT11), .B2(new_n391_), .ZN(new_n392_));
  XOR2_X1   g191(.A(G57gat), .B(G64gat), .Z(new_n393_));
  INV_X1    g192(.A(KEYINPUT11), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n392_), .A2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n391_), .A2(new_n390_), .A3(KEYINPUT11), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G85gat), .A2(G92gat), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(G85gat), .A2(G92gat), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT67), .ZN(new_n404_));
  NAND3_X1  g203(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n404_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G99gat), .A2(G106gat), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT6), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n411_), .A2(KEYINPUT67), .A3(new_n405_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n408_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT7), .ZN(new_n414_));
  INV_X1    g213(.A(G99gat), .ZN(new_n415_));
  INV_X1    g214(.A(G106gat), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n414_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  AOI211_X1 g219(.A(KEYINPUT8), .B(new_n403_), .C1(new_n413_), .C2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n411_), .A2(new_n405_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n423_), .B1(new_n419_), .B2(KEYINPUT69), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT69), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n417_), .A2(new_n425_), .A3(new_n418_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n403_), .B1(new_n424_), .B2(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT8), .B1(new_n427_), .B2(KEYINPUT70), .ZN(new_n428_));
  INV_X1    g227(.A(new_n418_), .ZN(new_n429_));
  NOR3_X1   g228(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT69), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n423_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n431_), .A2(new_n432_), .A3(new_n426_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n433_), .A2(KEYINPUT70), .A3(new_n402_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n422_), .B1(new_n428_), .B2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n415_), .A2(KEYINPUT10), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT10), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(G99gat), .ZN(new_n439_));
  AND3_X1   g238(.A1(new_n437_), .A2(new_n439_), .A3(KEYINPUT65), .ZN(new_n440_));
  AOI21_X1  g239(.A(KEYINPUT65), .B1(new_n437_), .B2(new_n439_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n416_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT66), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT9), .ZN(new_n444_));
  NOR3_X1   g243(.A1(new_n399_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT9), .B1(new_n400_), .B2(new_n401_), .ZN(new_n446_));
  AOI21_X1  g245(.A(KEYINPUT66), .B1(new_n399_), .B2(new_n444_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n445_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n442_), .A2(new_n413_), .A3(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT68), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT68), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n442_), .A2(new_n451_), .A3(new_n448_), .A4(new_n413_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n398_), .B1(new_n436_), .B2(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(KEYINPUT74), .B1(new_n455_), .B2(KEYINPUT12), .ZN(new_n456_));
  INV_X1    g255(.A(new_n398_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT8), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n433_), .A2(new_n402_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT70), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n458_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n421_), .B1(new_n461_), .B2(new_n434_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n457_), .B1(new_n462_), .B2(new_n453_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT74), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT12), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n463_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT73), .ZN(new_n467_));
  AOI211_X1 g266(.A(new_n467_), .B(new_n421_), .C1(new_n461_), .C2(new_n434_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n459_), .A2(new_n460_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n469_), .A2(KEYINPUT8), .A3(new_n434_), .ZN(new_n470_));
  AOI21_X1  g269(.A(KEYINPUT73), .B1(new_n470_), .B2(new_n422_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n454_), .B1(new_n468_), .B2(new_n471_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n398_), .A2(new_n465_), .ZN(new_n473_));
  AOI22_X1  g272(.A1(new_n456_), .A2(new_n466_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G230gat), .A2(G233gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT64), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n453_), .B1(new_n470_), .B2(new_n422_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n476_), .B1(new_n477_), .B2(new_n398_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n436_), .A2(new_n454_), .A3(new_n398_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT71), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n477_), .A2(KEYINPUT71), .A3(new_n398_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n455_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n476_), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT72), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(KEYINPUT71), .B1(new_n477_), .B2(new_n398_), .ZN(new_n486_));
  NOR4_X1   g285(.A1(new_n462_), .A2(new_n453_), .A3(new_n480_), .A4(new_n457_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n463_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT72), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n488_), .A2(new_n489_), .A3(new_n476_), .ZN(new_n490_));
  AOI221_X4 g289(.A(new_n389_), .B1(new_n474_), .B2(new_n478_), .C1(new_n485_), .C2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n389_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n485_), .A2(new_n490_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n472_), .A2(new_n473_), .ZN(new_n494_));
  NOR3_X1   g293(.A1(new_n455_), .A2(KEYINPUT74), .A3(KEYINPUT12), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n464_), .B1(new_n463_), .B2(new_n465_), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n494_), .B(new_n478_), .C1(new_n495_), .C2(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n492_), .B1(new_n493_), .B2(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n384_), .B1(new_n491_), .B2(new_n498_), .ZN(new_n499_));
  NOR3_X1   g298(.A1(new_n483_), .A2(KEYINPUT72), .A3(new_n484_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n489_), .B1(new_n488_), .B2(new_n476_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n497_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(new_n389_), .ZN(new_n503_));
  AOI22_X1  g302(.A1(new_n485_), .A2(new_n490_), .B1(new_n474_), .B2(new_n478_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(new_n492_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n503_), .A2(new_n505_), .A3(KEYINPUT13), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n499_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G229gat), .A2(G233gat), .ZN(new_n508_));
  XOR2_X1   g307(.A(G43gat), .B(G50gat), .Z(new_n509_));
  XNOR2_X1  g308(.A(G29gat), .B(G36gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  XOR2_X1   g313(.A(G1gat), .B(G8gat), .Z(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT81), .ZN(new_n516_));
  INV_X1    g315(.A(G15gat), .ZN(new_n517_));
  INV_X1    g316(.A(G22gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G15gat), .A2(G22gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G1gat), .A2(G8gat), .ZN(new_n521_));
  AOI22_X1  g320(.A1(new_n519_), .A2(new_n520_), .B1(KEYINPUT14), .B2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n516_), .B(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n514_), .A2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n513_), .B(KEYINPUT15), .ZN(new_n525_));
  OAI211_X1 g324(.A(new_n508_), .B(new_n524_), .C1(new_n525_), .C2(new_n523_), .ZN(new_n526_));
  XOR2_X1   g325(.A(new_n513_), .B(new_n523_), .Z(new_n527_));
  INV_X1    g326(.A(new_n508_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G113gat), .B(G141gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G169gat), .B(G197gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n526_), .A2(new_n529_), .A3(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n533_), .B1(new_n526_), .B2(new_n529_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n507_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G231gat), .A2(G233gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n398_), .B(new_n540_), .ZN(new_n541_));
  XOR2_X1   g340(.A(new_n541_), .B(new_n523_), .Z(new_n542_));
  XNOR2_X1  g341(.A(G127gat), .B(G155gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(G211gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(KEYINPUT16), .B(G183gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT17), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n542_), .A2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n541_), .B(new_n523_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n546_), .A2(KEYINPUT17), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  AND2_X1   g350(.A1(new_n548_), .A2(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT82), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT80), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G190gat), .B(G218gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G134gat), .B(G162gat), .ZN(new_n556_));
  XOR2_X1   g355(.A(new_n555_), .B(new_n556_), .Z(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT36), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n436_), .A2(new_n467_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n462_), .A2(KEYINPUT73), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n453_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G232gat), .A2(G233gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT34), .ZN(new_n563_));
  OAI22_X1  g362(.A1(new_n561_), .A2(new_n525_), .B1(KEYINPUT35), .B2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT78), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n565_), .B1(new_n477_), .B2(new_n514_), .ZN(new_n566_));
  NOR4_X1   g365(.A1(new_n462_), .A2(new_n513_), .A3(new_n453_), .A4(KEYINPUT78), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n563_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT35), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NOR3_X1   g370(.A1(new_n564_), .A2(new_n568_), .A3(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n571_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n525_), .ZN(new_n574_));
  AOI22_X1  g373(.A1(new_n574_), .A2(new_n472_), .B1(new_n570_), .B2(new_n569_), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n566_), .A2(new_n567_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n573_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n558_), .B1(new_n572_), .B2(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n571_), .B1(new_n564_), .B2(new_n568_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT36), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n575_), .A2(new_n576_), .A3(new_n573_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n579_), .A2(new_n580_), .A3(new_n581_), .A4(new_n557_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT37), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n578_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n558_), .B(KEYINPUT79), .Z(new_n585_));
  OAI21_X1  g384(.A(new_n585_), .B1(new_n572_), .B2(new_n577_), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n586_), .A2(new_n582_), .ZN(new_n587_));
  OAI211_X1 g386(.A(new_n554_), .B(new_n584_), .C1(new_n587_), .C2(new_n583_), .ZN(new_n588_));
  AND3_X1   g387(.A1(new_n578_), .A2(new_n583_), .A3(new_n582_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n583_), .B1(new_n586_), .B2(new_n582_), .ZN(new_n590_));
  OAI21_X1  g389(.A(KEYINPUT80), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n588_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NOR4_X1   g392(.A1(new_n383_), .A2(new_n539_), .A3(new_n553_), .A4(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(G1gat), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n594_), .A2(new_n595_), .A3(new_n351_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT38), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n382_), .A2(new_n362_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n330_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n363_), .B1(new_n600_), .B2(new_n328_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n539_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n578_), .A2(new_n582_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n605_), .A2(new_n553_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n602_), .A2(new_n603_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(G1gat), .B1(new_n608_), .B2(new_n380_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n596_), .A2(new_n597_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n598_), .A2(new_n609_), .A3(new_n610_), .ZN(G1324gat));
  INV_X1    g410(.A(G8gat), .ZN(new_n612_));
  INV_X1    g411(.A(new_n291_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n612_), .B1(new_n607_), .B2(new_n613_), .ZN(new_n614_));
  XOR2_X1   g413(.A(KEYINPUT101), .B(KEYINPUT39), .Z(new_n615_));
  OR2_X1    g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n594_), .A2(new_n612_), .A3(new_n613_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n614_), .A2(new_n615_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n616_), .A2(new_n617_), .A3(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(G1325gat));
  OAI21_X1  g420(.A(G15gat), .B1(new_n608_), .B2(new_n362_), .ZN(new_n622_));
  OR2_X1    g421(.A1(new_n622_), .A2(KEYINPUT41), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(KEYINPUT41), .ZN(new_n624_));
  INV_X1    g423(.A(new_n362_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n594_), .A2(new_n517_), .A3(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n623_), .A2(new_n624_), .A3(new_n626_), .ZN(G1326gat));
  AOI21_X1  g426(.A(new_n518_), .B1(new_n607_), .B2(new_n379_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n628_), .B(KEYINPUT42), .Z(new_n629_));
  NAND3_X1  g428(.A1(new_n594_), .A2(new_n518_), .A3(new_n379_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(G1327gat));
  NOR2_X1   g430(.A1(new_n383_), .A2(new_n539_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n553_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n633_), .A2(new_n604_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(G29gat), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n636_), .A2(new_n637_), .A3(new_n351_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n539_), .A2(new_n633_), .ZN(new_n639_));
  NOR3_X1   g438(.A1(new_n383_), .A2(KEYINPUT43), .A3(new_n592_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT43), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n641_), .B1(new_n602_), .B2(new_n593_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n639_), .B1(new_n640_), .B2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT44), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  OAI211_X1 g445(.A(KEYINPUT44), .B(new_n639_), .C1(new_n640_), .C2(new_n642_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n646_), .A2(new_n648_), .A3(new_n380_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n638_), .B1(new_n649_), .B2(new_n637_), .ZN(G1328gat));
  NOR2_X1   g449(.A1(new_n291_), .A2(G36gat), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n602_), .A2(new_n603_), .A3(new_n634_), .A4(new_n651_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT45), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT103), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT46), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n653_), .A2(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n645_), .A2(new_n613_), .A3(new_n647_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n657_), .B1(new_n658_), .B2(G36gat), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n654_), .A2(new_n655_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n659_), .A2(new_n661_), .ZN(new_n662_));
  AOI211_X1 g461(.A(new_n660_), .B(new_n657_), .C1(new_n658_), .C2(G36gat), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1329gat));
  NOR3_X1   g463(.A1(new_n635_), .A2(G43gat), .A3(new_n362_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n645_), .A2(new_n625_), .A3(new_n647_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n665_), .B1(new_n666_), .B2(G43gat), .ZN(new_n667_));
  XNOR2_X1  g466(.A(KEYINPUT104), .B(KEYINPUT47), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n668_), .ZN(new_n670_));
  AOI211_X1 g469(.A(new_n665_), .B(new_n670_), .C1(new_n666_), .C2(G43gat), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n669_), .A2(new_n671_), .ZN(G1330gat));
  INV_X1    g471(.A(G50gat), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n636_), .A2(new_n673_), .A3(new_n379_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n646_), .A2(new_n648_), .A3(new_n327_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n674_), .B1(new_n675_), .B2(new_n673_), .ZN(G1331gat));
  NOR2_X1   g475(.A1(new_n507_), .A2(new_n538_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n602_), .A2(new_n677_), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n678_), .A2(new_n633_), .A3(new_n592_), .ZN(new_n679_));
  INV_X1    g478(.A(G57gat), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n679_), .A2(new_n680_), .A3(new_n351_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n678_), .A2(new_n606_), .ZN(new_n682_));
  OAI21_X1  g481(.A(G57gat), .B1(new_n682_), .B2(new_n380_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n681_), .A2(new_n683_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT105), .ZN(G1332gat));
  OAI21_X1  g484(.A(G64gat), .B1(new_n682_), .B2(new_n291_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT48), .ZN(new_n687_));
  INV_X1    g486(.A(G64gat), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n679_), .A2(new_n688_), .A3(new_n613_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n689_), .ZN(G1333gat));
  OAI21_X1  g489(.A(G71gat), .B1(new_n682_), .B2(new_n362_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT49), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n362_), .A2(G71gat), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT106), .Z(new_n694_));
  NAND2_X1  g493(.A1(new_n679_), .A2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n692_), .A2(new_n695_), .ZN(G1334gat));
  INV_X1    g495(.A(G78gat), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n679_), .A2(new_n697_), .A3(new_n379_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n682_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n697_), .B1(new_n699_), .B2(new_n379_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n700_), .A2(new_n701_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n698_), .B1(new_n702_), .B2(new_n703_), .ZN(G1335gat));
  NAND2_X1  g503(.A1(new_n678_), .A2(new_n634_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(G85gat), .B1(new_n706_), .B2(new_n351_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n677_), .A2(new_n553_), .ZN(new_n708_));
  XOR2_X1   g507(.A(new_n708_), .B(KEYINPUT108), .Z(new_n709_));
  OAI21_X1  g508(.A(new_n709_), .B1(new_n640_), .B2(new_n642_), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT109), .Z(new_n711_));
  AND2_X1   g510(.A1(new_n351_), .A2(G85gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n707_), .B1(new_n711_), .B2(new_n712_), .ZN(G1336gat));
  AOI21_X1  g512(.A(G92gat), .B1(new_n706_), .B2(new_n613_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n613_), .A2(G92gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n711_), .B2(new_n715_), .ZN(G1337gat));
  OAI211_X1 g515(.A(new_n706_), .B(new_n625_), .C1(new_n441_), .C2(new_n440_), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n625_), .B(new_n709_), .C1(new_n640_), .C2(new_n642_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT110), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n718_), .A2(new_n719_), .A3(G99gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(new_n718_), .B2(G99gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n717_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g522(.A1(new_n706_), .A2(new_n416_), .A3(new_n379_), .ZN(new_n724_));
  OAI211_X1 g523(.A(new_n379_), .B(new_n709_), .C1(new_n640_), .C2(new_n642_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT52), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n725_), .A2(new_n726_), .A3(G106gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n725_), .B2(G106gat), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n724_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n729_), .B(new_n731_), .ZN(G1339gat));
  INV_X1    g531(.A(KEYINPUT54), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n553_), .A2(new_n538_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n499_), .A2(new_n506_), .A3(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT112), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n499_), .A2(new_n506_), .A3(new_n734_), .A4(KEYINPUT112), .ZN(new_n738_));
  AOI22_X1  g537(.A1(new_n737_), .A2(new_n738_), .B1(new_n591_), .B2(new_n588_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n733_), .B1(new_n739_), .B2(KEYINPUT113), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n737_), .A2(new_n738_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT114), .ZN(new_n742_));
  AND4_X1   g541(.A1(KEYINPUT113), .A2(new_n741_), .A3(new_n742_), .A4(new_n592_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n739_), .B2(KEYINPUT113), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n740_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n741_), .A2(KEYINPUT113), .A3(new_n592_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(KEYINPUT114), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n741_), .A2(new_n592_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT113), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n739_), .A2(KEYINPUT113), .A3(new_n742_), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n747_), .A2(new_n750_), .A3(new_n733_), .A4(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n745_), .A2(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n533_), .B1(new_n527_), .B2(new_n508_), .ZN(new_n754_));
  OR2_X1    g553(.A1(new_n754_), .A2(KEYINPUT116), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(KEYINPUT116), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n528_), .B(new_n524_), .C1(new_n525_), .C2(new_n523_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n755_), .A2(new_n756_), .A3(new_n757_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n758_), .A2(new_n534_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n759_), .B1(new_n491_), .B2(new_n498_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n537_), .B1(new_n504_), .B2(new_n492_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n481_), .A2(new_n482_), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n494_), .B(new_n762_), .C1(new_n495_), .C2(new_n496_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(new_n476_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT55), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n497_), .A2(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n474_), .A2(KEYINPUT55), .A3(new_n478_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n764_), .A2(new_n766_), .A3(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(KEYINPUT115), .B1(new_n768_), .B2(new_n389_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n761_), .B1(new_n769_), .B2(KEYINPUT56), .ZN(new_n770_));
  AOI22_X1  g569(.A1(new_n765_), .A2(new_n497_), .B1(new_n763_), .B2(new_n476_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n492_), .B1(new_n771_), .B2(new_n767_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT56), .ZN(new_n773_));
  NOR3_X1   g572(.A1(new_n772_), .A2(KEYINPUT115), .A3(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n760_), .B1(new_n770_), .B2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n775_), .A2(KEYINPUT57), .A3(new_n604_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(KEYINPUT117), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n604_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT57), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n759_), .A2(new_n505_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT118), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n768_), .A2(new_n782_), .A3(KEYINPUT56), .A4(new_n389_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n783_), .B1(new_n772_), .B2(KEYINPUT56), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n782_), .B1(new_n772_), .B2(KEYINPUT56), .ZN(new_n785_));
  OAI211_X1 g584(.A(KEYINPUT58), .B(new_n781_), .C1(new_n784_), .C2(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n781_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT58), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n592_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  AOI22_X1  g588(.A1(new_n777_), .A2(new_n780_), .B1(new_n786_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT117), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n773_), .B1(new_n772_), .B2(KEYINPUT115), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n769_), .A2(KEYINPUT56), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n792_), .A2(new_n793_), .A3(new_n761_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n605_), .B1(new_n794_), .B2(new_n760_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n791_), .B1(new_n795_), .B2(KEYINPUT57), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n795_), .A2(KEYINPUT57), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n633_), .B1(new_n790_), .B2(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(KEYINPUT119), .B1(new_n753_), .B2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n787_), .A2(new_n788_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n801_), .A2(new_n593_), .A3(new_n786_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n802_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n777_), .A2(new_n780_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n553_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT119), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n805_), .A2(new_n806_), .A3(new_n752_), .A4(new_n745_), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n800_), .A2(new_n807_), .ZN(new_n808_));
  AOI211_X1 g607(.A(new_n380_), .B(new_n362_), .C1(new_n329_), .C2(new_n330_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n808_), .A2(new_n538_), .A3(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(G113gat), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n802_), .A2(new_n780_), .A3(new_n776_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n553_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n745_), .A2(new_n752_), .A3(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT59), .ZN(new_n815_));
  AND2_X1   g614(.A1(new_n809_), .A2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n814_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n800_), .A2(new_n807_), .A3(new_n809_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n818_), .B1(new_n819_), .B2(KEYINPUT59), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n537_), .A2(new_n811_), .ZN(new_n821_));
  AOI22_X1  g620(.A1(new_n810_), .A2(new_n811_), .B1(new_n820_), .B2(new_n821_), .ZN(G1340gat));
  INV_X1    g621(.A(new_n507_), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n820_), .A2(new_n823_), .ZN(new_n824_));
  XOR2_X1   g623(.A(KEYINPUT120), .B(G120gat), .Z(new_n825_));
  OAI21_X1  g624(.A(new_n825_), .B1(new_n507_), .B2(KEYINPUT60), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(KEYINPUT60), .B2(new_n825_), .ZN(new_n827_));
  OAI22_X1  g626(.A1(new_n824_), .A2(new_n825_), .B1(new_n819_), .B2(new_n827_), .ZN(G1341gat));
  INV_X1    g627(.A(KEYINPUT122), .ZN(new_n829_));
  NOR2_X1   g628(.A1(KEYINPUT121), .A2(G127gat), .ZN(new_n830_));
  AND2_X1   g629(.A1(KEYINPUT121), .A2(G127gat), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n830_), .B1(new_n633_), .B2(new_n831_), .ZN(new_n832_));
  AOI211_X1 g631(.A(new_n818_), .B(new_n832_), .C1(new_n819_), .C2(KEYINPUT59), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n800_), .A2(new_n807_), .A3(new_n633_), .A4(new_n809_), .ZN(new_n834_));
  INV_X1    g633(.A(G127gat), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n829_), .B1(new_n833_), .B2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n819_), .A2(KEYINPUT59), .ZN(new_n839_));
  INV_X1    g638(.A(new_n832_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n839_), .A2(new_n817_), .A3(new_n840_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n841_), .A2(KEYINPUT122), .A3(new_n836_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n838_), .A2(new_n842_), .ZN(G1342gat));
  INV_X1    g642(.A(G134gat), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n592_), .A2(new_n844_), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n820_), .A2(new_n845_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n800_), .A2(new_n807_), .A3(new_n605_), .A4(new_n809_), .ZN(new_n847_));
  AND3_X1   g646(.A1(new_n847_), .A2(KEYINPUT123), .A3(new_n844_), .ZN(new_n848_));
  AOI21_X1  g647(.A(KEYINPUT123), .B1(new_n847_), .B2(new_n844_), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n846_), .A2(new_n848_), .A3(new_n849_), .ZN(G1343gat));
  NOR2_X1   g649(.A1(new_n327_), .A2(new_n625_), .ZN(new_n851_));
  AND3_X1   g650(.A1(new_n800_), .A2(new_n807_), .A3(new_n851_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n613_), .A2(new_n380_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n852_), .A2(new_n538_), .A3(new_n853_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g654(.A1(new_n852_), .A2(new_n823_), .A3(new_n853_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g656(.A1(new_n852_), .A2(new_n633_), .A3(new_n853_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(KEYINPUT61), .B(G155gat), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n858_), .B(new_n859_), .ZN(G1346gat));
  AND4_X1   g659(.A1(G162gat), .A2(new_n852_), .A3(new_n593_), .A4(new_n853_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n852_), .A2(new_n605_), .A3(new_n853_), .ZN(new_n862_));
  INV_X1    g661(.A(G162gat), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n861_), .B1(new_n862_), .B2(new_n863_), .ZN(G1347gat));
  XOR2_X1   g663(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n865_));
  NAND2_X1  g664(.A1(new_n613_), .A2(new_n363_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n814_), .A2(new_n538_), .A3(new_n327_), .A4(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n865_), .B1(new_n869_), .B2(new_n207_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT125), .ZN(new_n871_));
  INV_X1    g670(.A(new_n865_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n868_), .A2(G169gat), .A3(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n870_), .B1(new_n871_), .B2(new_n873_), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n873_), .A2(new_n871_), .ZN(new_n875_));
  OAI22_X1  g674(.A1(new_n874_), .A2(new_n875_), .B1(new_n210_), .B2(new_n868_), .ZN(G1348gat));
  AND2_X1   g675(.A1(new_n814_), .A2(new_n327_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(new_n867_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n208_), .B1(new_n878_), .B2(new_n507_), .ZN(new_n879_));
  NOR3_X1   g678(.A1(new_n866_), .A2(new_n208_), .A3(new_n507_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n808_), .A2(new_n327_), .A3(new_n880_), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n879_), .A2(new_n881_), .ZN(G1349gat));
  NAND4_X1  g681(.A1(new_n808_), .A2(new_n327_), .A3(new_n633_), .A4(new_n867_), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n866_), .A2(new_n238_), .A3(new_n553_), .ZN(new_n884_));
  AOI22_X1  g683(.A1(new_n883_), .A2(new_n235_), .B1(new_n877_), .B2(new_n884_), .ZN(G1350gat));
  OAI21_X1  g684(.A(G190gat), .B1(new_n878_), .B2(new_n592_), .ZN(new_n886_));
  NAND4_X1  g685(.A1(new_n877_), .A2(new_n239_), .A3(new_n605_), .A4(new_n867_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(KEYINPUT126), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT126), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n886_), .A2(new_n890_), .A3(new_n887_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n891_), .ZN(G1351gat));
  NOR2_X1   g691(.A1(new_n291_), .A2(new_n351_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n852_), .A2(new_n538_), .A3(new_n893_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g694(.A1(new_n852_), .A2(new_n823_), .A3(new_n893_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g696(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n852_), .A2(new_n893_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n899_), .B2(new_n553_), .ZN(new_n900_));
  XOR2_X1   g699(.A(KEYINPUT63), .B(G211gat), .Z(new_n901_));
  NAND4_X1  g700(.A1(new_n852_), .A2(new_n633_), .A3(new_n893_), .A4(new_n901_), .ZN(new_n902_));
  AND2_X1   g701(.A1(new_n900_), .A2(new_n902_), .ZN(G1354gat));
  XOR2_X1   g702(.A(KEYINPUT127), .B(G218gat), .Z(new_n904_));
  OR2_X1    g703(.A1(new_n592_), .A2(new_n904_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n899_), .A2(new_n905_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n852_), .A2(new_n605_), .A3(new_n893_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n906_), .B1(new_n907_), .B2(new_n904_), .ZN(G1355gat));
endmodule


