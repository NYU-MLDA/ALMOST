//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 1 1 0 0 0 1 1 0 1 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 1 0 1 0 1 0 1 0 1 1 1 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n807_, new_n808_, new_n809_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n898_, new_n900_, new_n901_,
    new_n903_, new_n904_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n917_,
    new_n918_, new_n920_, new_n921_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n932_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_;
  INV_X1    g000(.A(KEYINPUT13), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT8), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G99gat), .A2(G106gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT7), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT6), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT6), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n208_), .A2(G99gat), .A3(G106gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n207_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n205_), .A2(new_n210_), .ZN(new_n211_));
  XOR2_X1   g010(.A(G85gat), .B(G92gat), .Z(new_n212_));
  AOI21_X1  g011(.A(new_n203_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n210_), .B(KEYINPUT64), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(new_n205_), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n212_), .A2(new_n203_), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n213_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  XOR2_X1   g016(.A(KEYINPUT10), .B(G99gat), .Z(new_n218_));
  INV_X1    g017(.A(G106gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT9), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(G85gat), .A3(G92gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n212_), .A2(KEYINPUT9), .ZN(new_n223_));
  AND4_X1   g022(.A1(new_n214_), .A2(new_n220_), .A3(new_n222_), .A4(new_n223_), .ZN(new_n224_));
  OR3_X1    g023(.A1(new_n217_), .A2(KEYINPUT65), .A3(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT65), .B1(new_n217_), .B2(new_n224_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G57gat), .B(G64gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT11), .ZN(new_n228_));
  XOR2_X1   g027(.A(G71gat), .B(G78gat), .Z(new_n229_));
  OR2_X1    g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n228_), .A2(new_n229_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n227_), .A2(KEYINPUT11), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n230_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(new_n233_), .B(KEYINPUT66), .Z(new_n234_));
  NAND3_X1  g033(.A1(new_n225_), .A2(new_n226_), .A3(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n217_), .A2(new_n224_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT12), .ZN(new_n237_));
  OR3_X1    g036(.A1(new_n236_), .A2(new_n237_), .A3(new_n233_), .ZN(new_n238_));
  AND2_X1   g037(.A1(new_n235_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G230gat), .A2(G233gat), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n234_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n239_), .B(new_n240_), .C1(KEYINPUT12), .C2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n243_));
  INV_X1    g042(.A(new_n240_), .ZN(new_n244_));
  AND3_X1   g043(.A1(new_n225_), .A2(new_n226_), .A3(new_n234_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n244_), .B1(new_n245_), .B2(new_n241_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G120gat), .B(G148gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT5), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G176gat), .B(G204gat), .ZN(new_n249_));
  XOR2_X1   g048(.A(new_n248_), .B(new_n249_), .Z(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n242_), .A2(new_n243_), .A3(new_n246_), .A4(new_n251_), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n235_), .B(new_n238_), .C1(new_n241_), .C2(KEYINPUT12), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n246_), .B(new_n251_), .C1(new_n253_), .C2(new_n244_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT67), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n252_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n242_), .A2(new_n246_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(new_n250_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n256_), .A2(KEYINPUT68), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(KEYINPUT68), .B1(new_n256_), .B2(new_n258_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n202_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n256_), .A2(new_n258_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT68), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n265_), .A2(KEYINPUT13), .A3(new_n259_), .ZN(new_n266_));
  XOR2_X1   g065(.A(KEYINPUT73), .B(G1gat), .Z(new_n267_));
  XOR2_X1   g066(.A(KEYINPUT74), .B(G8gat), .Z(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(KEYINPUT14), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G15gat), .B(G22gat), .ZN(new_n271_));
  AND2_X1   g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G1gat), .B(G8gat), .ZN(new_n273_));
  OR2_X1    g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n270_), .A2(new_n271_), .A3(new_n273_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  XOR2_X1   g075(.A(G29gat), .B(G36gat), .Z(new_n277_));
  XOR2_X1   g076(.A(G43gat), .B(G50gat), .Z(new_n278_));
  XOR2_X1   g077(.A(new_n277_), .B(new_n278_), .Z(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n276_), .B(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G229gat), .A2(G233gat), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n281_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n276_), .ZN(new_n285_));
  XOR2_X1   g084(.A(new_n279_), .B(KEYINPUT15), .Z(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n276_), .A2(new_n280_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n287_), .A2(new_n288_), .A3(new_n282_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n284_), .A2(new_n289_), .ZN(new_n290_));
  XOR2_X1   g089(.A(G113gat), .B(G141gat), .Z(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT78), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT79), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G169gat), .B(G197gat), .ZN(new_n294_));
  XOR2_X1   g093(.A(new_n293_), .B(new_n294_), .Z(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n290_), .A2(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n284_), .A2(new_n289_), .A3(new_n295_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n262_), .A2(new_n266_), .A3(new_n299_), .ZN(new_n300_));
  XOR2_X1   g099(.A(G8gat), .B(G36gat), .Z(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G64gat), .B(G92gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT20), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G169gat), .A2(G176gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(KEYINPUT24), .ZN(new_n309_));
  OR2_X1    g108(.A1(new_n309_), .A2(KEYINPUT93), .ZN(new_n310_));
  INV_X1    g109(.A(G169gat), .ZN(new_n311_));
  INV_X1    g110(.A(G176gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n309_), .A2(KEYINPUT93), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n310_), .A2(new_n313_), .A3(new_n314_), .ZN(new_n315_));
  AND2_X1   g114(.A1(G183gat), .A2(G190gat), .ZN(new_n316_));
  AND2_X1   g115(.A1(KEYINPUT82), .A2(KEYINPUT23), .ZN(new_n317_));
  NOR2_X1   g116(.A1(KEYINPUT82), .A2(KEYINPUT23), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n316_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G183gat), .A2(G190gat), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT23), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n319_), .A2(new_n322_), .ZN(new_n323_));
  NOR3_X1   g122(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT26), .B(G190gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT25), .B(G183gat), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n324_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n315_), .A2(new_n323_), .A3(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n311_), .A2(KEYINPUT22), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT22), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(G169gat), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT94), .ZN(new_n332_));
  AND3_X1   g131(.A1(new_n329_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n332_), .B1(new_n329_), .B2(new_n331_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(new_n312_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n308_), .A2(KEYINPUT81), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT81), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n338_), .A2(G169gat), .A3(G176gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n336_), .A2(new_n341_), .ZN(new_n342_));
  OR2_X1    g141(.A1(KEYINPUT82), .A2(KEYINPUT23), .ZN(new_n343_));
  NAND2_X1  g142(.A1(KEYINPUT82), .A2(KEYINPUT23), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n316_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n320_), .A2(KEYINPUT23), .ZN(new_n346_));
  OAI21_X1  g145(.A(KEYINPUT83), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n320_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT83), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(G183gat), .ZN(new_n351_));
  INV_X1    g150(.A(G190gat), .ZN(new_n352_));
  AOI22_X1  g151(.A1(new_n347_), .A2(new_n350_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n328_), .B1(new_n342_), .B2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G211gat), .B(G218gat), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(G197gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(KEYINPUT92), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT92), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(G197gat), .ZN(new_n360_));
  INV_X1    g159(.A(G204gat), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n358_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT21), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n363_), .B1(G197gat), .B2(G204gat), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n356_), .B1(new_n362_), .B2(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n361_), .B1(new_n358_), .B2(new_n360_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(G197gat), .A2(G204gat), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n363_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n366_), .A2(new_n367_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n355_), .A2(new_n363_), .ZN(new_n370_));
  AOI22_X1  g169(.A1(new_n365_), .A2(new_n368_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n307_), .B1(new_n354_), .B2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G226gat), .A2(G233gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT19), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT84), .ZN(new_n377_));
  AOI21_X1  g176(.A(G176gat), .B1(new_n329_), .B2(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(KEYINPUT22), .B(G169gat), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n378_), .B1(new_n377_), .B2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n351_), .A2(new_n352_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n319_), .A2(new_n381_), .A3(new_n322_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n380_), .A2(new_n382_), .A3(new_n341_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n316_), .A2(new_n321_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n349_), .B1(new_n348_), .B2(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT82), .B(KEYINPUT23), .ZN(new_n386_));
  AOI21_X1  g185(.A(KEYINPUT83), .B1(new_n386_), .B2(new_n320_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n385_), .A2(new_n387_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n337_), .A2(new_n339_), .A3(new_n313_), .A4(KEYINPUT24), .ZN(new_n389_));
  INV_X1    g188(.A(new_n324_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT80), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n391_), .B1(new_n352_), .B2(KEYINPUT26), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n326_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT26), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(G190gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n352_), .A2(KEYINPUT26), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n391_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  OAI211_X1 g196(.A(new_n389_), .B(new_n390_), .C1(new_n393_), .C2(new_n397_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n383_), .B1(new_n388_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT85), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  OAI211_X1 g200(.A(KEYINPUT85), .B(new_n383_), .C1(new_n388_), .C2(new_n398_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n401_), .A2(new_n371_), .A3(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n373_), .A2(new_n376_), .A3(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n346_), .B1(new_n386_), .B2(new_n320_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n350_), .B1(new_n405_), .B2(new_n349_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n351_), .A2(KEYINPUT25), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT25), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(G183gat), .ZN(new_n409_));
  AND3_X1   g208(.A1(new_n392_), .A2(new_n407_), .A3(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n395_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n394_), .A2(G190gat), .ZN(new_n412_));
  OAI21_X1  g211(.A(KEYINPUT80), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n324_), .B1(new_n410_), .B2(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n406_), .A2(new_n414_), .A3(new_n389_), .ZN(new_n415_));
  AOI21_X1  g214(.A(KEYINPUT85), .B1(new_n415_), .B2(new_n383_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n402_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n372_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n340_), .B1(new_n335_), .B2(new_n312_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n381_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n420_));
  AND2_X1   g219(.A1(new_n323_), .A2(new_n327_), .ZN(new_n421_));
  AOI22_X1  g220(.A1(new_n419_), .A2(new_n420_), .B1(new_n421_), .B2(new_n315_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n307_), .B1(new_n422_), .B2(new_n371_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n376_), .B1(new_n418_), .B2(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n404_), .B1(new_n424_), .B2(KEYINPUT100), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n371_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n371_), .B(new_n328_), .C1(new_n342_), .C2(new_n353_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT20), .ZN(new_n428_));
  OAI211_X1 g227(.A(KEYINPUT100), .B(new_n375_), .C1(new_n426_), .C2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n306_), .B1(new_n425_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT102), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n418_), .A2(new_n376_), .A3(new_n423_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT95), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n373_), .A2(new_n403_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(new_n375_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT95), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n418_), .A2(new_n438_), .A3(new_n423_), .A4(new_n376_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n435_), .A2(new_n305_), .A3(new_n437_), .A4(new_n439_), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n440_), .A2(KEYINPUT27), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n375_), .B1(new_n426_), .B2(new_n428_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT100), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n444_), .A2(new_n429_), .A3(new_n404_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n445_), .A2(KEYINPUT102), .A3(new_n306_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n433_), .A2(new_n441_), .A3(new_n446_), .ZN(new_n447_));
  XOR2_X1   g246(.A(G78gat), .B(G106gat), .Z(new_n448_));
  AND3_X1   g247(.A1(KEYINPUT91), .A2(G228gat), .A3(G233gat), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n372_), .B1(KEYINPUT90), .B2(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(G141gat), .A2(G148gat), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT3), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G141gat), .A2(G148gat), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT2), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n453_), .A2(new_n456_), .A3(new_n457_), .A4(new_n458_), .ZN(new_n459_));
  OR2_X1    g258(.A1(G155gat), .A2(G162gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G155gat), .A2(G162gat), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n459_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n460_), .B1(KEYINPUT1), .B2(new_n461_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT89), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n461_), .A2(new_n464_), .A3(KEYINPUT1), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n464_), .B1(new_n461_), .B2(KEYINPUT1), .ZN(new_n467_));
  NOR3_X1   g266(.A1(new_n463_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n451_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(new_n454_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n462_), .B1(new_n468_), .B2(new_n470_), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n471_), .A2(KEYINPUT29), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n450_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT91), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n371_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT90), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n471_), .A2(new_n476_), .A3(KEYINPUT29), .ZN(new_n477_));
  AOI22_X1  g276(.A1(new_n475_), .A2(new_n477_), .B1(G228gat), .B2(G233gat), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n448_), .B1(new_n473_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NOR3_X1   g279(.A1(new_n473_), .A2(new_n478_), .A3(new_n448_), .ZN(new_n481_));
  OR3_X1    g280(.A1(new_n471_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n482_));
  OAI21_X1  g281(.A(KEYINPUT28), .B1(new_n471_), .B2(KEYINPUT29), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G22gat), .B(G50gat), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  AND3_X1   g284(.A1(new_n482_), .A2(new_n483_), .A3(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n485_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n487_));
  OAI22_X1  g286(.A1(new_n480_), .A2(new_n481_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n481_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n486_), .A2(new_n487_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n489_), .A2(new_n490_), .A3(new_n479_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n488_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G127gat), .B(G134gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G113gat), .B(G120gat), .ZN(new_n494_));
  XOR2_X1   g293(.A(new_n493_), .B(new_n494_), .Z(new_n495_));
  NOR2_X1   g294(.A1(new_n463_), .A2(new_n467_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n470_), .B1(new_n496_), .B2(new_n465_), .ZN(new_n497_));
  AND3_X1   g296(.A1(new_n459_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n495_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n493_), .B(new_n494_), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n500_), .B(new_n462_), .C1(new_n468_), .C2(new_n470_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n499_), .A2(new_n501_), .A3(KEYINPUT4), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G225gat), .A2(G233gat), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT4), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n471_), .A2(new_n505_), .A3(new_n495_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n502_), .A2(new_n504_), .A3(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n499_), .A2(new_n501_), .A3(new_n503_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT98), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G1gat), .B(G29gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G57gat), .B(G85gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n499_), .A2(new_n501_), .A3(KEYINPUT98), .A4(new_n503_), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n507_), .A2(new_n510_), .A3(new_n515_), .A4(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT101), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n507_), .A2(new_n510_), .A3(new_n516_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n515_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n519_), .B(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n492_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n435_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n437_), .A2(new_n439_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n306_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(new_n440_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT27), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n447_), .A2(new_n524_), .A3(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n445_), .A2(KEYINPUT32), .A3(new_n305_), .ZN(new_n532_));
  NOR3_X1   g331(.A1(new_n426_), .A2(new_n428_), .A3(new_n375_), .ZN(new_n533_));
  AOI22_X1  g332(.A1(new_n533_), .A2(new_n438_), .B1(new_n375_), .B2(new_n436_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n305_), .A2(KEYINPUT32), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(new_n535_), .A3(new_n435_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n523_), .A2(new_n532_), .A3(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT99), .ZN(new_n538_));
  INV_X1    g337(.A(new_n517_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT33), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n499_), .A2(new_n501_), .A3(new_n504_), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n521_), .A2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n502_), .A2(new_n503_), .A3(new_n506_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n540_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n538_), .B1(new_n539_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n539_), .A2(KEYINPUT33), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n539_), .A2(new_n538_), .A3(KEYINPUT33), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n547_), .A2(new_n527_), .A3(new_n440_), .A4(new_n548_), .ZN(new_n549_));
  AND2_X1   g348(.A1(new_n537_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n492_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n531_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  XOR2_X1   g351(.A(KEYINPUT87), .B(G43gat), .Z(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(KEYINPUT86), .B(KEYINPUT30), .ZN(new_n555_));
  AND3_X1   g354(.A1(new_n401_), .A2(new_n402_), .A3(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n555_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n557_));
  NOR3_X1   g356(.A1(new_n556_), .A2(new_n557_), .A3(G99gat), .ZN(new_n558_));
  INV_X1    g357(.A(G99gat), .ZN(new_n559_));
  INV_X1    g358(.A(new_n555_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n560_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n401_), .A2(new_n402_), .A3(new_n555_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n559_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n554_), .B1(new_n558_), .B2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G227gat), .A2(G233gat), .ZN(new_n565_));
  INV_X1    g364(.A(G15gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(G71gat), .ZN(new_n568_));
  OAI21_X1  g367(.A(G99gat), .B1(new_n556_), .B2(new_n557_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n561_), .A2(new_n559_), .A3(new_n562_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n569_), .A2(new_n553_), .A3(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n564_), .A2(new_n568_), .A3(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT88), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n568_), .B1(new_n564_), .B2(new_n571_), .ZN(new_n575_));
  OAI21_X1  g374(.A(KEYINPUT31), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n564_), .A2(new_n571_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n568_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT31), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n579_), .A2(new_n573_), .A3(new_n572_), .A4(new_n580_), .ZN(new_n581_));
  AND3_X1   g380(.A1(new_n576_), .A2(new_n495_), .A3(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n495_), .B1(new_n576_), .B2(new_n581_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n552_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n582_), .A2(new_n583_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n447_), .A2(new_n492_), .A3(new_n530_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT103), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n447_), .A2(new_n530_), .A3(KEYINPUT103), .A4(new_n492_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n523_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n585_), .A2(new_n590_), .A3(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n300_), .B1(new_n584_), .B2(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n286_), .B1(new_n224_), .B2(new_n217_), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n594_), .A2(KEYINPUT69), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n225_), .A2(new_n280_), .A3(new_n226_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n594_), .A2(KEYINPUT69), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n595_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(G232gat), .A2(G233gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT34), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n600_), .A2(KEYINPUT35), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(KEYINPUT35), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n594_), .A2(new_n603_), .ZN(new_n604_));
  AOI22_X1  g403(.A1(new_n598_), .A2(new_n601_), .B1(new_n596_), .B2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT36), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G190gat), .B(G218gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT70), .ZN(new_n608_));
  XOR2_X1   g407(.A(G134gat), .B(G162gat), .Z(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n605_), .A2(new_n606_), .A3(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(KEYINPUT36), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n611_), .B1(new_n613_), .B2(new_n605_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(KEYINPUT37), .ZN(new_n615_));
  XNOR2_X1  g414(.A(KEYINPUT72), .B(KEYINPUT37), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n605_), .A2(KEYINPUT71), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n612_), .B1(new_n605_), .B2(KEYINPUT71), .ZN(new_n618_));
  OAI211_X1 g417(.A(new_n611_), .B(new_n616_), .C1(new_n617_), .C2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n615_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(G231gat), .A2(G233gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n276_), .B(new_n621_), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n233_), .B(KEYINPUT75), .Z(new_n623_));
  AND2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n622_), .A2(new_n623_), .ZN(new_n625_));
  XOR2_X1   g424(.A(G127gat), .B(G155gat), .Z(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT16), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G183gat), .B(G211gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(new_n629_));
  XOR2_X1   g428(.A(KEYINPUT76), .B(KEYINPUT17), .Z(new_n630_));
  NOR4_X1   g429(.A1(new_n624_), .A2(new_n625_), .A3(new_n629_), .A4(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n622_), .B(new_n234_), .ZN(new_n632_));
  XOR2_X1   g431(.A(new_n629_), .B(KEYINPUT17), .Z(new_n633_));
  NOR2_X1   g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n631_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n620_), .A2(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT77), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n593_), .A2(new_n637_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n638_), .A2(new_n591_), .A3(new_n267_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n639_), .A2(KEYINPUT38), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT104), .Z(new_n641_));
  AOI21_X1  g440(.A(KEYINPUT27), .B1(new_n527_), .B2(new_n440_), .ZN(new_n642_));
  AOI21_X1  g441(.A(KEYINPUT102), .B1(new_n445_), .B2(new_n306_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n440_), .A2(KEYINPUT27), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n642_), .B1(new_n645_), .B2(new_n446_), .ZN(new_n646_));
  AOI21_X1  g445(.A(KEYINPUT103), .B1(new_n646_), .B2(new_n492_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n589_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n576_), .A2(new_n581_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(new_n500_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n576_), .A2(new_n495_), .A3(new_n581_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n651_), .A2(new_n591_), .A3(new_n652_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n584_), .B1(new_n649_), .B2(new_n653_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n611_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n300_), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n656_), .A2(new_n657_), .A3(new_n635_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(new_n523_), .ZN(new_n659_));
  AOI22_X1  g458(.A1(KEYINPUT38), .A2(new_n639_), .B1(new_n659_), .B2(G1gat), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n641_), .A2(new_n660_), .ZN(G1324gat));
  OR3_X1    g460(.A1(new_n638_), .A2(new_n646_), .A3(new_n268_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n646_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n658_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT39), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n664_), .A2(new_n665_), .A3(G8gat), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n665_), .B1(new_n664_), .B2(G8gat), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n662_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  XOR2_X1   g467(.A(new_n668_), .B(KEYINPUT40), .Z(G1325gat));
  NAND2_X1  g468(.A1(new_n658_), .A2(new_n585_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(G15gat), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(KEYINPUT105), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT105), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n670_), .A2(new_n673_), .A3(G15gat), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n672_), .A2(KEYINPUT41), .A3(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n585_), .A2(new_n566_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n675_), .B1(new_n638_), .B2(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(KEYINPUT41), .B1(new_n672_), .B2(new_n674_), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1326gat));
  OR3_X1    g478(.A1(new_n638_), .A2(G22gat), .A3(new_n492_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n658_), .A2(new_n551_), .ZN(new_n681_));
  XOR2_X1   g480(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n682_));
  AND3_X1   g481(.A1(new_n681_), .A2(G22gat), .A3(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n682_), .B1(new_n681_), .B2(G22gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n680_), .B1(new_n683_), .B2(new_n684_), .ZN(G1327gat));
  OR2_X1    g484(.A1(new_n655_), .A2(new_n635_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n593_), .A2(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(G29gat), .B1(new_n688_), .B2(new_n523_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n300_), .A2(new_n635_), .ZN(new_n690_));
  AOI211_X1 g489(.A(KEYINPUT43), .B(new_n620_), .C1(new_n592_), .C2(new_n584_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT43), .ZN(new_n692_));
  INV_X1    g491(.A(new_n620_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n692_), .B1(new_n654_), .B2(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n690_), .B1(new_n691_), .B2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  OAI211_X1 g497(.A(KEYINPUT44), .B(new_n690_), .C1(new_n691_), .C2(new_n694_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n698_), .A2(new_n700_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n523_), .A2(G29gat), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n689_), .B1(new_n701_), .B2(new_n702_), .ZN(G1328gat));
  INV_X1    g502(.A(KEYINPUT46), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n646_), .A2(G36gat), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n657_), .A2(new_n654_), .A3(new_n687_), .A4(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT45), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n706_), .B(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n697_), .A2(new_n663_), .A3(new_n699_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n708_), .B1(new_n709_), .B2(G36gat), .ZN(new_n710_));
  OAI211_X1 g509(.A(KEYINPUT108), .B(new_n704_), .C1(new_n710_), .C2(KEYINPUT107), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n709_), .A2(G36gat), .ZN(new_n713_));
  INV_X1    g512(.A(new_n708_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT107), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n712_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(KEYINPUT46), .B1(new_n710_), .B2(KEYINPUT108), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n711_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(G1329gat));
  NAND3_X1  g519(.A1(new_n593_), .A2(new_n585_), .A3(new_n687_), .ZN(new_n721_));
  INV_X1    g520(.A(G43gat), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT110), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT109), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n585_), .A2(G43gat), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n725_), .B1(new_n701_), .B2(new_n727_), .ZN(new_n728_));
  NOR4_X1   g527(.A1(new_n698_), .A2(new_n700_), .A3(KEYINPUT109), .A4(new_n726_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n724_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT47), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT47), .ZN(new_n732_));
  OAI211_X1 g531(.A(new_n732_), .B(new_n724_), .C1(new_n728_), .C2(new_n729_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(G1330gat));
  INV_X1    g533(.A(G50gat), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n688_), .A2(new_n735_), .A3(new_n551_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT111), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n697_), .A2(new_n737_), .A3(new_n551_), .A4(new_n699_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n738_), .A2(G50gat), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n697_), .A2(new_n551_), .A3(new_n699_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT111), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n739_), .A2(KEYINPUT112), .A3(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(KEYINPUT112), .B1(new_n739_), .B2(new_n741_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n736_), .B1(new_n742_), .B2(new_n743_), .ZN(G1331gat));
  NAND2_X1  g543(.A1(new_n262_), .A2(new_n266_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n637_), .A2(new_n745_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT113), .Z(new_n747_));
  INV_X1    g546(.A(new_n299_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n654_), .A2(new_n748_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT114), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n747_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(G57gat), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n752_), .A2(new_n753_), .A3(new_n523_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n745_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n755_), .A2(new_n299_), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n756_), .A2(new_n635_), .A3(new_n656_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n757_), .A2(new_n523_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n754_), .B1(new_n753_), .B2(new_n758_), .ZN(G1332gat));
  INV_X1    g558(.A(G64gat), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n663_), .A2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT48), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n757_), .A2(new_n663_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n762_), .B1(new_n763_), .B2(G64gat), .ZN(new_n764_));
  AOI211_X1 g563(.A(KEYINPUT48), .B(new_n760_), .C1(new_n757_), .C2(new_n663_), .ZN(new_n765_));
  OAI22_X1  g564(.A1(new_n751_), .A2(new_n761_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT115), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n766_), .B(new_n767_), .ZN(G1333gat));
  INV_X1    g567(.A(G71gat), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n769_), .B1(new_n757_), .B2(new_n585_), .ZN(new_n770_));
  XOR2_X1   g569(.A(new_n770_), .B(KEYINPUT49), .Z(new_n771_));
  NAND2_X1  g570(.A1(new_n585_), .A2(new_n769_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n771_), .B1(new_n751_), .B2(new_n772_), .ZN(G1334gat));
  INV_X1    g572(.A(G78gat), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n774_), .B1(new_n757_), .B2(new_n551_), .ZN(new_n775_));
  XOR2_X1   g574(.A(new_n775_), .B(KEYINPUT50), .Z(new_n776_));
  NAND2_X1  g575(.A1(new_n551_), .A2(new_n774_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n776_), .B1(new_n751_), .B2(new_n777_), .ZN(G1335gat));
  NOR2_X1   g577(.A1(new_n755_), .A2(new_n686_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n750_), .A2(KEYINPUT116), .A3(new_n779_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n749_), .A2(KEYINPUT114), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT114), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n782_), .B1(new_n654_), .B2(new_n748_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n779_), .B1(new_n781_), .B2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT116), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n780_), .A2(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(G85gat), .B1(new_n787_), .B2(new_n523_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT117), .ZN(new_n789_));
  OR2_X1    g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n789_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n654_), .A2(new_n693_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT43), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n654_), .A2(new_n692_), .A3(new_n693_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n635_), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n795_), .A2(new_n796_), .A3(new_n756_), .ZN(new_n797_));
  XOR2_X1   g596(.A(new_n797_), .B(KEYINPUT118), .Z(new_n798_));
  AND2_X1   g597(.A1(new_n523_), .A2(G85gat), .ZN(new_n799_));
  AOI22_X1  g598(.A1(new_n790_), .A2(new_n791_), .B1(new_n798_), .B2(new_n799_), .ZN(G1336gat));
  AOI21_X1  g599(.A(G92gat), .B1(new_n787_), .B2(new_n663_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT119), .ZN(new_n802_));
  OR2_X1    g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n801_), .A2(new_n802_), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n663_), .A2(G92gat), .ZN(new_n805_));
  AOI22_X1  g604(.A1(new_n803_), .A2(new_n804_), .B1(new_n798_), .B2(new_n805_), .ZN(G1337gat));
  AOI21_X1  g605(.A(new_n559_), .B1(new_n797_), .B2(new_n585_), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n585_), .A2(new_n218_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n807_), .B1(new_n787_), .B2(new_n808_), .ZN(new_n809_));
  XOR2_X1   g608(.A(new_n809_), .B(KEYINPUT51), .Z(G1338gat));
  NAND4_X1  g609(.A1(new_n795_), .A2(new_n551_), .A3(new_n796_), .A4(new_n756_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(G106gat), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(KEYINPUT52), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n811_), .A2(new_n814_), .A3(G106gat), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n813_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT120), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n492_), .A2(G106gat), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n817_), .B1(new_n787_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n818_), .ZN(new_n820_));
  AOI211_X1 g619(.A(KEYINPUT120), .B(new_n820_), .C1(new_n780_), .C2(new_n786_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n816_), .B1(new_n819_), .B2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(KEYINPUT53), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT53), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n824_), .B(new_n816_), .C1(new_n819_), .C2(new_n821_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n823_), .A2(new_n825_), .ZN(G1339gat));
  AND3_X1   g625(.A1(new_n585_), .A2(new_n590_), .A3(new_n523_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(KEYINPUT122), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n281_), .A2(new_n282_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n287_), .A2(new_n288_), .A3(new_n283_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n829_), .A2(new_n296_), .A3(new_n830_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n298_), .A2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n256_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT55), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n834_), .B1(new_n253_), .B2(new_n244_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n253_), .A2(new_n244_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n253_), .A2(new_n834_), .A3(new_n244_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n250_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT56), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  OAI211_X1 g640(.A(KEYINPUT56), .B(new_n250_), .C1(new_n837_), .C2(new_n838_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n833_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n693_), .B1(KEYINPUT58), .B2(new_n843_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n843_), .A2(KEYINPUT58), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n832_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n847_), .B1(new_n265_), .B2(new_n259_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n256_), .A2(new_n299_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n849_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n655_), .B1(new_n848_), .B2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(KEYINPUT121), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n846_), .B1(KEYINPUT57), .B2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n851_), .A2(KEYINPUT121), .A3(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n635_), .B1(new_n853_), .B2(new_n855_), .ZN(new_n856_));
  AOI211_X1 g655(.A(new_n299_), .B(new_n796_), .C1(new_n615_), .C2(new_n619_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n857_), .A2(new_n262_), .A3(new_n266_), .ZN(new_n858_));
  XOR2_X1   g657(.A(new_n858_), .B(KEYINPUT54), .Z(new_n859_));
  OAI21_X1  g658(.A(new_n828_), .B1(new_n856_), .B2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(G113gat), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n861_), .A2(new_n862_), .A3(new_n299_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT59), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n852_), .A2(KEYINPUT57), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n865_), .B(new_n855_), .C1(new_n845_), .C2(new_n844_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n859_), .B1(new_n866_), .B2(new_n796_), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n860_), .B(new_n864_), .C1(KEYINPUT123), .C2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n796_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n859_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT123), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n871_), .B(new_n828_), .C1(new_n872_), .C2(KEYINPUT59), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n748_), .B1(new_n868_), .B2(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n863_), .B1(new_n874_), .B2(new_n862_), .ZN(G1340gat));
  INV_X1    g674(.A(G120gat), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n876_), .B1(new_n755_), .B2(KEYINPUT60), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n861_), .B(new_n877_), .C1(KEYINPUT60), .C2(new_n876_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n755_), .B1(new_n868_), .B2(new_n873_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n879_), .B2(new_n876_), .ZN(G1341gat));
  INV_X1    g679(.A(G127gat), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n861_), .A2(new_n881_), .A3(new_n635_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n796_), .B1(new_n868_), .B2(new_n873_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n883_), .B2(new_n881_), .ZN(G1342gat));
  NAND2_X1  g683(.A1(new_n868_), .A2(new_n873_), .ZN(new_n885_));
  INV_X1    g684(.A(G134gat), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n620_), .A2(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n860_), .B2(new_n655_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(KEYINPUT124), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT124), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n890_), .B(new_n886_), .C1(new_n860_), .C2(new_n655_), .ZN(new_n891_));
  AOI22_X1  g690(.A1(new_n885_), .A2(new_n887_), .B1(new_n889_), .B2(new_n891_), .ZN(G1343gat));
  NOR4_X1   g691(.A1(new_n585_), .A2(new_n591_), .A3(new_n492_), .A4(new_n663_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n871_), .A2(new_n893_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n894_), .A2(new_n748_), .ZN(new_n895_));
  XOR2_X1   g694(.A(KEYINPUT125), .B(G141gat), .Z(new_n896_));
  XNOR2_X1  g695(.A(new_n895_), .B(new_n896_), .ZN(G1344gat));
  NAND3_X1  g696(.A1(new_n871_), .A2(new_n745_), .A3(new_n893_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g698(.A1(new_n894_), .A2(new_n796_), .ZN(new_n900_));
  XOR2_X1   g699(.A(KEYINPUT61), .B(G155gat), .Z(new_n901_));
  XNOR2_X1  g700(.A(new_n900_), .B(new_n901_), .ZN(G1346gat));
  OAI21_X1  g701(.A(G162gat), .B1(new_n894_), .B2(new_n620_), .ZN(new_n903_));
  OR2_X1    g702(.A1(new_n655_), .A2(G162gat), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n903_), .B1(new_n894_), .B2(new_n904_), .ZN(G1347gat));
  NOR2_X1   g704(.A1(new_n653_), .A2(new_n551_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n871_), .A2(new_n663_), .A3(new_n906_), .ZN(new_n907_));
  OAI21_X1  g706(.A(G169gat), .B1(new_n907_), .B2(new_n748_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT62), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n907_), .A2(new_n748_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n335_), .ZN(new_n912_));
  OAI211_X1 g711(.A(KEYINPUT62), .B(G169gat), .C1(new_n907_), .C2(new_n748_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n910_), .A2(new_n912_), .A3(new_n913_), .ZN(G1348gat));
  NOR2_X1   g713(.A1(new_n907_), .A2(new_n755_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(new_n312_), .ZN(G1349gat));
  NAND4_X1  g715(.A1(new_n871_), .A2(new_n663_), .A3(new_n635_), .A4(new_n906_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n917_), .A2(new_n326_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n918_), .B1(new_n351_), .B2(new_n917_), .ZN(G1350gat));
  OAI21_X1  g718(.A(G190gat), .B1(new_n907_), .B2(new_n620_), .ZN(new_n920_));
  OAI211_X1 g719(.A(new_n325_), .B(new_n611_), .C1(new_n617_), .C2(new_n618_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n920_), .B1(new_n907_), .B2(new_n921_), .ZN(G1351gat));
  INV_X1    g721(.A(KEYINPUT126), .ZN(new_n923_));
  NOR3_X1   g722(.A1(new_n585_), .A2(new_n523_), .A3(new_n492_), .ZN(new_n924_));
  NAND4_X1  g723(.A1(new_n871_), .A2(new_n663_), .A3(new_n299_), .A4(new_n924_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n923_), .B1(new_n925_), .B2(new_n357_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n924_), .ZN(new_n927_));
  NOR3_X1   g726(.A1(new_n867_), .A2(new_n646_), .A3(new_n927_), .ZN(new_n928_));
  NAND4_X1  g727(.A1(new_n928_), .A2(KEYINPUT126), .A3(G197gat), .A4(new_n299_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n925_), .A2(new_n357_), .ZN(new_n930_));
  AND3_X1   g729(.A1(new_n926_), .A2(new_n929_), .A3(new_n930_), .ZN(G1352gat));
  NAND2_X1  g730(.A1(new_n928_), .A2(new_n745_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g732(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n934_));
  AND2_X1   g733(.A1(new_n934_), .A2(KEYINPUT127), .ZN(new_n935_));
  AOI211_X1 g734(.A(new_n935_), .B(new_n796_), .C1(KEYINPUT63), .C2(G211gat), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n928_), .A2(new_n936_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n934_), .A2(KEYINPUT127), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n937_), .B(new_n938_), .ZN(G1354gat));
  INV_X1    g738(.A(new_n928_), .ZN(new_n940_));
  OAI21_X1  g739(.A(G218gat), .B1(new_n940_), .B2(new_n620_), .ZN(new_n941_));
  OR2_X1    g740(.A1(new_n655_), .A2(G218gat), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n941_), .B1(new_n940_), .B2(new_n942_), .ZN(G1355gat));
endmodule


