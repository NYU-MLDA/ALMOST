//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0 1 1 1 1 1 1 1 0 1 1 1 0 1 1 0 1 1 0 0 1 0 0 1 0 0 0 0 1 0 0 0 0 0 1 1 0 1 0 0 0 0 1 0 0 1 1 0 0 1 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n691_, new_n692_,
    new_n693_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n800_, new_n801_,
    new_n802_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n821_, new_n822_,
    new_n823_, new_n825_, new_n826_, new_n827_, new_n829_, new_n830_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n842_, new_n843_, new_n844_,
    new_n846_, new_n847_, new_n849_, new_n850_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_;
  INV_X1    g000(.A(KEYINPUT69), .ZN(new_n202_));
  NOR2_X1   g001(.A1(G99gat), .A2(G106gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  OAI22_X1  g004(.A1(KEYINPUT67), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  AND2_X1   g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT66), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n210_), .A2(KEYINPUT6), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT6), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n212_), .A2(KEYINPUT66), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n209_), .B1(new_n211_), .B2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(KEYINPUT66), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n210_), .A2(KEYINPUT6), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n215_), .A2(new_n216_), .A3(new_n208_), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n207_), .B1(new_n214_), .B2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(G85gat), .B(G92gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n202_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n219_), .ZN(new_n221_));
  AND3_X1   g020(.A1(new_n215_), .A2(new_n216_), .A3(new_n208_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n208_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  OAI211_X1 g023(.A(KEYINPUT69), .B(new_n221_), .C1(new_n224_), .C2(new_n207_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n220_), .A2(new_n225_), .A3(KEYINPUT8), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT70), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT68), .ZN(new_n228_));
  AOI21_X1  g027(.A(KEYINPUT8), .B1(new_n218_), .B2(new_n228_), .ZN(new_n229_));
  OAI211_X1 g028(.A(new_n229_), .B(new_n221_), .C1(new_n228_), .C2(new_n218_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT70), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n220_), .A2(new_n225_), .A3(new_n231_), .A4(KEYINPUT8), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n227_), .A2(new_n230_), .A3(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(G106gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT10), .B(G99gat), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT65), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n237_), .A2(G85gat), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT9), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n237_), .A2(new_n239_), .A3(G85gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n238_), .A2(new_n240_), .ZN(new_n241_));
  AOI22_X1  g040(.A1(new_n234_), .A2(new_n236_), .B1(new_n241_), .B2(G92gat), .ZN(new_n242_));
  OAI221_X1 g041(.A(new_n242_), .B1(new_n239_), .B2(new_n219_), .C1(new_n222_), .C2(new_n223_), .ZN(new_n243_));
  AND3_X1   g042(.A1(new_n233_), .A2(KEYINPUT71), .A3(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(KEYINPUT71), .B1(new_n233_), .B2(new_n243_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT73), .B(G43gat), .ZN(new_n247_));
  INV_X1    g046(.A(G50gat), .ZN(new_n248_));
  AND2_X1   g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n247_), .A2(new_n248_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G29gat), .B(G36gat), .ZN(new_n251_));
  OR3_X1    g050(.A1(new_n249_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n251_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(KEYINPUT74), .B1(new_n246_), .B2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT74), .ZN(new_n256_));
  INV_X1    g055(.A(new_n254_), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n256_), .B(new_n257_), .C1(new_n244_), .C2(new_n245_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n255_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n233_), .A2(new_n243_), .ZN(new_n260_));
  XOR2_X1   g059(.A(new_n254_), .B(KEYINPUT15), .Z(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G232gat), .A2(G233gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT34), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT35), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT75), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n259_), .A2(new_n262_), .A3(new_n268_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n265_), .A2(new_n266_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n270_), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n259_), .A2(new_n272_), .A3(new_n262_), .A4(new_n268_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT76), .B(G134gat), .ZN(new_n275_));
  INV_X1    g074(.A(G162gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G190gat), .B(G218gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT36), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n274_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT36), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n271_), .A2(new_n282_), .A3(new_n279_), .A4(new_n273_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n281_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT37), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n281_), .A2(KEYINPUT37), .A3(new_n283_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G15gat), .B(G22gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT77), .B(G8gat), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT14), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n289_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(G1gat), .ZN(new_n293_));
  INV_X1    g092(.A(G1gat), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n289_), .A2(new_n291_), .A3(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(G8gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G231gat), .A2(G233gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(G57gat), .B(G64gat), .Z(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT72), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT11), .ZN(new_n302_));
  XOR2_X1   g101(.A(G71gat), .B(G78gat), .Z(new_n303_));
  AND2_X1   g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT11), .ZN(new_n305_));
  NOR3_X1   g104(.A1(new_n301_), .A2(new_n305_), .A3(new_n303_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n299_), .B(new_n307_), .ZN(new_n308_));
  XOR2_X1   g107(.A(G127gat), .B(G155gat), .Z(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  XOR2_X1   g110(.A(G183gat), .B(G211gat), .Z(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT17), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  AND2_X1   g114(.A1(new_n313_), .A2(new_n314_), .ZN(new_n316_));
  NOR3_X1   g115(.A1(new_n308_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n317_), .B1(new_n315_), .B2(new_n308_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n288_), .A2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT79), .ZN(new_n321_));
  XOR2_X1   g120(.A(KEYINPUT26), .B(G190gat), .Z(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(KEYINPUT25), .B(G183gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(G169gat), .ZN(new_n326_));
  INV_X1    g125(.A(G176gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G169gat), .A2(G176gat), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n328_), .A2(KEYINPUT24), .A3(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n325_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT99), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G183gat), .A2(G190gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT23), .ZN(new_n334_));
  OR2_X1    g133(.A1(new_n328_), .A2(KEYINPUT24), .ZN(new_n335_));
  AND2_X1   g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n332_), .A2(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n334_), .B1(G183gat), .B2(G190gat), .ZN(new_n338_));
  INV_X1    g137(.A(new_n329_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT22), .B(G169gat), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n339_), .B1(new_n340_), .B2(new_n327_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n338_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n337_), .A2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT95), .B(G204gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT94), .B(G197gat), .ZN(new_n345_));
  AOI22_X1  g144(.A1(G197gat), .A2(new_n344_), .B1(new_n345_), .B2(G204gat), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT21), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT96), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  XOR2_X1   g149(.A(G211gat), .B(G218gat), .Z(new_n351_));
  OAI22_X1  g150(.A1(G197gat), .A2(new_n344_), .B1(new_n345_), .B2(G204gat), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n351_), .B1(new_n352_), .B2(KEYINPUT21), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n350_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n346_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n355_), .A2(KEYINPUT21), .A3(new_n351_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n354_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n343_), .A2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT84), .B(G190gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(KEYINPUT26), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n360_), .B1(KEYINPUT26), .B2(G190gat), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT83), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n361_), .B1(new_n362_), .B2(new_n324_), .ZN(new_n363_));
  INV_X1    g162(.A(G183gat), .ZN(new_n364_));
  AOI21_X1  g163(.A(KEYINPUT83), .B1(new_n364_), .B2(KEYINPUT25), .ZN(new_n365_));
  OAI211_X1 g164(.A(new_n336_), .B(new_n330_), .C1(new_n363_), .C2(new_n365_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n334_), .B1(G183gat), .B2(new_n359_), .ZN(new_n367_));
  OR2_X1    g166(.A1(new_n367_), .A2(KEYINPUT85), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(KEYINPUT85), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n368_), .A2(new_n341_), .A3(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n366_), .A2(new_n370_), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n358_), .B(KEYINPUT20), .C1(new_n357_), .C2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G226gat), .A2(G233gat), .ZN(new_n373_));
  XOR2_X1   g172(.A(new_n373_), .B(KEYINPUT98), .Z(new_n374_));
  XOR2_X1   g173(.A(new_n374_), .B(KEYINPUT19), .Z(new_n375_));
  NAND2_X1  g174(.A1(new_n372_), .A2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT18), .B(G64gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(G92gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G8gat), .B(G36gat), .ZN(new_n379_));
  XOR2_X1   g178(.A(new_n378_), .B(new_n379_), .Z(new_n380_));
  OR2_X1    g179(.A1(new_n343_), .A2(new_n357_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n375_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n357_), .A2(new_n371_), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n381_), .A2(KEYINPUT20), .A3(new_n382_), .A4(new_n383_), .ZN(new_n384_));
  AND3_X1   g183(.A1(new_n376_), .A2(new_n380_), .A3(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n380_), .B1(new_n376_), .B2(new_n384_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  XOR2_X1   g186(.A(G1gat), .B(G29gat), .Z(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT100), .B(KEYINPUT0), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  XOR2_X1   g189(.A(G57gat), .B(G85gat), .Z(new_n391_));
  XNOR2_X1  g190(.A(new_n390_), .B(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G127gat), .B(G134gat), .ZN(new_n393_));
  INV_X1    g192(.A(G113gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(G120gat), .ZN(new_n396_));
  NOR2_X1   g195(.A1(G141gat), .A2(G148gat), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G141gat), .A2(G148gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G155gat), .A2(G162gat), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT89), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n400_), .B(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(KEYINPUT1), .ZN(new_n403_));
  NOR2_X1   g202(.A1(G155gat), .A2(G162gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(KEYINPUT88), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n398_), .B(new_n399_), .C1(new_n403_), .C2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n399_), .A2(KEYINPUT90), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT2), .ZN(new_n409_));
  XOR2_X1   g208(.A(new_n397_), .B(KEYINPUT3), .Z(new_n410_));
  OAI211_X1 g209(.A(new_n405_), .B(new_n402_), .C1(new_n409_), .C2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n407_), .A2(KEYINPUT91), .A3(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(KEYINPUT91), .B1(new_n407_), .B2(new_n411_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n396_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT4), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n407_), .A2(new_n411_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n418_), .A2(new_n396_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n414_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(new_n412_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n419_), .B1(new_n421_), .B2(new_n396_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n417_), .B1(new_n422_), .B2(new_n416_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G225gat), .A2(G233gat), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n392_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n419_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n415_), .A2(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n425_), .B1(new_n424_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT33), .ZN(new_n429_));
  INV_X1    g228(.A(new_n424_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n427_), .A2(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n431_), .B1(new_n423_), .B2(new_n430_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n429_), .B1(new_n432_), .B2(new_n392_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n416_), .B1(new_n415_), .B2(new_n426_), .ZN(new_n434_));
  AOI21_X1  g233(.A(KEYINPUT4), .B1(new_n421_), .B2(new_n396_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n430_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n431_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n436_), .A2(new_n437_), .A3(new_n392_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n438_), .A2(KEYINPUT33), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n387_), .B(new_n428_), .C1(new_n433_), .C2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(KEYINPUT101), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n380_), .A2(KEYINPUT32), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n376_), .A2(new_n384_), .A3(new_n442_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n372_), .A2(new_n375_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n381_), .A2(KEYINPUT20), .A3(new_n383_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n444_), .B1(new_n375_), .B2(new_n445_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n432_), .A2(new_n392_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n438_), .ZN(new_n448_));
  OAI221_X1 g247(.A(new_n443_), .B1(new_n446_), .B2(new_n442_), .C1(new_n447_), .C2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n432_), .A2(new_n429_), .A3(new_n392_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n438_), .A2(KEYINPUT33), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT101), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n452_), .A2(new_n453_), .A3(new_n387_), .A4(new_n428_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n441_), .A2(new_n449_), .A3(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G228gat), .A2(G233gat), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n413_), .A2(new_n414_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT29), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n456_), .B(new_n357_), .C1(new_n457_), .C2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n357_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n460_), .B1(KEYINPUT29), .B2(new_n418_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n459_), .B1(new_n461_), .B2(new_n456_), .ZN(new_n462_));
  XOR2_X1   g261(.A(G78gat), .B(G106gat), .Z(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  AND2_X1   g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n462_), .A2(new_n464_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT97), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n468_), .B1(new_n462_), .B2(new_n464_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n457_), .A2(new_n458_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(KEYINPUT92), .B(KEYINPUT28), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT93), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n472_), .B(G22gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(G50gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n470_), .B(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n469_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n467_), .A2(new_n476_), .ZN(new_n477_));
  OAI22_X1  g276(.A1(new_n465_), .A2(new_n466_), .B1(new_n469_), .B2(new_n475_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n371_), .B(KEYINPUT30), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT87), .ZN(new_n482_));
  XOR2_X1   g281(.A(G15gat), .B(G43gat), .Z(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT86), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G71gat), .B(G99gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G227gat), .A2(G233gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n485_), .B(new_n486_), .ZN(new_n487_));
  XOR2_X1   g286(.A(new_n484_), .B(new_n487_), .Z(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n482_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n481_), .A2(KEYINPUT87), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(new_n488_), .ZN(new_n492_));
  XOR2_X1   g291(.A(new_n396_), .B(KEYINPUT31), .Z(new_n493_));
  AND3_X1   g292(.A1(new_n490_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n493_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n455_), .A2(new_n480_), .A3(new_n497_), .ZN(new_n498_));
  OR2_X1    g297(.A1(new_n387_), .A2(KEYINPUT27), .ZN(new_n499_));
  INV_X1    g298(.A(new_n385_), .ZN(new_n500_));
  XOR2_X1   g299(.A(new_n380_), .B(KEYINPUT102), .Z(new_n501_));
  OAI211_X1 g300(.A(new_n500_), .B(KEYINPUT27), .C1(new_n446_), .C2(new_n501_), .ZN(new_n502_));
  AND2_X1   g301(.A1(new_n499_), .A2(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n447_), .A2(new_n448_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n479_), .A2(new_n497_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n496_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n503_), .B(new_n504_), .C1(new_n505_), .C2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n498_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G229gat), .A2(G233gat), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n254_), .B(KEYINPUT80), .ZN(new_n511_));
  OAI21_X1  g310(.A(KEYINPUT81), .B1(new_n511_), .B2(new_n297_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT80), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n254_), .B(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT81), .ZN(new_n515_));
  INV_X1    g314(.A(new_n297_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n514_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n512_), .A2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n511_), .A2(new_n297_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n518_), .A2(KEYINPUT82), .A3(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(KEYINPUT82), .B1(new_n518_), .B2(new_n519_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n510_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n261_), .A2(new_n297_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n518_), .A2(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n525_), .A2(new_n510_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G113gat), .B(G141gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(new_n326_), .ZN(new_n529_));
  INV_X1    g328(.A(G197gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n523_), .A2(new_n527_), .A3(new_n532_), .ZN(new_n533_));
  NOR3_X1   g332(.A1(new_n511_), .A2(KEYINPUT81), .A3(new_n297_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n515_), .B1(new_n514_), .B2(new_n516_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n519_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT82), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n509_), .B1(new_n538_), .B2(new_n520_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n531_), .B1(new_n539_), .B2(new_n526_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n533_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT71), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n260_), .A2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n233_), .A2(KEYINPUT71), .A3(new_n243_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n544_), .A2(new_n545_), .A3(new_n307_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT12), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G230gat), .A2(G233gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT64), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n307_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n552_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n260_), .A2(new_n307_), .A3(KEYINPUT12), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n548_), .A2(new_n551_), .A3(new_n553_), .A4(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n546_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(new_n550_), .ZN(new_n557_));
  XOR2_X1   g356(.A(G120gat), .B(G148gat), .Z(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(G204gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT5), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(new_n327_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n555_), .A2(new_n557_), .A3(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n561_), .B1(new_n555_), .B2(new_n557_), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n565_), .A2(KEYINPUT13), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(KEYINPUT13), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n542_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  AND2_X1   g367(.A1(new_n508_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n321_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT103), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n504_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n321_), .A2(KEYINPUT103), .A3(new_n569_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n572_), .A2(new_n294_), .A3(new_n573_), .A4(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT38), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT105), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n575_), .A2(new_n576_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n284_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n581_), .A2(new_n319_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n569_), .A2(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT104), .ZN(new_n584_));
  OAI21_X1  g383(.A(G1gat), .B1(new_n584_), .B2(new_n504_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n575_), .A2(KEYINPUT105), .A3(new_n576_), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n579_), .A2(new_n580_), .A3(new_n585_), .A4(new_n586_), .ZN(G1324gat));
  OAI21_X1  g386(.A(G8gat), .B1(new_n583_), .B2(new_n503_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT107), .ZN(new_n589_));
  OR3_X1    g388(.A1(new_n588_), .A2(new_n589_), .A3(KEYINPUT39), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(KEYINPUT39), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(KEYINPUT106), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT106), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n588_), .A2(new_n593_), .A3(KEYINPUT39), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n589_), .B1(new_n588_), .B2(KEYINPUT39), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n590_), .A2(new_n592_), .A3(new_n594_), .A4(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n290_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n503_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n572_), .A2(new_n597_), .A3(new_n598_), .A4(new_n574_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n596_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT40), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(G1325gat));
  INV_X1    g401(.A(KEYINPUT41), .ZN(new_n603_));
  OAI21_X1  g402(.A(G15gat), .B1(new_n584_), .B2(new_n497_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(KEYINPUT108), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n604_), .A2(KEYINPUT108), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n603_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n607_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n609_), .A2(KEYINPUT41), .A3(new_n605_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n572_), .A2(new_n574_), .ZN(new_n611_));
  INV_X1    g410(.A(G15gat), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n611_), .A2(new_n612_), .A3(new_n496_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n608_), .A2(new_n610_), .A3(new_n613_), .ZN(G1326gat));
  XOR2_X1   g413(.A(new_n479_), .B(KEYINPUT109), .Z(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(G22gat), .B1(new_n584_), .B2(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT42), .ZN(new_n618_));
  INV_X1    g417(.A(G22gat), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n611_), .A2(new_n619_), .A3(new_n615_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n620_), .ZN(G1327gat));
  NOR2_X1   g420(.A1(new_n284_), .A2(new_n318_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n508_), .A2(new_n568_), .A3(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT111), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n508_), .A2(new_n568_), .A3(KEYINPUT111), .A4(new_n622_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(G29gat), .B1(new_n627_), .B2(new_n573_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT43), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n508_), .A2(new_n288_), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT110), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n288_), .A2(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n286_), .A2(KEYINPUT110), .A3(new_n287_), .ZN(new_n633_));
  AOI22_X1  g432(.A1(new_n632_), .A2(new_n633_), .B1(new_n507_), .B2(new_n498_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n630_), .B1(new_n634_), .B2(new_n629_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n635_), .A2(new_n568_), .A3(new_n319_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT44), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n635_), .A2(KEYINPUT44), .A3(new_n568_), .A4(new_n319_), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n638_), .A2(new_n573_), .A3(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n628_), .B1(new_n640_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g440(.A(G36gat), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n625_), .A2(new_n642_), .A3(new_n598_), .A4(new_n626_), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n643_), .A2(KEYINPUT112), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n643_), .A2(KEYINPUT112), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT45), .ZN(new_n646_));
  NOR3_X1   g445(.A1(new_n644_), .A2(new_n645_), .A3(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT112), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n627_), .A2(new_n648_), .A3(new_n642_), .A4(new_n598_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n643_), .A2(KEYINPUT112), .ZN(new_n650_));
  AOI21_X1  g449(.A(KEYINPUT45), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n647_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n638_), .A2(new_n598_), .A3(new_n639_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(G36gat), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n652_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT46), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n652_), .A2(new_n654_), .A3(KEYINPUT46), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(G1329gat));
  NAND4_X1  g458(.A1(new_n638_), .A2(G43gat), .A3(new_n496_), .A4(new_n639_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n627_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n661_), .A2(new_n497_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n660_), .B1(G43gat), .B2(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g463(.A1(new_n638_), .A2(G50gat), .A3(new_n479_), .A4(new_n639_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n248_), .B1(new_n661_), .B2(new_n616_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n665_), .A2(new_n666_), .ZN(G1331gat));
  NAND2_X1  g466(.A1(new_n508_), .A2(new_n542_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT113), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n566_), .A2(new_n567_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n669_), .A2(new_n671_), .A3(new_n321_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(G57gat), .B1(new_n673_), .B2(new_n573_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n670_), .A2(new_n541_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n675_), .A2(new_n508_), .A3(new_n582_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n677_), .A2(G57gat), .A3(new_n573_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT114), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n674_), .A2(new_n679_), .ZN(G1332gat));
  OAI21_X1  g479(.A(G64gat), .B1(new_n676_), .B2(new_n503_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT48), .ZN(new_n682_));
  OR2_X1    g481(.A1(new_n503_), .A2(G64gat), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n682_), .B1(new_n672_), .B2(new_n683_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT115), .ZN(G1333gat));
  OAI21_X1  g484(.A(G71gat), .B1(new_n676_), .B2(new_n497_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT49), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n497_), .A2(G71gat), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n687_), .B1(new_n672_), .B2(new_n688_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT116), .ZN(G1334gat));
  OAI21_X1  g489(.A(G78gat), .B1(new_n676_), .B2(new_n616_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT50), .ZN(new_n692_));
  OR2_X1    g491(.A1(new_n616_), .A2(G78gat), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n692_), .B1(new_n672_), .B2(new_n693_), .ZN(G1335gat));
  NAND3_X1  g493(.A1(new_n669_), .A2(new_n671_), .A3(new_n622_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(G85gat), .B1(new_n696_), .B2(new_n573_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n675_), .A2(new_n319_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT117), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n635_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT118), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(KEYINPUT118), .B1(new_n700_), .B2(new_n701_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n237_), .A2(G85gat), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n238_), .B1(new_n504_), .B2(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n697_), .B1(new_n706_), .B2(new_n708_), .ZN(G1336gat));
  AOI21_X1  g508(.A(G92gat), .B1(new_n696_), .B2(new_n598_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n503_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n711_), .B2(G92gat), .ZN(G1337gat));
  NAND2_X1  g511(.A1(new_n496_), .A2(new_n236_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n695_), .A2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n702_), .A2(new_n496_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n715_), .B2(G99gat), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT51), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n716_), .B(new_n717_), .ZN(G1338gat));
  NAND3_X1  g517(.A1(new_n699_), .A2(new_n635_), .A3(new_n479_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT52), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n719_), .A2(new_n720_), .A3(G106gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n719_), .B2(G106gat), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n479_), .A2(new_n234_), .ZN(new_n723_));
  OAI22_X1  g522(.A1(new_n721_), .A2(new_n722_), .B1(new_n695_), .B2(new_n723_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g524(.A(KEYINPUT55), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT120), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n550_), .B2(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(KEYINPUT12), .B1(new_n246_), .B2(new_n307_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n553_), .A2(new_n554_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n728_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n561_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n728_), .B1(new_n726_), .B2(new_n550_), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n548_), .A2(new_n553_), .A3(new_n554_), .A4(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n731_), .A2(new_n732_), .A3(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT56), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n731_), .A2(KEYINPUT56), .A3(new_n734_), .A4(new_n732_), .ZN(new_n738_));
  AND3_X1   g537(.A1(new_n737_), .A2(KEYINPUT121), .A3(new_n738_), .ZN(new_n739_));
  OAI211_X1 g538(.A(new_n541_), .B(new_n562_), .C1(KEYINPUT121), .C2(new_n738_), .ZN(new_n740_));
  OAI21_X1  g539(.A(KEYINPUT122), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n509_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n742_));
  OAI211_X1 g541(.A(new_n742_), .B(new_n531_), .C1(new_n509_), .C2(new_n525_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n743_), .A2(new_n533_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n565_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n738_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT121), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n563_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n737_), .A2(KEYINPUT121), .A3(new_n738_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT122), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n748_), .A2(new_n749_), .A3(new_n750_), .A4(new_n541_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n741_), .A2(new_n745_), .A3(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(new_n284_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT57), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n752_), .A2(KEYINPUT57), .A3(new_n284_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n737_), .A2(new_n738_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n757_), .A2(new_n562_), .A3(new_n744_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT58), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  OR2_X1    g559(.A1(new_n758_), .A2(new_n759_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n288_), .A2(new_n760_), .A3(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n755_), .A2(new_n756_), .A3(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT123), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n755_), .A2(KEYINPUT123), .A3(new_n756_), .A4(new_n762_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n765_), .A2(new_n319_), .A3(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n670_), .A2(new_n542_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(KEYINPUT119), .A2(KEYINPUT54), .ZN(new_n769_));
  NOR4_X1   g568(.A1(new_n768_), .A2(new_n288_), .A3(new_n319_), .A4(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n320_), .A2(new_n542_), .A3(new_n670_), .ZN(new_n771_));
  XOR2_X1   g570(.A(KEYINPUT119), .B(KEYINPUT54), .Z(new_n772_));
  AOI21_X1  g571(.A(new_n770_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n767_), .A2(new_n773_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n598_), .A2(new_n504_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n505_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n774_), .A2(new_n541_), .A3(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(new_n394_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n763_), .A2(new_n319_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n773_), .A2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT59), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n781_), .A2(new_n782_), .A3(new_n777_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n542_), .A2(new_n394_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n776_), .B1(new_n767_), .B2(new_n773_), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n783_), .B(new_n784_), .C1(new_n785_), .C2(new_n782_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n779_), .A2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(KEYINPUT124), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT124), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n779_), .A2(new_n786_), .A3(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n790_), .ZN(G1340gat));
  NAND2_X1  g590(.A1(new_n774_), .A2(new_n777_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT59), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n793_), .A2(new_n671_), .A3(new_n783_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(G120gat), .ZN(new_n795_));
  INV_X1    g594(.A(G120gat), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n796_), .B1(new_n670_), .B2(KEYINPUT60), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n785_), .B(new_n797_), .C1(KEYINPUT60), .C2(new_n796_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n795_), .A2(new_n798_), .ZN(G1341gat));
  AOI21_X1  g598(.A(G127gat), .B1(new_n785_), .B2(new_n318_), .ZN(new_n800_));
  OAI211_X1 g599(.A(G127gat), .B(new_n783_), .C1(new_n785_), .C2(new_n782_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n800_), .B1(new_n802_), .B2(new_n318_), .ZN(G1342gat));
  INV_X1    g602(.A(G134gat), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n804_), .B1(new_n792_), .B2(new_n284_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT125), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT125), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n807_), .B(new_n804_), .C1(new_n792_), .C2(new_n284_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n288_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n809_), .A2(new_n804_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n793_), .A2(new_n783_), .A3(new_n810_), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n806_), .A2(new_n808_), .A3(new_n811_), .ZN(G1343gat));
  NAND2_X1  g611(.A1(new_n774_), .A2(new_n506_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n775_), .ZN(new_n815_));
  OAI21_X1  g614(.A(G141gat), .B1(new_n815_), .B2(new_n542_), .ZN(new_n816_));
  NOR3_X1   g615(.A1(new_n813_), .A2(new_n504_), .A3(new_n598_), .ZN(new_n817_));
  INV_X1    g616(.A(G141gat), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n817_), .A2(new_n818_), .A3(new_n541_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n816_), .A2(new_n819_), .ZN(G1344gat));
  OAI21_X1  g619(.A(G148gat), .B1(new_n815_), .B2(new_n670_), .ZN(new_n821_));
  INV_X1    g620(.A(G148gat), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n817_), .A2(new_n822_), .A3(new_n671_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n823_), .ZN(G1345gat));
  NAND4_X1  g623(.A1(new_n774_), .A2(new_n506_), .A3(new_n318_), .A4(new_n775_), .ZN(new_n825_));
  XOR2_X1   g624(.A(KEYINPUT61), .B(G155gat), .Z(new_n826_));
  XNOR2_X1  g625(.A(new_n826_), .B(KEYINPUT126), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n825_), .B(new_n827_), .ZN(G1346gat));
  NAND2_X1  g627(.A1(new_n817_), .A2(new_n581_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n276_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n830_));
  AOI22_X1  g629(.A1(new_n829_), .A2(new_n276_), .B1(new_n817_), .B2(new_n830_), .ZN(G1347gat));
  INV_X1    g630(.A(KEYINPUT62), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n503_), .A2(new_n573_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n834_), .A2(new_n497_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n781_), .A2(new_n616_), .A3(new_n835_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n836_), .A2(new_n542_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n832_), .B1(new_n837_), .B2(new_n326_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n340_), .ZN(new_n839_));
  OAI211_X1 g638(.A(KEYINPUT62), .B(G169gat), .C1(new_n836_), .C2(new_n542_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n838_), .A2(new_n839_), .A3(new_n840_), .ZN(G1348gat));
  AOI21_X1  g640(.A(new_n479_), .B1(new_n767_), .B2(new_n773_), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n842_), .A2(G176gat), .A3(new_n671_), .A4(new_n835_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n327_), .B1(new_n836_), .B2(new_n670_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n843_), .A2(new_n844_), .ZN(G1349gat));
  NOR3_X1   g644(.A1(new_n836_), .A2(new_n324_), .A3(new_n319_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n842_), .A2(new_n318_), .A3(new_n835_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n846_), .B1(new_n364_), .B2(new_n847_), .ZN(G1350gat));
  OAI21_X1  g647(.A(G190gat), .B1(new_n836_), .B2(new_n809_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n581_), .A2(new_n323_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n849_), .B1(new_n836_), .B2(new_n850_), .ZN(G1351gat));
  XNOR2_X1  g650(.A(KEYINPUT127), .B(G197gat), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n814_), .A2(new_n833_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n853_), .B1(new_n854_), .B2(new_n542_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n813_), .A2(new_n834_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n856_), .A2(new_n541_), .A3(new_n852_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n857_), .ZN(G1352gat));
  OAI21_X1  g657(.A(G204gat), .B1(new_n854_), .B2(new_n670_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n856_), .A2(new_n671_), .A3(new_n344_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(G1353gat));
  OAI22_X1  g660(.A1(new_n854_), .A2(new_n319_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n862_));
  XNOR2_X1  g661(.A(KEYINPUT63), .B(G211gat), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n856_), .A2(new_n318_), .A3(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n864_), .ZN(G1354gat));
  NAND2_X1  g664(.A1(new_n856_), .A2(new_n581_), .ZN(new_n866_));
  INV_X1    g665(.A(G218gat), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n809_), .A2(new_n867_), .ZN(new_n868_));
  AOI22_X1  g667(.A1(new_n866_), .A2(new_n867_), .B1(new_n856_), .B2(new_n868_), .ZN(G1355gat));
endmodule


