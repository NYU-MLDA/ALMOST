//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 0 0 0 0 0 0 1 1 1 1 1 0 0 0 1 0 1 0 1 1 0 1 0 1 1 1 1 0 0 0 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n711_, new_n712_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n732_, new_n733_,
    new_n734_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n758_, new_n759_, new_n760_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n860_, new_n861_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n871_, new_n872_, new_n873_, new_n874_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n914_, new_n915_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n923_, new_n924_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n934_,
    new_n935_;
  INV_X1    g000(.A(G134gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(G127gat), .ZN(new_n203_));
  INV_X1    g002(.A(G127gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G134gat), .ZN(new_n205_));
  INV_X1    g004(.A(G120gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(G113gat), .ZN(new_n207_));
  INV_X1    g006(.A(G113gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(G120gat), .ZN(new_n209_));
  AND4_X1   g008(.A1(new_n203_), .A2(new_n205_), .A3(new_n207_), .A4(new_n209_), .ZN(new_n210_));
  AOI22_X1  g009(.A1(new_n203_), .A2(new_n205_), .B1(new_n207_), .B2(new_n209_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT31), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT24), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G183gat), .A2(G190gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT23), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT23), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n220_), .A2(G183gat), .A3(G190gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT79), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n219_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n218_), .ZN(new_n224_));
  AOI21_X1  g023(.A(KEYINPUT79), .B1(new_n224_), .B2(new_n220_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n217_), .B1(new_n223_), .B2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT80), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  OAI211_X1 g027(.A(KEYINPUT80), .B(new_n217_), .C1(new_n223_), .C2(new_n225_), .ZN(new_n229_));
  INV_X1    g028(.A(G183gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT25), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT25), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(G183gat), .ZN(new_n233_));
  INV_X1    g032(.A(G190gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT26), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT26), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(G190gat), .ZN(new_n237_));
  NAND4_X1  g036(.A1(new_n231_), .A2(new_n233_), .A3(new_n235_), .A4(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n215_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G169gat), .A2(G176gat), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(KEYINPUT24), .A3(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n238_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT78), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT78), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n238_), .A2(new_n241_), .A3(new_n244_), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n228_), .A2(new_n229_), .A3(new_n243_), .A4(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n219_), .A2(new_n221_), .A3(KEYINPUT81), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n230_), .A2(new_n234_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT81), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n224_), .A2(new_n249_), .A3(new_n220_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n247_), .A2(new_n248_), .A3(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT82), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n247_), .A2(new_n250_), .A3(KEYINPUT82), .A4(new_n248_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(KEYINPUT22), .B(G169gat), .ZN(new_n255_));
  INV_X1    g054(.A(G176gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  AND2_X1   g056(.A1(new_n257_), .A2(new_n240_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n253_), .A2(new_n254_), .A3(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n246_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G227gat), .A2(G233gat), .ZN(new_n261_));
  INV_X1    g060(.A(G71gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n261_), .B(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(G99gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n260_), .B(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G15gat), .B(G43gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT83), .ZN(new_n267_));
  XOR2_X1   g066(.A(new_n267_), .B(KEYINPUT30), .Z(new_n268_));
  XNOR2_X1  g067(.A(new_n265_), .B(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n214_), .B1(new_n269_), .B2(KEYINPUT84), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n270_), .B1(KEYINPUT84), .B2(new_n269_), .ZN(new_n271_));
  OR3_X1    g070(.A1(new_n269_), .A2(KEYINPUT84), .A3(new_n213_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(G155gat), .A2(G162gat), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G155gat), .A2(G162gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  OAI21_X1  g076(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NOR3_X1   g078(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n277_), .B1(new_n281_), .B2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(G141gat), .ZN(new_n287_));
  INV_X1    g086(.A(G148gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G141gat), .A2(G148gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n276_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT1), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n274_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n276_), .A2(KEYINPUT1), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n291_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n212_), .B1(new_n286_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT3), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n298_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT2), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n290_), .A2(new_n300_), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n299_), .A2(new_n301_), .A3(new_n282_), .A4(new_n278_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n302_), .A2(new_n276_), .A3(new_n275_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n203_), .A2(new_n205_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n207_), .A2(new_n209_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n203_), .A2(new_n205_), .A3(new_n207_), .A4(new_n209_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n293_), .A2(G155gat), .A3(G162gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n275_), .A2(new_n295_), .A3(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n310_), .A2(new_n290_), .A3(new_n289_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n303_), .A2(new_n308_), .A3(new_n311_), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n297_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G225gat), .A2(G233gat), .ZN(new_n314_));
  XOR2_X1   g113(.A(new_n314_), .B(KEYINPUT90), .Z(new_n315_));
  NOR2_X1   g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n297_), .A2(KEYINPUT4), .A3(new_n312_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT89), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n297_), .A2(new_n312_), .A3(KEYINPUT89), .A4(KEYINPUT4), .ZN(new_n320_));
  INV_X1    g119(.A(new_n297_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT4), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n319_), .A2(new_n320_), .A3(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n316_), .B1(new_n324_), .B2(new_n315_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G1gat), .B(G29gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G57gat), .B(G85gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT91), .B(KEYINPUT0), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n325_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n330_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n315_), .ZN(new_n333_));
  AOI22_X1  g132(.A1(new_n317_), .A2(new_n318_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n333_), .B1(new_n334_), .B2(new_n320_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n332_), .B1(new_n335_), .B2(new_n316_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n331_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT95), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT95), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n331_), .A2(new_n336_), .A3(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n273_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT27), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G8gat), .B(G36gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT18), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G64gat), .B(G92gat), .ZN(new_n348_));
  XOR2_X1   g147(.A(new_n347_), .B(new_n348_), .Z(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G226gat), .A2(G233gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT19), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n224_), .A2(KEYINPUT79), .A3(new_n220_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n221_), .A2(new_n222_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n353_), .A2(new_n354_), .A3(new_n219_), .ZN(new_n355_));
  AND2_X1   g154(.A1(new_n355_), .A2(new_n248_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n257_), .A2(new_n240_), .ZN(new_n357_));
  AND3_X1   g156(.A1(new_n240_), .A2(KEYINPUT88), .A3(KEYINPUT24), .ZN(new_n358_));
  AOI21_X1  g157(.A(KEYINPUT88), .B1(new_n240_), .B2(KEYINPUT24), .ZN(new_n359_));
  NOR3_X1   g158(.A1(new_n358_), .A2(new_n359_), .A3(new_n215_), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n238_), .A2(new_n247_), .A3(new_n250_), .A4(new_n217_), .ZN(new_n361_));
  OAI22_X1  g160(.A1(new_n356_), .A2(new_n357_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(G197gat), .ZN(new_n363_));
  INV_X1    g162(.A(G204gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G197gat), .A2(G204gat), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n365_), .A2(KEYINPUT21), .A3(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G211gat), .B(G218gat), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT86), .ZN(new_n369_));
  OR3_X1    g168(.A1(new_n367_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n369_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  AND2_X1   g171(.A1(new_n367_), .A2(new_n368_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n365_), .A2(new_n366_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT21), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n373_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n372_), .A2(new_n377_), .ZN(new_n378_));
  OAI21_X1  g177(.A(KEYINPUT20), .B1(new_n362_), .B2(new_n378_), .ZN(new_n379_));
  AOI22_X1  g178(.A1(new_n370_), .A2(new_n371_), .B1(new_n373_), .B2(new_n376_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n380_), .B1(new_n246_), .B2(new_n259_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n352_), .B1(new_n379_), .B2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT93), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  OAI211_X1 g183(.A(KEYINPUT93), .B(new_n352_), .C1(new_n379_), .C2(new_n381_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n243_), .A2(new_n229_), .A3(new_n245_), .ZN(new_n387_));
  AOI21_X1  g186(.A(KEYINPUT80), .B1(new_n355_), .B2(new_n217_), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n380_), .B(new_n259_), .C1(new_n387_), .C2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n389_), .A2(KEYINPUT87), .A3(KEYINPUT20), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n362_), .A2(new_n378_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(KEYINPUT87), .B1(new_n389_), .B2(KEYINPUT20), .ZN(new_n393_));
  NOR3_X1   g192(.A1(new_n392_), .A2(new_n352_), .A3(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n350_), .B1(new_n386_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT96), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n352_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n397_));
  OR3_X1    g196(.A1(new_n379_), .A2(new_n381_), .A3(new_n352_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n397_), .A2(new_n349_), .A3(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n395_), .A2(new_n396_), .A3(new_n399_), .ZN(new_n400_));
  AND2_X1   g199(.A1(new_n397_), .A2(new_n398_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n401_), .A2(KEYINPUT96), .A3(new_n349_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n345_), .B1(new_n400_), .B2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n397_), .A2(new_n398_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(new_n350_), .ZN(new_n405_));
  AOI21_X1  g204(.A(KEYINPUT27), .B1(new_n405_), .B2(new_n399_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n403_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n303_), .A2(new_n311_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(KEYINPUT29), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n378_), .A2(new_n409_), .ZN(new_n410_));
  XOR2_X1   g209(.A(G22gat), .B(G50gat), .Z(new_n411_));
  XOR2_X1   g210(.A(new_n410_), .B(new_n411_), .Z(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  OR3_X1    g212(.A1(new_n408_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n414_));
  OAI21_X1  g213(.A(KEYINPUT28), .B1(new_n408_), .B2(KEYINPUT29), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT85), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G228gat), .A2(G233gat), .ZN(new_n418_));
  INV_X1    g217(.A(G78gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(G106gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT85), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n414_), .A2(new_n424_), .A3(new_n415_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n417_), .A2(new_n423_), .A3(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n423_), .B1(new_n417_), .B2(new_n425_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n413_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n428_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n430_), .A2(new_n412_), .A3(new_n426_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n429_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n407_), .A2(KEYINPUT97), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n406_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n399_), .A2(new_n396_), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n399_), .A2(new_n396_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n436_), .B1(new_n437_), .B2(new_n395_), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n433_), .B(new_n435_), .C1(new_n438_), .C2(new_n345_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT97), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n344_), .B1(new_n434_), .B2(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT33), .B1(new_n325_), .B2(new_n330_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT33), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n444_), .B(new_n332_), .C1(new_n335_), .C2(new_n316_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n334_), .A2(new_n333_), .A3(new_n320_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n332_), .B1(new_n315_), .B2(new_n313_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n405_), .A2(new_n446_), .A3(new_n399_), .A4(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT92), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  AOI22_X1  g251(.A1(new_n443_), .A2(new_n445_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n453_), .A2(KEYINPUT92), .A3(new_n399_), .A4(new_n405_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n349_), .A2(KEYINPUT32), .ZN(new_n455_));
  AOI22_X1  g254(.A1(new_n401_), .A2(new_n455_), .B1(new_n336_), .B2(new_n331_), .ZN(new_n456_));
  OAI211_X1 g255(.A(KEYINPUT32), .B(new_n349_), .C1(new_n386_), .C2(new_n394_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n452_), .A2(new_n454_), .A3(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(new_n433_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT94), .ZN(new_n461_));
  AOI22_X1  g260(.A1(new_n450_), .A2(new_n451_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n432_), .B1(new_n462_), .B2(new_n454_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT94), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n341_), .A2(new_n432_), .ZN(new_n466_));
  OR3_X1    g265(.A1(new_n403_), .A2(new_n466_), .A3(new_n406_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n461_), .A2(new_n465_), .A3(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n442_), .B1(new_n468_), .B2(new_n273_), .ZN(new_n469_));
  XOR2_X1   g268(.A(G85gat), .B(G92gat), .Z(new_n470_));
  INV_X1    g269(.A(KEYINPUT64), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT9), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n470_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  XOR2_X1   g274(.A(KEYINPUT10), .B(G99gat), .Z(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(new_n421_), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n471_), .A2(new_n472_), .A3(G85gat), .A4(G92gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G99gat), .A2(G106gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT6), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT6), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n481_), .A2(G99gat), .A3(G106gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n475_), .A2(new_n477_), .A3(new_n478_), .A4(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT8), .ZN(new_n485_));
  AND3_X1   g284(.A1(new_n480_), .A2(new_n482_), .A3(KEYINPUT65), .ZN(new_n486_));
  AOI21_X1  g285(.A(KEYINPUT65), .B1(new_n480_), .B2(new_n482_), .ZN(new_n487_));
  OAI21_X1  g286(.A(KEYINPUT66), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT65), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n483_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT66), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n480_), .A2(new_n482_), .A3(KEYINPUT65), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n490_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(G99gat), .A2(G106gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT7), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n488_), .A2(new_n493_), .A3(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n485_), .B1(new_n496_), .B2(new_n470_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n470_), .A2(new_n485_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n498_), .B1(new_n483_), .B2(new_n495_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n484_), .B1(new_n497_), .B2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G29gat), .B(G36gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G43gat), .B(G50gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT15), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n500_), .A2(new_n504_), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n484_), .B(new_n503_), .C1(new_n497_), .C2(new_n499_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G232gat), .A2(G233gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT34), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n505_), .B(new_n506_), .C1(KEYINPUT35), .C2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(KEYINPUT35), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G190gat), .B(G218gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G134gat), .B(G162gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n514_), .A2(KEYINPUT36), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n511_), .A2(new_n515_), .ZN(new_n516_));
  XOR2_X1   g315(.A(new_n514_), .B(KEYINPUT36), .Z(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n516_), .B1(new_n511_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n469_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT11), .ZN(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT67), .B(G71gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(new_n419_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n523_), .A2(new_n419_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n522_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G57gat), .B(G64gat), .ZN(new_n528_));
  XOR2_X1   g327(.A(KEYINPUT67), .B(G71gat), .Z(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(G78gat), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n530_), .A2(KEYINPUT11), .A3(new_n524_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n527_), .A2(new_n528_), .A3(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n528_), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n530_), .A2(KEYINPUT11), .A3(new_n524_), .A4(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n532_), .A2(new_n534_), .ZN(new_n535_));
  OAI211_X1 g334(.A(new_n484_), .B(new_n535_), .C1(new_n497_), .C2(new_n499_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT68), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n535_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n500_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  AND2_X1   g340(.A1(G230gat), .A2(G233gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n536_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n544_), .A2(new_n542_), .ZN(new_n545_));
  AOI21_X1  g344(.A(KEYINPUT12), .B1(new_n540_), .B2(KEYINPUT69), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT69), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT12), .ZN(new_n548_));
  AOI211_X1 g347(.A(new_n547_), .B(new_n548_), .C1(new_n500_), .C2(new_n539_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n545_), .B1(new_n546_), .B2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n543_), .A2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G120gat), .B(G148gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT5), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G176gat), .B(G204gat), .ZN(new_n554_));
  XOR2_X1   g353(.A(new_n553_), .B(new_n554_), .Z(new_n555_));
  NAND2_X1  g354(.A1(new_n551_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n555_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n543_), .A2(new_n550_), .A3(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n556_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT13), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n556_), .A2(KEYINPUT13), .A3(new_n558_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G15gat), .B(G22gat), .ZN(new_n564_));
  INV_X1    g363(.A(G1gat), .ZN(new_n565_));
  INV_X1    g364(.A(G8gat), .ZN(new_n566_));
  OAI21_X1  g365(.A(KEYINPUT14), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n564_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G1gat), .B(G8gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G231gat), .A2(G233gat), .ZN(new_n571_));
  XOR2_X1   g370(.A(new_n570_), .B(new_n571_), .Z(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(new_n539_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  XOR2_X1   g373(.A(G127gat), .B(G155gat), .Z(new_n575_));
  XNOR2_X1  g374(.A(G183gat), .B(G211gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(KEYINPUT70), .B(KEYINPUT16), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n574_), .A2(KEYINPUT17), .A3(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT71), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n579_), .B(KEYINPUT17), .Z(new_n582_));
  NAND2_X1  g381(.A1(new_n573_), .A2(new_n582_), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n583_), .B(KEYINPUT72), .Z(new_n584_));
  NAND2_X1  g383(.A1(new_n581_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G229gat), .A2(G233gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n503_), .B(KEYINPUT74), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(new_n570_), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n588_), .A2(KEYINPUT75), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(KEYINPUT75), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n586_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n504_), .A2(new_n570_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT76), .ZN(new_n594_));
  INV_X1    g393(.A(new_n570_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n587_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n594_), .A2(new_n596_), .A3(new_n586_), .ZN(new_n597_));
  XOR2_X1   g396(.A(G113gat), .B(G141gat), .Z(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT77), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G169gat), .B(G197gat), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n599_), .B(new_n600_), .Z(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n592_), .A2(new_n597_), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n597_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n601_), .B1(new_n591_), .B2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n603_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NOR3_X1   g406(.A1(new_n563_), .A2(new_n585_), .A3(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n521_), .A2(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(G1gat), .B1(new_n609_), .B2(new_n341_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n519_), .A2(KEYINPUT37), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n519_), .A2(KEYINPUT37), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n585_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT73), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n617_), .A2(new_n563_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n469_), .A2(new_n607_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NOR3_X1   g419(.A1(new_n620_), .A2(G1gat), .A3(new_n341_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n621_), .A2(new_n622_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n610_), .B1(new_n623_), .B2(new_n624_), .ZN(G1324gat));
  INV_X1    g424(.A(KEYINPUT39), .ZN(new_n626_));
  INV_X1    g425(.A(new_n609_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n407_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n626_), .B1(new_n629_), .B2(G8gat), .ZN(new_n630_));
  AOI211_X1 g429(.A(KEYINPUT39), .B(new_n566_), .C1(new_n627_), .C2(new_n628_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n628_), .A2(new_n566_), .ZN(new_n632_));
  OAI22_X1  g431(.A1(new_n630_), .A2(new_n631_), .B1(new_n620_), .B2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT40), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(G1325gat));
  OAI21_X1  g434(.A(G15gat), .B1(new_n609_), .B2(new_n273_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT41), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n636_), .A2(new_n637_), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n273_), .A2(G15gat), .ZN(new_n640_));
  OAI22_X1  g439(.A1(new_n638_), .A2(new_n639_), .B1(new_n620_), .B2(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT99), .ZN(G1326gat));
  INV_X1    g441(.A(KEYINPUT42), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n627_), .A2(new_n432_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n643_), .B1(new_n644_), .B2(G22gat), .ZN(new_n645_));
  INV_X1    g444(.A(G22gat), .ZN(new_n646_));
  AOI211_X1 g445(.A(KEYINPUT42), .B(new_n646_), .C1(new_n627_), .C2(new_n432_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n432_), .A2(new_n646_), .ZN(new_n648_));
  OAI22_X1  g447(.A1(new_n645_), .A2(new_n647_), .B1(new_n620_), .B2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT100), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(G1327gat));
  NOR2_X1   g450(.A1(new_n615_), .A2(new_n519_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n653_), .A2(new_n563_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n619_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(G29gat), .B1(new_n656_), .B2(new_n342_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT101), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(KEYINPUT43), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n614_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n273_), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n403_), .A2(new_n466_), .A3(new_n406_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n663_), .B1(new_n460_), .B2(KEYINPUT94), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n662_), .B1(new_n664_), .B2(new_n465_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n661_), .B1(new_n665_), .B2(new_n442_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n658_), .A2(KEYINPUT43), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n660_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(KEYINPUT102), .A2(KEYINPUT43), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n669_), .B1(new_n665_), .B2(new_n442_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n467_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n460_), .A2(KEYINPUT94), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n273_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n441_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n439_), .A2(new_n440_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n343_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n673_), .A2(KEYINPUT102), .A3(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n670_), .A2(new_n661_), .A3(new_n677_), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n563_), .A2(new_n615_), .A3(new_n607_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n668_), .A2(new_n678_), .A3(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT44), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n682_), .A2(G29gat), .A3(new_n342_), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n668_), .A2(new_n678_), .A3(KEYINPUT44), .A4(new_n679_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n657_), .B1(new_n683_), .B2(new_n684_), .ZN(G1328gat));
  NOR2_X1   g484(.A1(KEYINPUT103), .A2(KEYINPUT46), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT104), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n407_), .A2(G36gat), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n656_), .A2(KEYINPUT45), .A3(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT45), .ZN(new_n691_));
  INV_X1    g490(.A(new_n689_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n691_), .B1(new_n655_), .B2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n690_), .A2(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n407_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(new_n684_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n694_), .B1(new_n696_), .B2(G36gat), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT103), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT46), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n688_), .B1(new_n697_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(G36gat), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n702_), .B1(new_n695_), .B2(new_n684_), .ZN(new_n703_));
  OAI221_X1 g502(.A(new_n687_), .B1(new_n698_), .B2(new_n699_), .C1(new_n703_), .C2(new_n694_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n701_), .A2(new_n704_), .ZN(G1329gat));
  NAND4_X1  g504(.A1(new_n682_), .A2(new_n684_), .A3(G43gat), .A4(new_n662_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n655_), .A2(new_n273_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n706_), .B1(G43gat), .B2(new_n707_), .ZN(new_n708_));
  XOR2_X1   g507(.A(KEYINPUT105), .B(KEYINPUT47), .Z(new_n709_));
  XNOR2_X1  g508(.A(new_n708_), .B(new_n709_), .ZN(G1330gat));
  AOI21_X1  g509(.A(G50gat), .B1(new_n656_), .B2(new_n432_), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n682_), .A2(G50gat), .A3(new_n432_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n711_), .B1(new_n712_), .B2(new_n684_), .ZN(G1331gat));
  NOR2_X1   g512(.A1(new_n585_), .A2(new_n606_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n563_), .A2(new_n714_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n521_), .A2(new_n715_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(KEYINPUT107), .B(G57gat), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n716_), .A2(new_n342_), .A3(new_n717_), .ZN(new_n718_));
  XOR2_X1   g517(.A(new_n718_), .B(KEYINPUT108), .Z(new_n719_));
  INV_X1    g518(.A(new_n563_), .ZN(new_n720_));
  OR4_X1    g519(.A1(new_n469_), .A2(new_n617_), .A3(new_n606_), .A4(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n341_), .B1(new_n721_), .B2(KEYINPUT106), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n722_), .B1(KEYINPUT106), .B2(new_n721_), .ZN(new_n723_));
  INV_X1    g522(.A(G57gat), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n719_), .B1(new_n723_), .B2(new_n724_), .ZN(G1332gat));
  NAND2_X1  g524(.A1(new_n521_), .A2(new_n715_), .ZN(new_n726_));
  OAI21_X1  g525(.A(G64gat), .B1(new_n726_), .B2(new_n407_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(KEYINPUT109), .B(KEYINPUT48), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n727_), .B(new_n728_), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n407_), .A2(G64gat), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n729_), .B1(new_n721_), .B2(new_n730_), .ZN(G1333gat));
  OAI21_X1  g530(.A(G71gat), .B1(new_n726_), .B2(new_n273_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT49), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n662_), .A2(new_n262_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n733_), .B1(new_n721_), .B2(new_n734_), .ZN(G1334gat));
  NAND2_X1  g534(.A1(new_n716_), .A2(new_n432_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n736_), .A2(G78gat), .A3(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n737_), .B1(new_n736_), .B2(G78gat), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n432_), .A2(new_n419_), .ZN(new_n740_));
  OAI22_X1  g539(.A1(new_n738_), .A2(new_n739_), .B1(new_n721_), .B2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT111), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n741_), .B(new_n742_), .ZN(G1335gat));
  NAND2_X1  g542(.A1(new_n668_), .A2(new_n678_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT112), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n563_), .A2(new_n585_), .A3(new_n607_), .ZN(new_n747_));
  OR2_X1    g546(.A1(new_n747_), .A2(KEYINPUT113), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(KEYINPUT113), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n668_), .A2(KEYINPUT112), .A3(new_n678_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n746_), .A2(new_n750_), .A3(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(G85gat), .B1(new_n752_), .B2(new_n341_), .ZN(new_n753_));
  NOR4_X1   g552(.A1(new_n469_), .A2(new_n606_), .A3(new_n720_), .A4(new_n653_), .ZN(new_n754_));
  INV_X1    g553(.A(G85gat), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n754_), .A2(new_n755_), .A3(new_n342_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n753_), .A2(new_n756_), .ZN(G1336gat));
  OAI21_X1  g556(.A(G92gat), .B1(new_n752_), .B2(new_n407_), .ZN(new_n758_));
  INV_X1    g557(.A(G92gat), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n754_), .A2(new_n759_), .A3(new_n628_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(G1337gat));
  OAI21_X1  g560(.A(G99gat), .B1(new_n752_), .B2(new_n273_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n754_), .A2(new_n662_), .A3(new_n476_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(KEYINPUT51), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT51), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n762_), .A2(new_n766_), .A3(new_n763_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n765_), .A2(new_n767_), .ZN(G1338gat));
  OAI21_X1  g567(.A(new_n667_), .B1(new_n469_), .B2(new_n614_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n433_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n678_), .A2(new_n659_), .A3(new_n769_), .A4(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT114), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n668_), .A2(new_n678_), .A3(KEYINPUT114), .A4(new_n770_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT115), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n421_), .B1(new_n775_), .B2(KEYINPUT52), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n773_), .A2(new_n774_), .A3(new_n776_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n775_), .A2(KEYINPUT52), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n778_), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n773_), .A2(new_n774_), .A3(new_n776_), .A4(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n754_), .A2(new_n421_), .A3(new_n432_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n779_), .A2(new_n781_), .A3(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT53), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n779_), .A2(new_n785_), .A3(new_n781_), .A4(new_n782_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(G1339gat));
  AOI211_X1 g586(.A(new_n341_), .B(new_n273_), .C1(new_n434_), .C2(new_n441_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT57), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n606_), .A2(new_n558_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n538_), .B1(new_n546_), .B2(new_n549_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n542_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n550_), .A2(new_n793_), .ZN(new_n794_));
  OAI211_X1 g593(.A(KEYINPUT55), .B(new_n545_), .C1(new_n546_), .C2(new_n549_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n792_), .A2(new_n794_), .A3(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(new_n555_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT116), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT56), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n790_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT116), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n801_), .B1(new_n796_), .B2(new_n555_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT56), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n589_), .A2(new_n590_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n586_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n586_), .B1(new_n587_), .B2(new_n595_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n602_), .B1(new_n594_), .B2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n805_), .A2(new_n807_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n603_), .A2(new_n808_), .ZN(new_n809_));
  AOI22_X1  g608(.A1(new_n800_), .A2(new_n803_), .B1(new_n559_), .B2(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n789_), .B1(new_n810_), .B2(new_n520_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n809_), .A2(new_n558_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n797_), .A2(KEYINPUT117), .A3(KEYINPUT56), .ZN(new_n813_));
  OR2_X1    g612(.A1(KEYINPUT117), .A2(KEYINPUT56), .ZN(new_n814_));
  NAND2_X1  g613(.A1(KEYINPUT117), .A2(KEYINPUT56), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n796_), .A2(new_n555_), .A3(new_n814_), .A4(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n812_), .A2(new_n813_), .A3(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT58), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n812_), .A2(new_n813_), .A3(KEYINPUT58), .A4(new_n816_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n819_), .A2(new_n661_), .A3(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n559_), .A2(new_n809_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n803_), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n606_), .B(new_n558_), .C1(new_n802_), .C2(KEYINPUT56), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n822_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n825_), .A2(KEYINPUT57), .A3(new_n519_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n811_), .A2(new_n821_), .A3(new_n826_), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n827_), .A2(new_n585_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n614_), .A2(new_n714_), .ZN(new_n829_));
  OR3_X1    g628(.A1(new_n829_), .A2(KEYINPUT54), .A3(new_n563_), .ZN(new_n830_));
  OAI21_X1  g629(.A(KEYINPUT54), .B1(new_n829_), .B2(new_n563_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n788_), .B1(new_n828_), .B2(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n208_), .B1(new_n834_), .B2(new_n607_), .ZN(new_n835_));
  OR2_X1    g634(.A1(new_n835_), .A2(KEYINPUT118), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(KEYINPUT118), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n834_), .A2(KEYINPUT59), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT59), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT119), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n827_), .A2(new_n840_), .A3(new_n585_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n832_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n840_), .B1(new_n827_), .B2(new_n585_), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n839_), .B(new_n788_), .C1(new_n842_), .C2(new_n843_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n838_), .A2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n606_), .A2(G113gat), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(KEYINPUT120), .ZN(new_n847_));
  AOI22_X1  g646(.A1(new_n836_), .A2(new_n837_), .B1(new_n845_), .B2(new_n847_), .ZN(G1340gat));
  INV_X1    g647(.A(new_n834_), .ZN(new_n849_));
  XOR2_X1   g648(.A(KEYINPUT121), .B(G120gat), .Z(new_n850_));
  OAI21_X1  g649(.A(new_n850_), .B1(new_n720_), .B2(KEYINPUT60), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n849_), .B(new_n851_), .C1(KEYINPUT60), .C2(new_n850_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n845_), .A2(new_n563_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n853_), .B2(new_n850_), .ZN(G1341gat));
  NOR2_X1   g653(.A1(new_n585_), .A2(new_n204_), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n838_), .B(new_n844_), .C1(KEYINPUT122), .C2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(G127gat), .B1(new_n856_), .B2(KEYINPUT122), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n856_), .A2(new_n615_), .A3(new_n849_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(G1342gat));
  NAND3_X1  g658(.A1(new_n849_), .A2(new_n202_), .A3(new_n520_), .ZN(new_n860_));
  AND2_X1   g659(.A1(new_n845_), .A2(new_n661_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(new_n861_), .B2(new_n202_), .ZN(G1343gat));
  NOR2_X1   g661(.A1(new_n828_), .A2(new_n833_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n863_), .A2(new_n662_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n628_), .A2(new_n341_), .A3(new_n433_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n867_), .A2(new_n287_), .A3(new_n606_), .ZN(new_n868_));
  OAI21_X1  g667(.A(G141gat), .B1(new_n866_), .B2(new_n607_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(G1344gat));
  XNOR2_X1  g669(.A(KEYINPUT123), .B(G148gat), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n867_), .A2(new_n563_), .A3(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n871_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n873_), .B1(new_n866_), .B2(new_n720_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n872_), .A2(new_n874_), .ZN(G1345gat));
  XNOR2_X1  g674(.A(KEYINPUT61), .B(G155gat), .ZN(new_n876_));
  OR3_X1    g675(.A1(new_n866_), .A2(new_n585_), .A3(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n866_), .B2(new_n585_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(G1346gat));
  OR3_X1    g678(.A1(new_n866_), .A2(G162gat), .A3(new_n519_), .ZN(new_n880_));
  OAI21_X1  g679(.A(G162gat), .B1(new_n866_), .B2(new_n614_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(G1347gat));
  INV_X1    g681(.A(KEYINPUT62), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n344_), .A2(new_n432_), .A3(new_n407_), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n606_), .B(new_n884_), .C1(new_n842_), .C2(new_n843_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT124), .ZN(new_n886_));
  AND3_X1   g685(.A1(new_n885_), .A2(new_n886_), .A3(G169gat), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n886_), .B1(new_n885_), .B2(G169gat), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n883_), .B1(new_n887_), .B2(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n885_), .A2(G169gat), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(KEYINPUT124), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n885_), .A2(new_n886_), .A3(G169gat), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n891_), .A2(KEYINPUT62), .A3(new_n892_), .ZN(new_n893_));
  OR2_X1    g692(.A1(new_n842_), .A2(new_n843_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n884_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n896_), .A2(new_n255_), .A3(new_n606_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n889_), .A2(new_n893_), .A3(new_n897_), .ZN(G1348gat));
  NOR2_X1   g697(.A1(new_n863_), .A2(new_n432_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n344_), .A2(new_n407_), .ZN(new_n900_));
  NAND4_X1  g699(.A1(new_n899_), .A2(G176gat), .A3(new_n563_), .A4(new_n900_), .ZN(new_n901_));
  OAI211_X1 g700(.A(new_n563_), .B(new_n884_), .C1(new_n842_), .C2(new_n843_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(new_n256_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n901_), .A2(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT125), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n901_), .A2(KEYINPUT125), .A3(new_n903_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(G1349gat));
  NAND3_X1  g707(.A1(new_n899_), .A2(new_n615_), .A3(new_n900_), .ZN(new_n909_));
  OR2_X1    g708(.A1(new_n909_), .A2(KEYINPUT126), .ZN(new_n910_));
  AOI21_X1  g709(.A(G183gat), .B1(new_n909_), .B2(KEYINPUT126), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n585_), .B1(new_n231_), .B2(new_n233_), .ZN(new_n912_));
  AOI22_X1  g711(.A1(new_n910_), .A2(new_n911_), .B1(new_n896_), .B2(new_n912_), .ZN(G1350gat));
  OAI21_X1  g712(.A(G190gat), .B1(new_n895_), .B2(new_n614_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n520_), .A2(new_n235_), .A3(new_n237_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n914_), .B1(new_n895_), .B2(new_n915_), .ZN(G1351gat));
  NOR2_X1   g715(.A1(new_n407_), .A2(new_n466_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n864_), .A2(new_n917_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  AOI21_X1  g718(.A(G197gat), .B1(new_n919_), .B2(new_n606_), .ZN(new_n920_));
  NOR3_X1   g719(.A1(new_n918_), .A2(new_n363_), .A3(new_n607_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n920_), .A2(new_n921_), .ZN(G1352gat));
  NAND3_X1  g721(.A1(new_n919_), .A2(new_n364_), .A3(new_n563_), .ZN(new_n923_));
  OAI21_X1  g722(.A(G204gat), .B1(new_n918_), .B2(new_n720_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(new_n924_), .ZN(G1353gat));
  NOR2_X1   g724(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n926_));
  INV_X1    g725(.A(new_n926_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n585_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n928_));
  XOR2_X1   g727(.A(new_n928_), .B(KEYINPUT127), .Z(new_n929_));
  INV_X1    g728(.A(new_n929_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n927_), .B1(new_n919_), .B2(new_n930_), .ZN(new_n931_));
  NOR3_X1   g730(.A1(new_n918_), .A2(new_n926_), .A3(new_n929_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n931_), .A2(new_n932_), .ZN(G1354gat));
  OR3_X1    g732(.A1(new_n918_), .A2(G218gat), .A3(new_n519_), .ZN(new_n934_));
  OAI21_X1  g733(.A(G218gat), .B1(new_n918_), .B2(new_n614_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n934_), .A2(new_n935_), .ZN(G1355gat));
endmodule


