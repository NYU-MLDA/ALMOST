//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 0 1 1 0 0 0 1 1 1 0 1 0 0 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 0 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n809_, new_n810_, new_n811_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n856_, new_n858_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n958_, new_n959_,
    new_n960_, new_n961_, new_n963_, new_n964_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n971_, new_n972_, new_n973_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n986_, new_n987_, new_n988_,
    new_n990_, new_n991_, new_n992_, new_n994_, new_n995_, new_n997_,
    new_n998_, new_n999_, new_n1000_, new_n1002_, new_n1003_, new_n1004_,
    new_n1005_, new_n1006_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_,
    new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1023_, new_n1024_;
  XNOR2_X1  g000(.A(G22gat), .B(G50gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(KEYINPUT89), .A2(KEYINPUT3), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT2), .ZN(new_n209_));
  INV_X1    g008(.A(G141gat), .ZN(new_n210_));
  INV_X1    g009(.A(G148gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n209_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n213_));
  OAI22_X1  g012(.A1(KEYINPUT89), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n208_), .A2(new_n212_), .A3(new_n213_), .A4(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT87), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT87), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(G155gat), .A3(G162gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  OR2_X1    g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221_));
  AND3_X1   g020(.A1(new_n215_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n220_), .A2(KEYINPUT1), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT88), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT1), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n217_), .A2(new_n219_), .A3(new_n225_), .ZN(new_n226_));
  AND2_X1   g025(.A1(new_n226_), .A2(new_n221_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n225_), .B1(new_n217_), .B2(new_n219_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT88), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n224_), .A2(new_n227_), .A3(new_n230_), .ZN(new_n231_));
  OR2_X1    g030(.A1(new_n206_), .A2(KEYINPUT86), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n206_), .A2(KEYINPUT86), .ZN(new_n233_));
  AOI22_X1  g032(.A1(new_n232_), .A2(new_n233_), .B1(G141gat), .B2(G148gat), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n222_), .B1(new_n231_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT29), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n205_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  OAI211_X1 g036(.A(new_n221_), .B(new_n226_), .C1(new_n228_), .C2(new_n229_), .ZN(new_n238_));
  AOI211_X1 g037(.A(KEYINPUT88), .B(new_n225_), .C1(new_n217_), .C2(new_n219_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n234_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n222_), .ZN(new_n241_));
  AND4_X1   g040(.A1(new_n236_), .A2(new_n240_), .A3(new_n241_), .A4(new_n205_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n203_), .B1(new_n237_), .B2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n240_), .A2(new_n241_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n204_), .B1(new_n244_), .B2(KEYINPUT29), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n235_), .A2(new_n236_), .A3(new_n205_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n245_), .A2(new_n202_), .A3(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT92), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n243_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT93), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n236_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n251_));
  AND2_X1   g050(.A1(G197gat), .A2(G204gat), .ZN(new_n252_));
  NOR2_X1   g051(.A1(G197gat), .A2(G204gat), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT91), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT21), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G211gat), .B(G218gat), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n254_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n254_), .A2(new_n256_), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n252_), .A2(new_n253_), .ZN(new_n259_));
  XOR2_X1   g058(.A(G211gat), .B(G218gat), .Z(new_n260_));
  AOI21_X1  g059(.A(new_n255_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n257_), .B1(new_n258_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(G228gat), .ZN(new_n263_));
  INV_X1    g062(.A(G233gat), .ZN(new_n264_));
  OAI22_X1  g063(.A1(new_n251_), .A2(new_n262_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G78gat), .B(G106gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n261_), .A2(new_n258_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n257_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n263_), .A2(new_n264_), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n269_), .B(new_n270_), .C1(new_n235_), .C2(new_n236_), .ZN(new_n271_));
  AND3_X1   g070(.A1(new_n265_), .A2(new_n266_), .A3(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n266_), .B1(new_n265_), .B2(new_n271_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n243_), .A2(new_n247_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(KEYINPUT92), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT93), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n243_), .A2(new_n247_), .A3(new_n248_), .A4(new_n277_), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n250_), .A2(new_n274_), .A3(new_n276_), .A4(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n250_), .A2(new_n278_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n274_), .A2(new_n276_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G183gat), .A2(G190gat), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT23), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(G169gat), .ZN(new_n289_));
  INV_X1    g088(.A(G176gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G169gat), .A2(G176gat), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n291_), .A2(KEYINPUT24), .A3(new_n292_), .ZN(new_n293_));
  OR3_X1    g092(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n294_));
  AND3_X1   g093(.A1(new_n288_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT82), .ZN(new_n296_));
  INV_X1    g095(.A(G183gat), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT81), .B1(new_n297_), .B2(KEYINPUT25), .ZN(new_n298_));
  INV_X1    g097(.A(G190gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT26), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT26), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(G190gat), .ZN(new_n302_));
  AND3_X1   g101(.A1(new_n298_), .A2(new_n300_), .A3(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT25), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(G183gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n297_), .A2(KEYINPUT25), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT81), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n296_), .B1(new_n303_), .B2(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n298_), .A2(new_n300_), .A3(new_n302_), .ZN(new_n311_));
  AOI21_X1  g110(.A(KEYINPUT81), .B1(new_n305_), .B2(new_n306_), .ZN(new_n312_));
  NOR3_X1   g111(.A1(new_n311_), .A2(new_n312_), .A3(KEYINPUT82), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n295_), .B1(new_n310_), .B2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n289_), .A2(KEYINPUT22), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT22), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(G169gat), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n315_), .A2(new_n317_), .A3(new_n290_), .ZN(new_n318_));
  AOI21_X1  g117(.A(KEYINPUT83), .B1(new_n318_), .B2(new_n292_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(G183gat), .A2(G190gat), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n287_), .A2(new_n320_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  AND3_X1   g121(.A1(new_n318_), .A2(KEYINPUT83), .A3(new_n292_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n314_), .A2(KEYINPUT30), .A3(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT30), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n288_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n303_), .A2(new_n309_), .A3(new_n296_), .ZN(new_n329_));
  OAI21_X1  g128(.A(KEYINPUT82), .B1(new_n311_), .B2(new_n312_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n328_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  NOR3_X1   g130(.A1(new_n323_), .A2(new_n319_), .A3(new_n321_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n327_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT84), .ZN(new_n334_));
  AND3_X1   g133(.A1(new_n326_), .A2(new_n333_), .A3(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n334_), .B1(new_n326_), .B2(new_n333_), .ZN(new_n336_));
  INV_X1    g135(.A(G227gat), .ZN(new_n337_));
  OAI22_X1  g136(.A1(new_n335_), .A2(new_n336_), .B1(new_n337_), .B2(new_n264_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G15gat), .B(G43gat), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NOR3_X1   g139(.A1(new_n331_), .A2(new_n332_), .A3(new_n327_), .ZN(new_n341_));
  AOI21_X1  g140(.A(KEYINPUT30), .B1(new_n314_), .B2(new_n325_), .ZN(new_n342_));
  OAI21_X1  g141(.A(KEYINPUT84), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n337_), .A2(new_n264_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n326_), .A2(new_n333_), .A3(new_n334_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n343_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  AND3_X1   g145(.A1(new_n338_), .A2(new_n340_), .A3(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n340_), .B1(new_n338_), .B2(new_n346_), .ZN(new_n348_));
  INV_X1    g147(.A(G127gat), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n349_), .A2(G134gat), .ZN(new_n350_));
  INV_X1    g149(.A(G134gat), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n351_), .A2(G127gat), .ZN(new_n352_));
  INV_X1    g151(.A(G113gat), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n353_), .A2(G120gat), .ZN(new_n354_));
  INV_X1    g153(.A(G120gat), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n355_), .A2(G113gat), .ZN(new_n356_));
  OAI22_X1  g155(.A1(new_n350_), .A2(new_n352_), .B1(new_n354_), .B2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G127gat), .B(G134gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G113gat), .B(G120gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n357_), .A2(new_n360_), .A3(KEYINPUT85), .ZN(new_n361_));
  OR3_X1    g160(.A1(new_n358_), .A2(new_n359_), .A3(KEYINPUT85), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT31), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G71gat), .B(G99gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NOR3_X1   g166(.A1(new_n347_), .A2(new_n348_), .A3(new_n367_), .ZN(new_n368_));
  AND3_X1   g167(.A1(new_n343_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n344_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n339_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n338_), .A2(new_n340_), .A3(new_n346_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n366_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  OAI211_X1 g172(.A(new_n279_), .B(new_n282_), .C1(new_n368_), .C2(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n371_), .A2(new_n366_), .A3(new_n372_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n367_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n376_));
  AND4_X1   g175(.A1(new_n276_), .A2(new_n250_), .A3(new_n274_), .A4(new_n278_), .ZN(new_n377_));
  AOI22_X1  g176(.A1(new_n250_), .A2(new_n278_), .B1(new_n274_), .B2(new_n276_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n375_), .B(new_n376_), .C1(new_n377_), .C2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n374_), .A2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(KEYINPUT100), .B(KEYINPUT27), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G8gat), .B(G36gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT18), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(G64gat), .ZN(new_n384_));
  INV_X1    g183(.A(G92gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT95), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n314_), .A2(new_n262_), .A3(new_n325_), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n285_), .B(new_n286_), .C1(G183gat), .C2(G190gat), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n389_), .A2(new_n318_), .A3(new_n292_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(KEYINPUT94), .ZN(new_n391_));
  INV_X1    g190(.A(new_n292_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT22), .B(G169gat), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n392_), .B1(new_n393_), .B2(new_n290_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT94), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n394_), .A2(new_n395_), .A3(new_n389_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n300_), .A2(new_n302_), .A3(new_n305_), .A4(new_n306_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n288_), .A2(new_n397_), .A3(new_n294_), .A4(new_n293_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n391_), .A2(new_n396_), .A3(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n269_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n388_), .A2(new_n400_), .A3(KEYINPUT20), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G226gat), .A2(G233gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(KEYINPUT19), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n269_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n262_), .A2(new_n396_), .A3(new_n398_), .A4(new_n391_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT20), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n403_), .A2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n405_), .A2(new_n406_), .A3(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT96), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT96), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n405_), .A2(new_n406_), .A3(new_n411_), .A4(new_n408_), .ZN(new_n412_));
  AOI22_X1  g211(.A1(new_n387_), .A2(new_n404_), .B1(new_n410_), .B2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n401_), .A2(KEYINPUT95), .A3(new_n403_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n386_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n404_), .A2(new_n387_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n410_), .A2(new_n412_), .ZN(new_n417_));
  AND4_X1   g216(.A1(new_n386_), .A2(new_n416_), .A3(new_n417_), .A4(new_n414_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n381_), .B1(new_n415_), .B2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G225gat), .A2(G233gat), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n244_), .A2(new_n363_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n357_), .A2(new_n360_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n235_), .A2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n422_), .A2(new_n424_), .A3(KEYINPUT4), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT97), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n361_), .A2(new_n362_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n427_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT4), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n426_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NOR4_X1   g229(.A1(new_n235_), .A2(KEYINPUT97), .A3(new_n427_), .A4(KEYINPUT4), .ZN(new_n431_));
  OAI211_X1 g230(.A(new_n421_), .B(new_n425_), .C1(new_n430_), .C2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(KEYINPUT98), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n244_), .A2(new_n429_), .A3(new_n363_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT97), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n428_), .A2(new_n426_), .A3(new_n429_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT98), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n437_), .A2(new_n438_), .A3(new_n421_), .A4(new_n425_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n422_), .A2(new_n424_), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT99), .B1(new_n440_), .B2(new_n421_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT99), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n422_), .A2(new_n424_), .A3(new_n442_), .A4(new_n420_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n441_), .A2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n433_), .A2(new_n439_), .A3(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G1gat), .B(G29gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(KEYINPUT0), .ZN(new_n447_));
  INV_X1    g246(.A(G57gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n447_), .B(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(G85gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n449_), .B(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n445_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n451_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n433_), .A2(new_n453_), .A3(new_n439_), .A4(new_n444_), .ZN(new_n454_));
  OR2_X1    g253(.A1(new_n401_), .A2(new_n403_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n262_), .A2(new_n390_), .A3(new_n398_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n405_), .A2(KEYINPUT20), .A3(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(new_n403_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n455_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n386_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n416_), .A2(new_n417_), .A3(new_n414_), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n461_), .B(KEYINPUT27), .C1(new_n460_), .C2(new_n462_), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n419_), .A2(new_n452_), .A3(new_n454_), .A4(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n380_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT33), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n454_), .A2(new_n467_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n415_), .A2(new_n418_), .ZN(new_n469_));
  AOI22_X1  g268(.A1(new_n432_), .A2(KEYINPUT98), .B1(new_n441_), .B2(new_n443_), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n470_), .A2(KEYINPUT33), .A3(new_n453_), .A4(new_n439_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n437_), .A2(new_n420_), .A3(new_n425_), .ZN(new_n472_));
  OAI211_X1 g271(.A(new_n472_), .B(new_n451_), .C1(new_n420_), .C2(new_n440_), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n468_), .A2(new_n469_), .A3(new_n471_), .A4(new_n473_), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n455_), .A2(new_n458_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n386_), .A2(KEYINPUT32), .ZN(new_n476_));
  MUX2_X1   g275(.A(new_n475_), .B(new_n462_), .S(new_n476_), .Z(new_n477_));
  INV_X1    g276(.A(new_n454_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n453_), .B1(new_n470_), .B2(new_n439_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n477_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n474_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n376_), .A2(new_n375_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n282_), .A2(new_n279_), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n481_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n466_), .A2(new_n485_), .ZN(new_n486_));
  XOR2_X1   g285(.A(G120gat), .B(G148gat), .Z(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(G204gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(KEYINPUT5), .B(G176gat), .ZN(new_n489_));
  XOR2_X1   g288(.A(new_n488_), .B(new_n489_), .Z(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT8), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n450_), .A2(new_n385_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(G85gat), .A2(G92gat), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(G99gat), .A2(G106gat), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT7), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G99gat), .A2(G106gat), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT6), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n495_), .B1(new_n498_), .B2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n496_), .B(KEYINPUT7), .ZN(new_n503_));
  OR2_X1    g302(.A1(KEYINPUT65), .A2(KEYINPUT6), .ZN(new_n504_));
  NAND2_X1  g303(.A1(KEYINPUT65), .A2(KEYINPUT6), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n499_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n504_), .A2(new_n499_), .A3(new_n505_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n503_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  NOR3_X1   g309(.A1(new_n493_), .A2(new_n492_), .A3(new_n494_), .ZN(new_n511_));
  AOI22_X1  g310(.A1(new_n492_), .A2(new_n502_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G71gat), .B(G78gat), .ZN(new_n513_));
  XOR2_X1   g312(.A(G57gat), .B(G64gat), .Z(new_n514_));
  INV_X1    g313(.A(KEYINPUT11), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n513_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G57gat), .B(G64gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(KEYINPUT11), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n517_), .A2(new_n513_), .A3(KEYINPUT11), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n493_), .A2(KEYINPUT9), .ZN(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT64), .B(G85gat), .ZN(new_n523_));
  AND2_X1   g322(.A1(new_n523_), .A2(G92gat), .ZN(new_n524_));
  OAI21_X1  g323(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n522_), .B1(new_n524_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(G106gat), .ZN(new_n528_));
  XOR2_X1   g327(.A(KEYINPUT10), .B(G99gat), .Z(new_n529_));
  AOI21_X1  g328(.A(new_n501_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n527_), .A2(new_n530_), .ZN(new_n531_));
  AND3_X1   g330(.A1(new_n512_), .A2(new_n521_), .A3(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n519_), .A2(KEYINPUT68), .A3(new_n520_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(KEYINPUT68), .B1(new_n519_), .B2(new_n520_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT12), .ZN(new_n536_));
  NOR3_X1   g335(.A1(new_n534_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n502_), .A2(new_n492_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n510_), .A2(new_n511_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n531_), .A2(new_n538_), .A3(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n532_), .B1(new_n537_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G230gat), .A2(G233gat), .ZN(new_n542_));
  INV_X1    g341(.A(new_n521_), .ZN(new_n543_));
  AOI21_X1  g342(.A(KEYINPUT12), .B1(new_n540_), .B2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(KEYINPUT69), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT69), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n521_), .B1(new_n512_), .B2(new_n531_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n546_), .B1(new_n547_), .B2(KEYINPUT12), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n541_), .A2(new_n542_), .A3(new_n545_), .A4(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n512_), .A2(new_n521_), .A3(new_n531_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n550_), .B1(new_n547_), .B2(KEYINPUT66), .ZN(new_n551_));
  OR3_X1    g350(.A1(new_n540_), .A2(KEYINPUT66), .A3(new_n543_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n542_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n549_), .B1(KEYINPUT67), .B2(new_n553_), .ZN(new_n554_));
  AND2_X1   g353(.A1(new_n553_), .A2(KEYINPUT67), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n491_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT67), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n551_), .A2(new_n552_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n557_), .B1(new_n558_), .B2(new_n542_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n553_), .A2(KEYINPUT67), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n559_), .A2(new_n560_), .A3(new_n549_), .A4(new_n490_), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n556_), .A2(KEYINPUT13), .A3(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(KEYINPUT13), .B1(new_n556_), .B2(new_n561_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G43gat), .B(G50gat), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(G36gat), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(G29gat), .ZN(new_n567_));
  INV_X1    g366(.A(G29gat), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(G36gat), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT70), .ZN(new_n570_));
  AND3_X1   g369(.A1(new_n567_), .A2(new_n569_), .A3(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n570_), .B1(new_n567_), .B2(new_n569_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n565_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n567_), .A2(new_n569_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(KEYINPUT70), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n567_), .A2(new_n569_), .A3(new_n570_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n575_), .A2(new_n564_), .A3(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n573_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT15), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G15gat), .B(G22gat), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G1gat), .A2(G8gat), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(KEYINPUT14), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(G1gat), .ZN(new_n585_));
  INV_X1    g384(.A(G8gat), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT75), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n587_), .A2(new_n588_), .A3(new_n582_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n588_), .B1(new_n587_), .B2(new_n582_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n584_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G1gat), .B(G8gat), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(KEYINPUT75), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n594_), .A2(new_n583_), .A3(new_n581_), .A4(new_n589_), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n592_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n573_), .A2(new_n577_), .A3(KEYINPUT15), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n580_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(G229gat), .A2(G233gat), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n592_), .A2(new_n595_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(new_n578_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n598_), .A2(new_n599_), .A3(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT79), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT79), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n598_), .A2(new_n604_), .A3(new_n599_), .A4(new_n601_), .ZN(new_n605_));
  OR3_X1    g404(.A1(new_n600_), .A2(new_n578_), .A3(KEYINPUT78), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n592_), .A2(new_n595_), .A3(new_n573_), .A4(new_n577_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n601_), .A2(KEYINPUT78), .A3(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n599_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n606_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n603_), .A2(new_n605_), .A3(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G113gat), .B(G141gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(G169gat), .ZN(new_n613_));
  INV_X1    g412(.A(G197gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n611_), .A2(new_n616_), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n603_), .A2(new_n605_), .A3(new_n610_), .A4(new_n615_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT80), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n617_), .A2(KEYINPUT80), .A3(new_n618_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NOR3_X1   g423(.A1(new_n562_), .A2(new_n563_), .A3(new_n624_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n486_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n578_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n540_), .A2(new_n627_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n580_), .A2(new_n597_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n628_), .B1(new_n540_), .B2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(G232gat), .A2(G233gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT34), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(KEYINPUT35), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n540_), .A2(new_n597_), .A3(new_n580_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT71), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n633_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n632_), .A2(KEYINPUT35), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n630_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(G190gat), .B(G218gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(G134gat), .B(G162gat), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n639_), .B(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n641_), .A2(KEYINPUT36), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n634_), .B1(new_n540_), .B2(new_n627_), .ZN(new_n644_));
  AOI21_X1  g443(.A(KEYINPUT71), .B1(new_n629_), .B2(new_n540_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n644_), .B1(new_n645_), .B2(new_n633_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n641_), .A2(KEYINPUT36), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n638_), .A2(new_n643_), .A3(new_n646_), .A4(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT73), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT74), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n648_), .A2(new_n649_), .A3(new_n650_), .A4(KEYINPUT37), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n651_), .B1(new_n649_), .B2(new_n648_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n638_), .A2(new_n646_), .ZN(new_n653_));
  AOI21_X1  g452(.A(KEYINPUT72), .B1(new_n653_), .B2(new_n642_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT72), .ZN(new_n655_));
  AOI211_X1 g454(.A(new_n655_), .B(new_n643_), .C1(new_n638_), .C2(new_n646_), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n654_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n652_), .A2(new_n657_), .ZN(new_n658_));
  OAI211_X1 g457(.A(new_n650_), .B(new_n648_), .C1(new_n654_), .C2(new_n656_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n658_), .B1(new_n660_), .B2(KEYINPUT37), .ZN(new_n661_));
  XNOR2_X1  g460(.A(G127gat), .B(G155gat), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT16), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n662_), .B(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(G183gat), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n662_), .B(KEYINPUT16), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(new_n297_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n665_), .A2(new_n667_), .A3(G211gat), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(G211gat), .B1(new_n665_), .B2(new_n667_), .ZN(new_n670_));
  OAI21_X1  g469(.A(KEYINPUT17), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n596_), .A2(G231gat), .A3(G233gat), .ZN(new_n672_));
  INV_X1    g471(.A(G231gat), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n600_), .B1(new_n673_), .B2(new_n264_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n672_), .A2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(new_n543_), .ZN(new_n676_));
  OR3_X1    g475(.A1(new_n669_), .A2(KEYINPUT17), .A3(new_n670_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n672_), .A2(new_n674_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(new_n521_), .ZN(new_n679_));
  AND4_X1   g478(.A1(new_n671_), .A2(new_n676_), .A3(new_n677_), .A4(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT76), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n681_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT68), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n521_), .A2(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n684_), .A2(KEYINPUT76), .A3(new_n533_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n675_), .A2(new_n682_), .A3(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT77), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n671_), .A2(new_n687_), .ZN(new_n688_));
  OAI211_X1 g487(.A(KEYINPUT77), .B(KEYINPUT17), .C1(new_n669_), .C2(new_n670_), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n686_), .A2(new_n688_), .A3(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n682_), .A2(new_n685_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(new_n678_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n680_), .B1(new_n690_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n661_), .A2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n626_), .A2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT101), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n626_), .A2(KEYINPUT101), .A3(new_n695_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n452_), .A2(new_n454_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n700_), .A2(new_n585_), .A3(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT38), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n648_), .B1(new_n654_), .B2(new_n656_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT102), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  OAI211_X1 g506(.A(KEYINPUT102), .B(new_n648_), .C1(new_n654_), .C2(new_n656_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n709_), .A2(new_n694_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n486_), .A2(new_n710_), .A3(new_n625_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n701_), .ZN(new_n712_));
  OAI21_X1  g511(.A(G1gat), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT103), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n702_), .A2(new_n714_), .A3(new_n703_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n716_));
  OAI211_X1 g515(.A(new_n704_), .B(new_n713_), .C1(new_n715_), .C2(new_n716_), .ZN(G1324gat));
  NAND2_X1  g516(.A1(new_n419_), .A2(new_n463_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(G8gat), .B1(new_n711_), .B2(new_n719_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT39), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n698_), .A2(new_n586_), .A3(new_n718_), .A4(new_n699_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(KEYINPUT104), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT104), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n721_), .A2(new_n725_), .A3(new_n722_), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n724_), .A2(KEYINPUT40), .A3(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(KEYINPUT40), .B1(new_n724_), .B2(new_n726_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1325gat));
  INV_X1    g528(.A(G15gat), .ZN(new_n730_));
  INV_X1    g529(.A(new_n482_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n700_), .A2(new_n730_), .A3(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT105), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n733_), .ZN(new_n735_));
  OAI21_X1  g534(.A(G15gat), .B1(new_n711_), .B2(new_n482_), .ZN(new_n736_));
  XOR2_X1   g535(.A(new_n736_), .B(KEYINPUT41), .Z(new_n737_));
  NAND3_X1  g536(.A1(new_n734_), .A2(new_n735_), .A3(new_n737_), .ZN(G1326gat));
  INV_X1    g537(.A(G22gat), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n483_), .B(KEYINPUT106), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n700_), .A2(new_n739_), .A3(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n740_), .ZN(new_n742_));
  OAI21_X1  g541(.A(G22gat), .B1(new_n711_), .B2(new_n742_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(KEYINPUT107), .B(KEYINPUT42), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n743_), .B(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n741_), .A2(new_n745_), .ZN(G1327gat));
  NAND2_X1  g545(.A1(new_n709_), .A2(new_n694_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT110), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n747_), .B(new_n748_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n749_), .A2(new_n626_), .ZN(new_n750_));
  AOI21_X1  g549(.A(G29gat), .B1(new_n750_), .B2(new_n701_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT43), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT37), .ZN(new_n754_));
  AOI22_X1  g553(.A1(new_n657_), .A2(new_n652_), .B1(new_n659_), .B2(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n755_), .B1(new_n466_), .B2(new_n485_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n753_), .B1(new_n756_), .B2(KEYINPUT108), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n482_), .A2(new_n483_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n758_), .B1(new_n480_), .B2(new_n474_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n464_), .B1(new_n374_), .B2(new_n379_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n661_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT108), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n761_), .A2(new_n762_), .A3(KEYINPUT43), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n757_), .A2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n625_), .A2(new_n694_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  AND4_X1   g565(.A1(new_n752_), .A2(new_n764_), .A3(KEYINPUT44), .A4(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n765_), .B1(new_n757_), .B2(new_n763_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n752_), .B1(new_n768_), .B2(KEYINPUT44), .ZN(new_n769_));
  OR2_X1    g568(.A1(new_n767_), .A2(new_n769_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n768_), .A2(KEYINPUT44), .ZN(new_n771_));
  NOR3_X1   g570(.A1(new_n771_), .A2(new_n568_), .A3(new_n712_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n751_), .B1(new_n770_), .B2(new_n772_), .ZN(G1328gat));
  INV_X1    g572(.A(KEYINPUT111), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT46), .ZN(new_n775_));
  AOI21_X1  g574(.A(KEYINPUT112), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n756_), .A2(KEYINPUT108), .A3(new_n753_), .ZN(new_n778_));
  AOI21_X1  g577(.A(KEYINPUT43), .B1(new_n761_), .B2(new_n762_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n766_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT44), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n719_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n782_), .B1(new_n767_), .B2(new_n769_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(G36gat), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n719_), .A2(G36gat), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n749_), .A2(new_n626_), .A3(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT45), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT45), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n749_), .A2(new_n626_), .A3(new_n788_), .A4(new_n785_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n775_), .A2(KEYINPUT112), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n777_), .B1(new_n784_), .B2(new_n793_), .ZN(new_n794_));
  AOI211_X1 g593(.A(new_n776_), .B(new_n792_), .C1(new_n783_), .C2(G36gat), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n794_), .A2(new_n795_), .ZN(G1329gat));
  INV_X1    g595(.A(new_n771_), .ZN(new_n797_));
  INV_X1    g596(.A(G43gat), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n482_), .A2(new_n798_), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n797_), .B(new_n799_), .C1(new_n767_), .C2(new_n769_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n749_), .A2(new_n626_), .A3(new_n731_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(new_n798_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(KEYINPUT113), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n800_), .A2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(KEYINPUT47), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT47), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n800_), .A2(new_n806_), .A3(new_n803_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n805_), .A2(new_n807_), .ZN(G1330gat));
  AOI21_X1  g607(.A(G50gat), .B1(new_n750_), .B2(new_n740_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n483_), .ZN(new_n810_));
  AND3_X1   g609(.A1(new_n797_), .A2(G50gat), .A3(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n809_), .B1(new_n811_), .B2(new_n770_), .ZN(G1331gat));
  NOR2_X1   g611(.A1(new_n562_), .A2(new_n563_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n813_), .A2(new_n623_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n486_), .A2(new_n710_), .A3(new_n814_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n815_), .B(KEYINPUT114), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(G57gat), .B1(new_n817_), .B2(new_n712_), .ZN(new_n818_));
  AND3_X1   g617(.A1(new_n695_), .A2(new_n486_), .A3(new_n814_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n819_), .A2(new_n448_), .A3(new_n701_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n820_), .ZN(G1332gat));
  INV_X1    g620(.A(G64gat), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n819_), .A2(new_n822_), .A3(new_n718_), .ZN(new_n823_));
  OAI21_X1  g622(.A(G64gat), .B1(new_n817_), .B2(new_n719_), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n824_), .A2(KEYINPUT48), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n824_), .A2(KEYINPUT48), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n823_), .B1(new_n825_), .B2(new_n826_), .ZN(G1333gat));
  INV_X1    g626(.A(G71gat), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n819_), .A2(new_n828_), .A3(new_n731_), .ZN(new_n829_));
  OAI21_X1  g628(.A(G71gat), .B1(new_n817_), .B2(new_n482_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n830_), .A2(KEYINPUT49), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n830_), .A2(KEYINPUT49), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n829_), .B1(new_n831_), .B2(new_n832_), .ZN(G1334gat));
  INV_X1    g632(.A(G78gat), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n819_), .A2(new_n834_), .A3(new_n740_), .ZN(new_n835_));
  OAI21_X1  g634(.A(G78gat), .B1(new_n817_), .B2(new_n742_), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n836_), .A2(KEYINPUT50), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n836_), .A2(KEYINPUT50), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n835_), .B1(new_n837_), .B2(new_n838_), .ZN(G1335gat));
  AND3_X1   g638(.A1(new_n749_), .A2(new_n486_), .A3(new_n814_), .ZN(new_n840_));
  AOI21_X1  g639(.A(G85gat), .B1(new_n840_), .B2(new_n701_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n764_), .A2(KEYINPUT115), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n814_), .A2(new_n694_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT115), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n757_), .A2(new_n845_), .A3(new_n763_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n842_), .A2(new_n844_), .A3(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n701_), .A2(new_n523_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n841_), .B1(new_n848_), .B2(new_n849_), .ZN(G1336gat));
  OAI21_X1  g649(.A(G92gat), .B1(new_n847_), .B2(new_n719_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n840_), .A2(new_n385_), .A3(new_n718_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(G1337gat));
  OAI21_X1  g652(.A(G99gat), .B1(new_n847_), .B2(new_n482_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n840_), .A2(new_n529_), .A3(new_n731_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g656(.A1(new_n840_), .A2(new_n528_), .A3(new_n810_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT52), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n843_), .A2(new_n483_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n764_), .A2(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n859_), .B1(new_n861_), .B2(G106gat), .ZN(new_n862_));
  AOI211_X1 g661(.A(KEYINPUT52), .B(new_n528_), .C1(new_n764_), .C2(new_n860_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n858_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g664(.A(new_n379_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n712_), .A2(new_n718_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n556_), .A2(new_n561_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT13), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n621_), .A2(new_n693_), .A3(new_n622_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT116), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n556_), .A2(KEYINPUT13), .A3(new_n561_), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n621_), .A2(new_n693_), .A3(KEYINPUT116), .A4(new_n622_), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n870_), .A2(new_n873_), .A3(new_n874_), .A4(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(KEYINPUT117), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT117), .ZN(new_n878_));
  NAND4_X1  g677(.A1(new_n813_), .A2(new_n878_), .A3(new_n875_), .A4(new_n873_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n755_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT118), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT54), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n881_), .A2(new_n882_), .A3(new_n883_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n880_), .A2(KEYINPUT118), .A3(new_n755_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(KEYINPUT54), .ZN(new_n886_));
  AOI21_X1  g685(.A(KEYINPUT118), .B1(new_n880_), .B2(new_n755_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n884_), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n540_), .A2(KEYINPUT12), .A3(new_n684_), .A4(new_n533_), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n550_), .B(new_n889_), .C1(new_n544_), .C2(KEYINPUT69), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n547_), .A2(new_n546_), .A3(KEYINPUT12), .ZN(new_n891_));
  INV_X1    g690(.A(new_n542_), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n890_), .A2(new_n891_), .A3(new_n892_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n890_), .B2(new_n891_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n893_), .B1(KEYINPUT55), .B2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT55), .ZN(new_n896_));
  NOR4_X1   g695(.A1(new_n890_), .A2(new_n891_), .A3(new_n896_), .A4(new_n892_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n491_), .B1(new_n895_), .B2(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(KEYINPUT56), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT56), .ZN(new_n900_));
  OAI211_X1 g699(.A(new_n900_), .B(new_n491_), .C1(new_n895_), .C2(new_n897_), .ZN(new_n901_));
  NAND4_X1  g700(.A1(new_n899_), .A2(new_n623_), .A3(new_n561_), .A4(new_n901_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n606_), .A2(new_n608_), .A3(new_n599_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n598_), .A2(new_n609_), .A3(new_n601_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n903_), .A2(new_n616_), .A3(new_n904_), .ZN(new_n905_));
  AND2_X1   g704(.A1(new_n618_), .A2(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n868_), .A2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n902_), .A2(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n709_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT57), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n912_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(KEYINPUT119), .A2(KEYINPUT58), .ZN(new_n914_));
  NAND4_X1  g713(.A1(new_n899_), .A2(new_n561_), .A3(new_n906_), .A4(new_n901_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n755_), .B1(new_n914_), .B2(new_n915_), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n554_), .A2(new_n555_), .A3(new_n491_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n917_), .B1(new_n898_), .B2(KEYINPUT56), .ZN(new_n918_));
  INV_X1    g717(.A(new_n914_), .ZN(new_n919_));
  NAND4_X1  g718(.A1(new_n918_), .A2(new_n906_), .A3(new_n901_), .A4(new_n919_), .ZN(new_n920_));
  AOI22_X1  g719(.A1(new_n910_), .A2(new_n911_), .B1(new_n916_), .B2(new_n920_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n693_), .B1(new_n913_), .B2(new_n921_), .ZN(new_n922_));
  OAI211_X1 g721(.A(new_n866_), .B(new_n867_), .C1(new_n888_), .C2(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(KEYINPUT59), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n915_), .A2(new_n914_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n925_), .A2(new_n661_), .A3(new_n920_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n709_), .B1(new_n902_), .B2(new_n907_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n926_), .B1(KEYINPUT57), .B2(new_n927_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n694_), .B1(new_n928_), .B2(new_n912_), .ZN(new_n929_));
  OAI211_X1 g728(.A(new_n929_), .B(new_n884_), .C1(new_n887_), .C2(new_n886_), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT59), .ZN(new_n931_));
  NAND4_X1  g730(.A1(new_n930_), .A2(new_n931_), .A3(new_n866_), .A4(new_n867_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n924_), .A2(new_n623_), .A3(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(G113gat), .ZN(new_n934_));
  AND2_X1   g733(.A1(new_n930_), .A2(new_n867_), .ZN(new_n935_));
  NAND4_X1  g734(.A1(new_n935_), .A2(new_n353_), .A3(new_n866_), .A4(new_n623_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n934_), .A2(new_n936_), .ZN(G1340gat));
  INV_X1    g736(.A(new_n813_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n924_), .A2(new_n938_), .A3(new_n932_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(KEYINPUT120), .B(G120gat), .ZN(new_n940_));
  INV_X1    g739(.A(new_n940_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n939_), .A2(new_n941_), .ZN(new_n942_));
  OR2_X1    g741(.A1(new_n940_), .A2(KEYINPUT60), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n940_), .B1(new_n813_), .B2(KEYINPUT60), .ZN(new_n944_));
  NAND4_X1  g743(.A1(new_n935_), .A2(new_n866_), .A3(new_n943_), .A4(new_n944_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n942_), .A2(new_n945_), .ZN(G1341gat));
  XOR2_X1   g745(.A(KEYINPUT121), .B(G127gat), .Z(new_n947_));
  NAND2_X1  g746(.A1(new_n693_), .A2(new_n947_), .ZN(new_n948_));
  XOR2_X1   g747(.A(new_n948_), .B(KEYINPUT122), .Z(new_n949_));
  NAND3_X1  g748(.A1(new_n924_), .A2(new_n932_), .A3(new_n949_), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n349_), .B1(new_n923_), .B2(new_n694_), .ZN(new_n951_));
  AND2_X1   g750(.A1(new_n950_), .A2(new_n951_), .ZN(G1342gat));
  NAND2_X1  g751(.A1(new_n661_), .A2(G134gat), .ZN(new_n953_));
  XNOR2_X1  g752(.A(new_n953_), .B(KEYINPUT123), .ZN(new_n954_));
  NAND3_X1  g753(.A1(new_n924_), .A2(new_n932_), .A3(new_n954_), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n351_), .B1(new_n923_), .B2(new_n909_), .ZN(new_n956_));
  AND2_X1   g755(.A1(new_n955_), .A2(new_n956_), .ZN(G1343gat));
  INV_X1    g756(.A(new_n374_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n935_), .A2(new_n958_), .ZN(new_n959_));
  OAI21_X1  g758(.A(G141gat), .B1(new_n959_), .B2(new_n624_), .ZN(new_n960_));
  NAND4_X1  g759(.A1(new_n935_), .A2(new_n210_), .A3(new_n958_), .A4(new_n623_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n960_), .A2(new_n961_), .ZN(G1344gat));
  OAI21_X1  g761(.A(G148gat), .B1(new_n959_), .B2(new_n813_), .ZN(new_n963_));
  NAND4_X1  g762(.A1(new_n935_), .A2(new_n211_), .A3(new_n958_), .A4(new_n938_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n963_), .A2(new_n964_), .ZN(G1345gat));
  XNOR2_X1  g764(.A(KEYINPUT61), .B(G155gat), .ZN(new_n966_));
  OAI21_X1  g765(.A(new_n966_), .B1(new_n959_), .B2(new_n694_), .ZN(new_n967_));
  INV_X1    g766(.A(new_n966_), .ZN(new_n968_));
  NAND4_X1  g767(.A1(new_n935_), .A2(new_n693_), .A3(new_n958_), .A4(new_n968_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n967_), .A2(new_n969_), .ZN(G1346gat));
  OAI21_X1  g769(.A(G162gat), .B1(new_n959_), .B2(new_n755_), .ZN(new_n971_));
  NOR2_X1   g770(.A1(new_n909_), .A2(G162gat), .ZN(new_n972_));
  NAND3_X1  g771(.A1(new_n935_), .A2(new_n958_), .A3(new_n972_), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n971_), .A2(new_n973_), .ZN(G1347gat));
  NOR2_X1   g773(.A1(new_n719_), .A2(new_n701_), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n975_), .A2(new_n731_), .ZN(new_n976_));
  NOR2_X1   g775(.A1(new_n976_), .A2(new_n740_), .ZN(new_n977_));
  NAND3_X1  g776(.A1(new_n930_), .A2(new_n623_), .A3(new_n977_), .ZN(new_n978_));
  NAND2_X1  g777(.A1(new_n978_), .A2(G169gat), .ZN(new_n979_));
  INV_X1    g778(.A(KEYINPUT62), .ZN(new_n980_));
  NAND2_X1  g779(.A1(new_n979_), .A2(new_n980_), .ZN(new_n981_));
  AND2_X1   g780(.A1(new_n930_), .A2(new_n977_), .ZN(new_n982_));
  NAND3_X1  g781(.A1(new_n982_), .A2(new_n393_), .A3(new_n623_), .ZN(new_n983_));
  NAND3_X1  g782(.A1(new_n978_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n984_));
  NAND3_X1  g783(.A1(new_n981_), .A2(new_n983_), .A3(new_n984_), .ZN(G1348gat));
  AOI21_X1  g784(.A(G176gat), .B1(new_n982_), .B2(new_n938_), .ZN(new_n986_));
  AND2_X1   g785(.A1(new_n930_), .A2(new_n483_), .ZN(new_n987_));
  NOR3_X1   g786(.A1(new_n976_), .A2(new_n290_), .A3(new_n813_), .ZN(new_n988_));
  AOI21_X1  g787(.A(new_n986_), .B1(new_n987_), .B2(new_n988_), .ZN(G1349gat));
  NAND4_X1  g788(.A1(new_n987_), .A2(new_n693_), .A3(new_n731_), .A4(new_n975_), .ZN(new_n990_));
  NAND2_X1  g789(.A1(new_n693_), .A2(new_n307_), .ZN(new_n991_));
  INV_X1    g790(.A(new_n991_), .ZN(new_n992_));
  AOI22_X1  g791(.A1(new_n990_), .A2(new_n297_), .B1(new_n982_), .B2(new_n992_), .ZN(G1350gat));
  NAND4_X1  g792(.A1(new_n982_), .A2(new_n300_), .A3(new_n302_), .A4(new_n709_), .ZN(new_n994_));
  AND2_X1   g793(.A1(new_n982_), .A2(new_n661_), .ZN(new_n995_));
  OAI21_X1  g794(.A(new_n994_), .B1(new_n995_), .B2(new_n299_), .ZN(G1351gat));
  NAND2_X1  g795(.A1(new_n975_), .A2(new_n958_), .ZN(new_n997_));
  INV_X1    g796(.A(new_n997_), .ZN(new_n998_));
  NAND2_X1  g797(.A1(new_n930_), .A2(new_n998_), .ZN(new_n999_));
  NOR2_X1   g798(.A1(new_n999_), .A2(new_n624_), .ZN(new_n1000_));
  XNOR2_X1  g799(.A(new_n1000_), .B(new_n614_), .ZN(G1352gat));
  NOR2_X1   g800(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n1002_));
  AND2_X1   g801(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n1003_));
  OAI22_X1  g802(.A1(new_n999_), .A2(new_n813_), .B1(new_n1002_), .B2(new_n1003_), .ZN(new_n1004_));
  AND2_X1   g803(.A1(new_n930_), .A2(new_n998_), .ZN(new_n1005_));
  NAND2_X1  g804(.A1(new_n1005_), .A2(new_n938_), .ZN(new_n1006_));
  OAI21_X1  g805(.A(new_n1004_), .B1(new_n1006_), .B2(new_n1003_), .ZN(G1353gat));
  NAND2_X1  g806(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1008_));
  NAND2_X1  g807(.A1(new_n693_), .A2(new_n1008_), .ZN(new_n1009_));
  INV_X1    g808(.A(new_n1009_), .ZN(new_n1010_));
  NAND3_X1  g809(.A1(new_n930_), .A2(new_n998_), .A3(new_n1010_), .ZN(new_n1011_));
  NOR2_X1   g810(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1012_));
  XNOR2_X1  g811(.A(new_n1012_), .B(KEYINPUT125), .ZN(new_n1013_));
  NAND2_X1  g812(.A1(new_n1011_), .A2(new_n1013_), .ZN(new_n1014_));
  INV_X1    g813(.A(KEYINPUT127), .ZN(new_n1015_));
  NAND2_X1  g814(.A1(new_n1014_), .A2(new_n1015_), .ZN(new_n1016_));
  NAND3_X1  g815(.A1(new_n1011_), .A2(KEYINPUT127), .A3(new_n1013_), .ZN(new_n1017_));
  INV_X1    g816(.A(KEYINPUT126), .ZN(new_n1018_));
  INV_X1    g817(.A(new_n1013_), .ZN(new_n1019_));
  NAND4_X1  g818(.A1(new_n1005_), .A2(new_n1018_), .A3(new_n1019_), .A4(new_n1010_), .ZN(new_n1020_));
  OAI21_X1  g819(.A(KEYINPUT126), .B1(new_n1011_), .B2(new_n1013_), .ZN(new_n1021_));
  AOI22_X1  g820(.A1(new_n1016_), .A2(new_n1017_), .B1(new_n1020_), .B2(new_n1021_), .ZN(G1354gat));
  OAI21_X1  g821(.A(G218gat), .B1(new_n999_), .B2(new_n755_), .ZN(new_n1023_));
  OR2_X1    g822(.A1(new_n909_), .A2(G218gat), .ZN(new_n1024_));
  OAI21_X1  g823(.A(new_n1023_), .B1(new_n999_), .B2(new_n1024_), .ZN(G1355gat));
endmodule


