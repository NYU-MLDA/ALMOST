//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 1 1 1 1 0 0 0 0 1 1 1 1 0 1 0 1 0 1 0 1 1 1 0 0 0 1 0 1 0 1 0 0 0 0 0 1 1 0 1 0 0 0 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n704_, new_n705_, new_n706_, new_n707_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n807_, new_n808_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_, new_n910_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n917_, new_n918_,
    new_n920_, new_n921_, new_n922_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n958_, new_n959_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n966_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n975_, new_n976_,
    new_n977_, new_n978_, new_n979_, new_n980_, new_n981_, new_n982_,
    new_n983_, new_n984_;
  INV_X1    g000(.A(KEYINPUT103), .ZN(new_n202_));
  NOR2_X1   g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT1), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(new_n206_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT1), .ZN(new_n209_));
  INV_X1    g008(.A(G141gat), .ZN(new_n210_));
  INV_X1    g009(.A(G148gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G141gat), .A2(G148gat), .ZN(new_n213_));
  NAND4_X1  g012(.A1(new_n207_), .A2(new_n209_), .A3(new_n212_), .A4(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n210_), .A2(new_n211_), .A3(KEYINPUT3), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT3), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n216_), .B1(G141gat), .B2(G148gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  AND3_X1   g017(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n219_));
  AOI21_X1  g018(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  AND2_X1   g020(.A1(new_n218_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT87), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n204_), .A2(new_n223_), .A3(new_n206_), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT87), .B1(new_n208_), .B2(new_n203_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n214_), .B1(new_n222_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT88), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n218_), .A2(new_n221_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n230_), .A2(new_n225_), .A3(new_n224_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n231_), .A2(KEYINPUT88), .A3(new_n214_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G127gat), .B(G134gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G113gat), .B(G120gat), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n234_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(KEYINPUT86), .A3(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT86), .ZN(new_n238_));
  AND2_X1   g037(.A1(new_n233_), .A2(new_n234_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n233_), .A2(new_n234_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n238_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n237_), .A2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n229_), .A2(new_n232_), .A3(new_n242_), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n231_), .B(new_n214_), .C1(new_n239_), .C2(new_n240_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n243_), .A2(KEYINPUT4), .A3(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT101), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n243_), .A2(new_n244_), .A3(KEYINPUT101), .A4(KEYINPUT4), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(KEYINPUT102), .B(KEYINPUT4), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n229_), .A2(new_n242_), .A3(new_n232_), .A4(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G225gat), .A2(G233gat), .ZN(new_n252_));
  AND2_X1   g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n249_), .A2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G1gat), .B(G29gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT0), .ZN(new_n256_));
  INV_X1    g055(.A(G57gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(G85gat), .ZN(new_n259_));
  AND2_X1   g058(.A1(new_n243_), .A2(new_n244_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n252_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n259_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n254_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n251_), .A2(new_n261_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n249_), .A2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n243_), .A2(new_n244_), .A3(new_n252_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n259_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT33), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n266_), .A2(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n264_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n269_), .B1(new_n272_), .B2(new_n268_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n263_), .A2(new_n271_), .A3(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT22), .B(G169gat), .ZN(new_n275_));
  INV_X1    g074(.A(G176gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G169gat), .A2(G176gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT84), .ZN(new_n280_));
  AND3_X1   g079(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n281_));
  AOI21_X1  g080(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  OR2_X1    g082(.A1(G183gat), .A2(G190gat), .ZN(new_n284_));
  AOI22_X1  g083(.A1(new_n279_), .A2(new_n280_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n278_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n286_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT84), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT25), .B(G183gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT26), .B(G190gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(new_n283_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(G169gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(new_n276_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(new_n278_), .ZN(new_n296_));
  MUX2_X1   g095(.A(new_n295_), .B(new_n296_), .S(KEYINPUT24), .Z(new_n297_));
  AOI22_X1  g096(.A1(new_n285_), .A2(new_n288_), .B1(new_n293_), .B2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(G204gat), .ZN(new_n299_));
  OAI21_X1  g098(.A(KEYINPUT92), .B1(new_n299_), .B2(G197gat), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT92), .ZN(new_n301_));
  INV_X1    g100(.A(G197gat), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n301_), .A2(new_n302_), .A3(G204gat), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT21), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n299_), .A2(G197gat), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n300_), .A2(new_n303_), .A3(new_n304_), .A4(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G211gat), .B(G218gat), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT91), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n308_), .B1(new_n299_), .B2(G197gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n302_), .A2(KEYINPUT91), .A3(G204gat), .ZN(new_n310_));
  AND3_X1   g109(.A1(new_n309_), .A2(new_n310_), .A3(new_n305_), .ZN(new_n311_));
  OAI211_X1 g110(.A(new_n306_), .B(new_n307_), .C1(new_n311_), .C2(new_n304_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n307_), .A2(new_n304_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n300_), .A2(new_n303_), .A3(new_n305_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n312_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(KEYINPUT99), .B1(new_n298_), .B2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n293_), .A2(new_n297_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n288_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n283_), .A2(new_n284_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n321_), .B1(new_n287_), .B2(KEYINPUT84), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n319_), .B1(new_n320_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT99), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n323_), .A2(new_n324_), .A3(new_n316_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n318_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT98), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT97), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n287_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n321_), .B1(new_n287_), .B2(new_n328_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n327_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n279_), .A2(KEYINPUT97), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n333_), .A2(KEYINPUT98), .A3(new_n321_), .A4(new_n329_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(KEYINPUT96), .B(KEYINPUT24), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n296_), .A2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n335_), .A2(new_n294_), .A3(new_n276_), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n336_), .A2(new_n283_), .A3(new_n291_), .A4(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n332_), .A2(new_n334_), .A3(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(KEYINPUT100), .B1(new_n339_), .B2(new_n316_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n338_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n333_), .A2(new_n321_), .A3(new_n329_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n341_), .B1(new_n342_), .B2(new_n327_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT100), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n343_), .A2(new_n344_), .A3(new_n317_), .A4(new_n334_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G226gat), .A2(G233gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT19), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT20), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n326_), .A2(new_n340_), .A3(new_n345_), .A4(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n317_), .B1(new_n343_), .B2(new_n334_), .ZN(new_n351_));
  OAI21_X1  g150(.A(KEYINPUT20), .B1(new_n323_), .B2(new_n316_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n347_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n350_), .A2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G8gat), .B(G36gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT18), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(G64gat), .ZN(new_n357_));
  INV_X1    g156(.A(G92gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n354_), .A2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n350_), .A2(new_n359_), .A3(new_n353_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n202_), .B1(new_n274_), .B2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n339_), .A2(new_n316_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n347_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n348_), .B1(new_n298_), .B2(new_n317_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n365_), .A2(new_n366_), .A3(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n338_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n369_));
  OAI21_X1  g168(.A(KEYINPUT20), .B1(new_n369_), .B2(new_n316_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n370_), .B1(new_n318_), .B2(new_n325_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n368_), .B1(new_n371_), .B2(new_n366_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n350_), .A2(KEYINPUT104), .A3(new_n353_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n359_), .A2(KEYINPUT32), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n373_), .A2(new_n374_), .A3(new_n376_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n375_), .B1(new_n354_), .B2(KEYINPUT104), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n268_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n266_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n259_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n267_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n382_), .B1(new_n272_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n381_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n379_), .A2(new_n385_), .ZN(new_n386_));
  AND3_X1   g185(.A1(new_n350_), .A2(new_n359_), .A3(new_n353_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n359_), .B1(new_n350_), .B2(new_n353_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  AOI22_X1  g188(.A1(new_n266_), .A2(new_n270_), .B1(new_n254_), .B2(new_n262_), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n389_), .A2(new_n390_), .A3(KEYINPUT103), .A4(new_n273_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n364_), .A2(new_n386_), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT94), .ZN(new_n393_));
  AOI22_X1  g192(.A1(new_n227_), .A2(KEYINPUT29), .B1(new_n312_), .B2(new_n315_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G228gat), .A2(G233gat), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n393_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n395_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT29), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n398_), .B1(new_n231_), .B2(new_n214_), .ZN(new_n399_));
  OAI211_X1 g198(.A(KEYINPUT94), .B(new_n397_), .C1(new_n317_), .C2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n396_), .A2(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n229_), .A2(KEYINPUT29), .A3(new_n232_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT93), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n395_), .B(KEYINPUT90), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n404_), .B1(new_n312_), .B2(new_n315_), .ZN(new_n405_));
  AND3_X1   g204(.A1(new_n402_), .A2(new_n403_), .A3(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n403_), .B1(new_n402_), .B2(new_n405_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n401_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G78gat), .B(G106gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n409_), .ZN(new_n411_));
  OAI211_X1 g210(.A(new_n401_), .B(new_n411_), .C1(new_n406_), .C2(new_n407_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n229_), .A2(new_n232_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(new_n398_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G22gat), .B(G50gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT28), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n416_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n413_), .A2(new_n398_), .A3(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n410_), .A2(new_n412_), .A3(new_n420_), .ZN(new_n421_));
  AND3_X1   g220(.A1(new_n410_), .A2(KEYINPUT95), .A3(new_n412_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT89), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n420_), .A2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n417_), .A2(KEYINPUT89), .A3(new_n419_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT95), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n408_), .A2(new_n427_), .A3(new_n409_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n426_), .A2(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n421_), .B1(new_n422_), .B2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n392_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT107), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n385_), .A2(KEYINPUT105), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT105), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n381_), .A2(new_n384_), .A3(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n430_), .A2(new_n434_), .A3(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n362_), .A2(KEYINPUT106), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT27), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n439_), .B1(new_n372_), .B2(new_n360_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT106), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n350_), .A2(new_n441_), .A3(new_n353_), .A4(new_n359_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n438_), .A2(new_n440_), .A3(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n439_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n433_), .B1(new_n437_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n436_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n435_), .B1(new_n381_), .B2(new_n384_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n443_), .A2(new_n444_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n449_), .A2(new_n450_), .A3(KEYINPUT107), .A4(new_n430_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n432_), .A2(new_n446_), .A3(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(G227gat), .ZN(new_n453_));
  INV_X1    g252(.A(G233gat), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n298_), .B(KEYINPUT30), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT85), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n323_), .B(KEYINPUT30), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT85), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n455_), .B1(new_n457_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G71gat), .B(G99gat), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n457_), .A2(new_n460_), .A3(new_n455_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n462_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n465_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n463_), .B1(new_n467_), .B2(new_n461_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n242_), .B(KEYINPUT31), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G15gat), .B(G43gat), .ZN(new_n471_));
  XOR2_X1   g270(.A(new_n470_), .B(new_n471_), .Z(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n469_), .A2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n466_), .A2(new_n468_), .A3(new_n472_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n452_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT108), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT108), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n452_), .A2(new_n480_), .A3(new_n477_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n476_), .A2(new_n449_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n450_), .A2(KEYINPUT109), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT109), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n445_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  NOR3_X1   g285(.A1(new_n482_), .A2(new_n486_), .A3(new_n430_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n479_), .A2(new_n481_), .A3(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT13), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT72), .ZN(new_n491_));
  NOR2_X1   g290(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n492_), .A2(G85gat), .A3(G92gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G85gat), .B(G92gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n493_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT65), .ZN(new_n497_));
  XNOR2_X1  g296(.A(KEYINPUT10), .B(G99gat), .ZN(new_n498_));
  OR2_X1    g297(.A1(new_n498_), .A2(G106gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G99gat), .A2(G106gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT6), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n497_), .A2(new_n499_), .A3(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT8), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT66), .ZN(new_n504_));
  INV_X1    g303(.A(G99gat), .ZN(new_n505_));
  INV_X1    g304(.A(G106gat), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n504_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT7), .ZN(new_n508_));
  OAI21_X1  g307(.A(KEYINPUT66), .B1(G99gat), .B2(G106gat), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n507_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT67), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n505_), .A2(new_n506_), .ZN(new_n513_));
  AOI22_X1  g312(.A1(new_n510_), .A2(new_n511_), .B1(KEYINPUT7), .B2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(KEYINPUT68), .B(KEYINPUT6), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT69), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n516_), .B1(G99gat), .B2(G106gat), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n500_), .A2(KEYINPUT69), .ZN(new_n518_));
  OR3_X1    g317(.A1(new_n515_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n515_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n512_), .A2(new_n514_), .A3(new_n519_), .A4(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n494_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n503_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n512_), .A2(new_n514_), .A3(new_n501_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n494_), .A2(KEYINPUT8), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n502_), .B1(new_n523_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G57gat), .B(G64gat), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n529_), .A2(KEYINPUT11), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G71gat), .B(G78gat), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n529_), .A2(KEYINPUT11), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n529_), .A2(new_n531_), .A3(KEYINPUT11), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT70), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n528_), .A2(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n527_), .A2(new_n537_), .ZN(new_n540_));
  OAI211_X1 g339(.A(G230gat), .B(G233gat), .C1(new_n539_), .C2(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(KEYINPUT12), .B1(new_n527_), .B2(new_n537_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G230gat), .A2(G233gat), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n528_), .A2(new_n538_), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n527_), .A2(KEYINPUT12), .A3(new_n535_), .A4(new_n534_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n543_), .A2(new_n544_), .A3(new_n545_), .A4(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n541_), .A2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G120gat), .B(G148gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(new_n299_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(KEYINPUT5), .B(G176gat), .ZN(new_n551_));
  XOR2_X1   g350(.A(new_n550_), .B(new_n551_), .Z(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n491_), .B1(new_n548_), .B2(new_n553_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n541_), .A2(new_n547_), .A3(KEYINPUT72), .A4(new_n552_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT73), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n552_), .B(KEYINPUT71), .Z(new_n558_));
  NAND2_X1  g357(.A1(new_n548_), .A2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n556_), .A2(new_n557_), .A3(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n557_), .B1(new_n556_), .B2(new_n559_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n490_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n556_), .A2(new_n559_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT73), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n565_), .A2(KEYINPUT13), .A3(new_n560_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G15gat), .B(G22gat), .ZN(new_n567_));
  INV_X1    g366(.A(G1gat), .ZN(new_n568_));
  INV_X1    g367(.A(G8gat), .ZN(new_n569_));
  OAI21_X1  g368(.A(KEYINPUT14), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n567_), .A2(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G1gat), .B(G8gat), .ZN(new_n572_));
  XOR2_X1   g371(.A(new_n571_), .B(new_n572_), .Z(new_n573_));
  XNOR2_X1  g372(.A(G29gat), .B(G36gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G43gat), .B(G50gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n573_), .A2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n571_), .B(new_n572_), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n574_), .B(new_n575_), .Z(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n577_), .A2(KEYINPUT79), .A3(new_n580_), .ZN(new_n581_));
  OR3_X1    g380(.A1(new_n573_), .A2(KEYINPUT79), .A3(new_n576_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G229gat), .A2(G233gat), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n581_), .A2(new_n582_), .A3(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT80), .ZN(new_n586_));
  INV_X1    g385(.A(new_n577_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT15), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n576_), .A2(KEYINPUT74), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n576_), .A2(KEYINPUT74), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n588_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n576_), .A2(KEYINPUT74), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n593_), .A2(KEYINPUT15), .A3(new_n589_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n587_), .B1(new_n595_), .B2(new_n578_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT81), .ZN(new_n597_));
  AND3_X1   g396(.A1(new_n596_), .A2(new_n597_), .A3(new_n583_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n597_), .B1(new_n596_), .B2(new_n583_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n586_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G113gat), .B(G141gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(G169gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(new_n302_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n600_), .A2(new_n604_), .ZN(new_n605_));
  OAI211_X1 g404(.A(new_n586_), .B(new_n603_), .C1(new_n598_), .C2(new_n599_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT82), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT83), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n606_), .A2(new_n607_), .A3(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n608_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n605_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n606_), .A2(new_n607_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(KEYINPUT83), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n614_), .A2(new_n600_), .A3(new_n604_), .A4(new_n609_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n612_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n563_), .A2(new_n566_), .A3(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(G231gat), .A2(G233gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n578_), .B(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n537_), .B(new_n620_), .ZN(new_n621_));
  XOR2_X1   g420(.A(G183gat), .B(G211gat), .Z(new_n622_));
  XNOR2_X1  g421(.A(G127gat), .B(G155gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  XOR2_X1   g423(.A(KEYINPUT77), .B(KEYINPUT16), .Z(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT17), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n621_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n620_), .A2(new_n536_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n629_), .A2(KEYINPUT17), .A3(new_n626_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n620_), .A2(new_n536_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n628_), .A2(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT78), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT35), .ZN(new_n635_));
  NAND2_X1  g434(.A1(G232gat), .A2(G233gat), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT34), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  AOI22_X1  g437(.A1(new_n528_), .A2(new_n576_), .B1(new_n635_), .B2(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n595_), .A2(new_n527_), .A3(KEYINPUT75), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(KEYINPUT75), .B1(new_n595_), .B2(new_n527_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n639_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n638_), .A2(new_n635_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n642_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(new_n640_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n644_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n647_), .A2(new_n648_), .A3(new_n639_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n645_), .A2(new_n649_), .A3(KEYINPUT76), .ZN(new_n650_));
  XNOR2_X1  g449(.A(G190gat), .B(G218gat), .ZN(new_n651_));
  XNOR2_X1  g450(.A(G134gat), .B(G162gat), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n651_), .B(new_n652_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n653_), .A2(KEYINPUT36), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n650_), .A2(new_n655_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n645_), .A2(new_n649_), .A3(KEYINPUT76), .A4(new_n654_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n653_), .A2(KEYINPUT36), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n659_), .B1(new_n645_), .B2(new_n649_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(KEYINPUT37), .B1(new_n658_), .B2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT37), .ZN(new_n663_));
  AOI211_X1 g462(.A(new_n663_), .B(new_n660_), .C1(new_n656_), .C2(new_n657_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n634_), .B1(new_n662_), .B2(new_n664_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n618_), .A2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n489_), .A2(new_n666_), .ZN(new_n667_));
  NOR3_X1   g466(.A1(new_n667_), .A2(G1gat), .A3(new_n449_), .ZN(new_n668_));
  XOR2_X1   g467(.A(new_n668_), .B(KEYINPUT38), .Z(new_n669_));
  AND3_X1   g468(.A1(new_n452_), .A2(new_n480_), .A3(new_n477_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n480_), .B1(new_n452_), .B2(new_n477_), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n670_), .A2(new_n671_), .A3(new_n487_), .ZN(new_n672_));
  AND3_X1   g471(.A1(new_n658_), .A2(KEYINPUT110), .A3(new_n661_), .ZN(new_n673_));
  AOI21_X1  g472(.A(KEYINPUT110), .B1(new_n658_), .B2(new_n661_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n672_), .A2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n633_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n618_), .A2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(G1gat), .B1(new_n680_), .B2(new_n449_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n669_), .A2(new_n681_), .ZN(G1324gat));
  NAND4_X1  g481(.A1(new_n489_), .A2(new_n569_), .A3(new_n486_), .A4(new_n666_), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n489_), .A2(new_n679_), .A3(new_n675_), .A4(new_n486_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT39), .ZN(new_n685_));
  AND3_X1   g484(.A1(new_n684_), .A2(new_n685_), .A3(G8gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n685_), .B1(new_n684_), .B2(G8gat), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n683_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(KEYINPUT111), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT111), .ZN(new_n690_));
  OAI211_X1 g489(.A(new_n690_), .B(new_n683_), .C1(new_n686_), .C2(new_n687_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n691_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(KEYINPUT112), .B(KEYINPUT40), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n692_), .A2(new_n694_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n689_), .A2(new_n693_), .A3(new_n691_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(G1325gat));
  OAI21_X1  g496(.A(G15gat), .B1(new_n680_), .B2(new_n477_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(KEYINPUT113), .B(KEYINPUT41), .ZN(new_n699_));
  OR2_X1    g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n698_), .A2(new_n699_), .ZN(new_n701_));
  OR3_X1    g500(.A1(new_n667_), .A2(G15gat), .A3(new_n477_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n700_), .A2(new_n701_), .A3(new_n702_), .ZN(G1326gat));
  OR3_X1    g502(.A1(new_n667_), .A2(G22gat), .A3(new_n431_), .ZN(new_n704_));
  OAI21_X1  g503(.A(G22gat), .B1(new_n680_), .B2(new_n431_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n705_), .A2(KEYINPUT42), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n705_), .A2(KEYINPUT42), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n704_), .B1(new_n706_), .B2(new_n707_), .ZN(G1327gat));
  NAND2_X1  g507(.A1(new_n489_), .A2(new_n676_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n618_), .A2(new_n634_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n449_), .ZN(new_n714_));
  AOI21_X1  g513(.A(G29gat), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n662_), .A2(new_n664_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT43), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT114), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n718_), .B1(new_n716_), .B2(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n487_), .B1(new_n478_), .B2(KEYINPUT108), .ZN(new_n721_));
  AOI211_X1 g520(.A(new_n717_), .B(new_n720_), .C1(new_n721_), .C2(new_n481_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n720_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n723_), .B1(new_n489_), .B2(new_n716_), .ZN(new_n724_));
  OAI211_X1 g523(.A(KEYINPUT44), .B(new_n711_), .C1(new_n722_), .C2(new_n724_), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n725_), .A2(G29gat), .A3(new_n714_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n711_), .B1(new_n722_), .B2(new_n724_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n715_), .B1(new_n726_), .B2(new_n729_), .ZN(G1328gat));
  INV_X1    g529(.A(KEYINPUT46), .ZN(new_n731_));
  INV_X1    g530(.A(G36gat), .ZN(new_n732_));
  INV_X1    g531(.A(new_n486_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n711_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n720_), .B1(new_n672_), .B2(new_n717_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n489_), .A2(new_n716_), .A3(new_n723_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n734_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n733_), .B1(new_n737_), .B2(KEYINPUT44), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n732_), .B1(new_n738_), .B2(new_n729_), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n710_), .A2(new_n732_), .A3(new_n486_), .A4(new_n711_), .ZN(new_n740_));
  XOR2_X1   g539(.A(KEYINPUT115), .B(KEYINPUT45), .Z(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n740_), .B(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n731_), .B1(new_n739_), .B2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n725_), .A2(new_n486_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n737_), .A2(KEYINPUT44), .ZN(new_n746_));
  OAI21_X1  g545(.A(G36gat), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n740_), .B(new_n741_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n747_), .A2(KEYINPUT46), .A3(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n744_), .A2(new_n749_), .ZN(G1329gat));
  INV_X1    g549(.A(G43gat), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n751_), .B1(new_n712_), .B2(new_n477_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n725_), .A2(G43gat), .A3(new_n476_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n752_), .B1(new_n753_), .B2(new_n746_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(KEYINPUT47), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT47), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n756_), .B(new_n752_), .C1(new_n753_), .C2(new_n746_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(G1330gat));
  OR3_X1    g557(.A1(new_n712_), .A2(G50gat), .A3(new_n431_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT116), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n725_), .A2(new_n430_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n760_), .B1(new_n761_), .B2(new_n746_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(G50gat), .ZN(new_n763_));
  NOR3_X1   g562(.A1(new_n761_), .A2(new_n746_), .A3(new_n760_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n759_), .B1(new_n763_), .B2(new_n764_), .ZN(G1331gat));
  AND2_X1   g564(.A1(new_n563_), .A2(new_n566_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n766_), .A2(new_n617_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n634_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n677_), .ZN(new_n771_));
  NOR3_X1   g570(.A1(new_n771_), .A2(new_n257_), .A3(new_n449_), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n768_), .A2(new_n672_), .A3(new_n665_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n449_), .B1(new_n773_), .B2(KEYINPUT117), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n774_), .B1(KEYINPUT117), .B2(new_n773_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n772_), .B1(new_n775_), .B2(new_n257_), .ZN(G1332gat));
  INV_X1    g575(.A(G64gat), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n773_), .A2(new_n777_), .A3(new_n486_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT48), .ZN(new_n779_));
  INV_X1    g578(.A(new_n771_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(new_n486_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n779_), .B1(new_n781_), .B2(G64gat), .ZN(new_n782_));
  AOI211_X1 g581(.A(KEYINPUT48), .B(new_n777_), .C1(new_n780_), .C2(new_n486_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n778_), .B1(new_n782_), .B2(new_n783_), .ZN(G1333gat));
  INV_X1    g583(.A(G71gat), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n773_), .A2(new_n785_), .A3(new_n476_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT49), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n780_), .A2(new_n476_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n787_), .B1(new_n788_), .B2(G71gat), .ZN(new_n789_));
  AOI211_X1 g588(.A(KEYINPUT49), .B(new_n785_), .C1(new_n780_), .C2(new_n476_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n786_), .B1(new_n789_), .B2(new_n790_), .ZN(G1334gat));
  INV_X1    g590(.A(G78gat), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n773_), .A2(new_n792_), .A3(new_n430_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT50), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n780_), .A2(new_n430_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n794_), .B1(new_n795_), .B2(G78gat), .ZN(new_n796_));
  AOI211_X1 g595(.A(KEYINPUT50), .B(new_n792_), .C1(new_n780_), .C2(new_n430_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n793_), .B1(new_n796_), .B2(new_n797_), .ZN(G1335gat));
  NAND2_X1  g597(.A1(new_n767_), .A2(new_n769_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n799_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(G85gat), .B1(new_n801_), .B2(new_n449_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n709_), .A2(new_n799_), .ZN(new_n803_));
  INV_X1    g602(.A(G85gat), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n803_), .A2(new_n804_), .A3(new_n714_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n802_), .A2(new_n805_), .ZN(G1336gat));
  OAI21_X1  g605(.A(G92gat), .B1(new_n801_), .B2(new_n733_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n803_), .A2(new_n358_), .A3(new_n486_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(G1337gat));
  INV_X1    g608(.A(KEYINPUT51), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT118), .ZN(new_n811_));
  INV_X1    g610(.A(new_n799_), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n476_), .B(new_n812_), .C1(new_n722_), .C2(new_n724_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(G99gat), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n477_), .A2(new_n498_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  NOR3_X1   g615(.A1(new_n709_), .A2(new_n799_), .A3(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n811_), .B1(new_n814_), .B2(new_n818_), .ZN(new_n819_));
  AOI211_X1 g618(.A(KEYINPUT118), .B(new_n817_), .C1(new_n813_), .C2(G99gat), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n810_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n505_), .B1(new_n800_), .B2(new_n476_), .ZN(new_n822_));
  OAI21_X1  g621(.A(KEYINPUT118), .B1(new_n822_), .B2(new_n817_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n814_), .A2(new_n818_), .A3(new_n811_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(KEYINPUT51), .A3(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n821_), .A2(new_n825_), .ZN(G1338gat));
  NAND3_X1  g625(.A1(new_n803_), .A2(new_n506_), .A3(new_n430_), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n430_), .B(new_n812_), .C1(new_n722_), .C2(new_n724_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT52), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n828_), .A2(new_n829_), .A3(G106gat), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n829_), .B1(new_n828_), .B2(G106gat), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n827_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT53), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT53), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n834_), .B(new_n827_), .C1(new_n830_), .C2(new_n831_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n835_), .ZN(G1339gat));
  INV_X1    g635(.A(KEYINPUT59), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n733_), .A2(new_n431_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n476_), .A2(new_n714_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n612_), .A2(new_n615_), .A3(new_n556_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n545_), .A2(new_n546_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n843_), .A2(KEYINPUT55), .A3(new_n544_), .A4(new_n543_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT55), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n547_), .A2(new_n845_), .ZN(new_n846_));
  OAI211_X1 g645(.A(G230gat), .B(G233gat), .C1(new_n842_), .C2(new_n542_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n844_), .A2(new_n846_), .A3(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT120), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n844_), .A2(new_n846_), .A3(KEYINPUT120), .A4(new_n847_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n558_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT56), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n852_), .A2(KEYINPUT56), .A3(new_n558_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n841_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n596_), .A2(new_n584_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n581_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n858_), .A2(new_n604_), .A3(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n606_), .A2(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n861_), .B1(new_n565_), .B2(new_n560_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n675_), .B1(new_n857_), .B2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(KEYINPUT57), .ZN(new_n864_));
  INV_X1    g663(.A(new_n861_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n865_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n866_));
  AND3_X1   g665(.A1(new_n852_), .A2(KEYINPUT56), .A3(new_n558_), .ZN(new_n867_));
  AOI21_X1  g666(.A(KEYINPUT56), .B1(new_n852_), .B2(new_n558_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n866_), .B1(new_n869_), .B2(new_n841_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT57), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n870_), .A2(new_n871_), .A3(new_n675_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n864_), .A2(new_n872_), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n556_), .B(new_n865_), .C1(new_n867_), .C2(new_n868_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT58), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n717_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n876_), .B1(new_n875_), .B2(new_n874_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n634_), .B1(new_n873_), .B2(new_n877_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n563_), .A2(new_n566_), .A3(new_n616_), .ZN(new_n879_));
  OAI21_X1  g678(.A(KEYINPUT54), .B1(new_n879_), .B2(new_n665_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(KEYINPUT119), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT119), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n882_), .B(KEYINPUT54), .C1(new_n879_), .C2(new_n665_), .ZN(new_n883_));
  OR3_X1    g682(.A1(new_n879_), .A2(KEYINPUT54), .A3(new_n665_), .ZN(new_n884_));
  AND3_X1   g683(.A1(new_n881_), .A2(new_n883_), .A3(new_n884_), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n837_), .B(new_n840_), .C1(new_n878_), .C2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n840_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n863_), .A2(KEYINPUT57), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n871_), .B1(new_n870_), .B2(new_n675_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n877_), .B1(new_n888_), .B2(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(new_n678_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n881_), .A2(new_n883_), .A3(new_n884_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n887_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n886_), .B1(new_n893_), .B2(new_n837_), .ZN(new_n894_));
  OAI21_X1  g693(.A(G113gat), .B1(new_n894_), .B2(new_n616_), .ZN(new_n895_));
  INV_X1    g694(.A(G113gat), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n893_), .A2(new_n896_), .A3(new_n617_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n897_), .ZN(G1340gat));
  OAI21_X1  g697(.A(G120gat), .B1(new_n894_), .B2(new_n766_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT60), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n900_), .B1(new_n766_), .B2(G120gat), .ZN(new_n901_));
  OAI211_X1 g700(.A(new_n893_), .B(new_n901_), .C1(new_n900_), .C2(G120gat), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n899_), .A2(new_n902_), .ZN(G1341gat));
  OAI21_X1  g702(.A(G127gat), .B1(new_n894_), .B2(new_n678_), .ZN(new_n904_));
  INV_X1    g703(.A(G127gat), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n893_), .A2(new_n905_), .A3(new_n634_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n904_), .A2(new_n906_), .ZN(G1342gat));
  OAI21_X1  g706(.A(G134gat), .B1(new_n894_), .B2(new_n717_), .ZN(new_n908_));
  INV_X1    g707(.A(G134gat), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n893_), .A2(new_n909_), .A3(new_n676_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n908_), .A2(new_n910_), .ZN(G1343gat));
  AOI21_X1  g710(.A(new_n633_), .B1(new_n873_), .B2(new_n877_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n912_), .A2(new_n885_), .ZN(new_n913_));
  NAND4_X1  g712(.A1(new_n733_), .A2(new_n714_), .A3(new_n477_), .A4(new_n430_), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n913_), .A2(new_n616_), .A3(new_n914_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(new_n210_), .ZN(G1344gat));
  NOR3_X1   g715(.A1(new_n913_), .A2(new_n766_), .A3(new_n914_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(KEYINPUT121), .B(G148gat), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n917_), .B(new_n918_), .ZN(G1345gat));
  NOR3_X1   g718(.A1(new_n913_), .A2(new_n769_), .A3(new_n914_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(KEYINPUT61), .B(G155gat), .ZN(new_n921_));
  INV_X1    g720(.A(new_n921_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n920_), .B(new_n922_), .ZN(G1346gat));
  NOR2_X1   g722(.A1(new_n913_), .A2(new_n914_), .ZN(new_n924_));
  AOI21_X1  g723(.A(G162gat), .B1(new_n924_), .B2(new_n676_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n716_), .A2(G162gat), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(KEYINPUT122), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n925_), .B1(new_n924_), .B2(new_n927_), .ZN(G1347gat));
  NOR3_X1   g727(.A1(new_n733_), .A2(new_n482_), .A3(new_n430_), .ZN(new_n929_));
  OAI211_X1 g728(.A(new_n617_), .B(new_n929_), .C1(new_n878_), .C2(new_n885_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n930_), .A2(G169gat), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT62), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(new_n932_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n930_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n934_));
  INV_X1    g733(.A(new_n275_), .ZN(new_n935_));
  OAI211_X1 g734(.A(new_n933_), .B(new_n934_), .C1(new_n935_), .C2(new_n930_), .ZN(G1348gat));
  NAND2_X1  g735(.A1(new_n891_), .A2(new_n892_), .ZN(new_n937_));
  INV_X1    g736(.A(KEYINPUT124), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n766_), .A2(new_n276_), .ZN(new_n939_));
  NAND4_X1  g738(.A1(new_n937_), .A2(new_n938_), .A3(new_n929_), .A4(new_n939_), .ZN(new_n940_));
  OAI211_X1 g739(.A(new_n929_), .B(new_n939_), .C1(new_n912_), .C2(new_n885_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n941_), .A2(KEYINPUT124), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n940_), .A2(new_n942_), .ZN(new_n943_));
  INV_X1    g742(.A(new_n766_), .ZN(new_n944_));
  OAI211_X1 g743(.A(new_n944_), .B(new_n929_), .C1(new_n878_), .C2(new_n885_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n945_), .A2(new_n276_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n946_), .A2(KEYINPUT123), .ZN(new_n947_));
  INV_X1    g746(.A(KEYINPUT123), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n945_), .A2(new_n948_), .A3(new_n276_), .ZN(new_n949_));
  AND3_X1   g748(.A1(new_n943_), .A2(new_n947_), .A3(new_n949_), .ZN(G1349gat));
  OR2_X1    g749(.A1(new_n878_), .A2(new_n885_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n951_), .A2(new_n929_), .ZN(new_n952_));
  INV_X1    g751(.A(new_n952_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n678_), .A2(new_n289_), .ZN(new_n954_));
  INV_X1    g753(.A(G183gat), .ZN(new_n955_));
  NAND3_X1  g754(.A1(new_n937_), .A2(new_n634_), .A3(new_n929_), .ZN(new_n956_));
  AOI22_X1  g755(.A1(new_n953_), .A2(new_n954_), .B1(new_n955_), .B2(new_n956_), .ZN(G1350gat));
  OAI21_X1  g756(.A(G190gat), .B1(new_n952_), .B2(new_n717_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n676_), .A2(new_n290_), .ZN(new_n959_));
  OAI21_X1  g758(.A(new_n958_), .B1(new_n952_), .B2(new_n959_), .ZN(G1351gat));
  NOR3_X1   g759(.A1(new_n733_), .A2(new_n476_), .A3(new_n437_), .ZN(new_n961_));
  INV_X1    g760(.A(new_n961_), .ZN(new_n962_));
  AOI21_X1  g761(.A(new_n962_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n963_), .A2(new_n617_), .ZN(new_n964_));
  XNOR2_X1  g763(.A(new_n964_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g764(.A1(new_n963_), .A2(new_n944_), .ZN(new_n966_));
  XNOR2_X1  g765(.A(new_n966_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g766(.A(new_n678_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n968_));
  OAI211_X1 g767(.A(new_n961_), .B(new_n968_), .C1(new_n912_), .C2(new_n885_), .ZN(new_n969_));
  NOR2_X1   g768(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n970_));
  AND3_X1   g769(.A1(new_n969_), .A2(KEYINPUT125), .A3(new_n970_), .ZN(new_n971_));
  AOI21_X1  g770(.A(KEYINPUT125), .B1(new_n969_), .B2(new_n970_), .ZN(new_n972_));
  NOR2_X1   g771(.A1(new_n969_), .A2(new_n970_), .ZN(new_n973_));
  NOR3_X1   g772(.A1(new_n971_), .A2(new_n972_), .A3(new_n973_), .ZN(G1354gat));
  INV_X1    g773(.A(KEYINPUT127), .ZN(new_n975_));
  AOI21_X1  g774(.A(G218gat), .B1(new_n963_), .B2(new_n676_), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n716_), .A2(G218gat), .ZN(new_n977_));
  XNOR2_X1  g776(.A(new_n977_), .B(KEYINPUT126), .ZN(new_n978_));
  INV_X1    g777(.A(new_n978_), .ZN(new_n979_));
  NOR3_X1   g778(.A1(new_n913_), .A2(new_n962_), .A3(new_n979_), .ZN(new_n980_));
  OAI21_X1  g779(.A(new_n975_), .B1(new_n976_), .B2(new_n980_), .ZN(new_n981_));
  NAND2_X1  g780(.A1(new_n963_), .A2(new_n978_), .ZN(new_n982_));
  NOR3_X1   g781(.A1(new_n913_), .A2(new_n675_), .A3(new_n962_), .ZN(new_n983_));
  OAI211_X1 g782(.A(KEYINPUT127), .B(new_n982_), .C1(new_n983_), .C2(G218gat), .ZN(new_n984_));
  NAND2_X1  g783(.A1(new_n981_), .A2(new_n984_), .ZN(G1355gat));
endmodule


