//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 0 0 0 0 0 0 0 0 1 0 1 0 1 0 0 1 0 0 1 1 0 0 0 1 0 0 1 0 0 0 1 1 0 1 1 1 0 0 0 1 0 1 0 1 0 1 0 0 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n891_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n898_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n911_, new_n912_, new_n913_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n927_, new_n928_, new_n930_,
    new_n931_, new_n932_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n941_, new_n942_, new_n943_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  INV_X1    g001(.A(G113gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G120gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n202_), .B(G113gat), .ZN(new_n206_));
  INV_X1    g005(.A(G120gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n205_), .A2(new_n208_), .ZN(new_n209_));
  XOR2_X1   g008(.A(G155gat), .B(G162gat), .Z(new_n210_));
  NAND2_X1  g009(.A1(G141gat), .A2(G148gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT2), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT77), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT3), .ZN(new_n216_));
  OAI211_X1 g015(.A(new_n213_), .B(new_n214_), .C1(new_n215_), .C2(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(G141gat), .A2(G148gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n219_));
  OAI22_X1  g018(.A1(KEYINPUT77), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n210_), .B1(new_n217_), .B2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n218_), .B(KEYINPUT76), .ZN(new_n223_));
  AND3_X1   g022(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n224_));
  AOI21_X1  g023(.A(KEYINPUT1), .B1(G155gat), .B2(G162gat), .ZN(new_n225_));
  OAI22_X1  g024(.A1(new_n224_), .A2(new_n225_), .B1(G155gat), .B2(G162gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n223_), .A2(new_n226_), .A3(new_n211_), .ZN(new_n227_));
  AND3_X1   g026(.A1(new_n222_), .A2(new_n227_), .A3(KEYINPUT78), .ZN(new_n228_));
  AOI21_X1  g027(.A(KEYINPUT78), .B1(new_n222_), .B2(new_n227_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n209_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT90), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n222_), .A2(new_n227_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n232_), .A2(new_n205_), .A3(new_n208_), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n230_), .A2(new_n231_), .A3(KEYINPUT4), .A4(new_n233_), .ZN(new_n234_));
  AND3_X1   g033(.A1(new_n230_), .A2(KEYINPUT4), .A3(new_n233_), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT90), .B1(new_n230_), .B2(KEYINPUT4), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n234_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G225gat), .A2(G233gat), .ZN(new_n238_));
  XOR2_X1   g037(.A(new_n238_), .B(KEYINPUT91), .Z(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n230_), .A2(new_n233_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n241_), .A2(new_n239_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n240_), .A2(new_n243_), .ZN(new_n244_));
  XOR2_X1   g043(.A(KEYINPUT92), .B(KEYINPUT0), .Z(new_n245_));
  XNOR2_X1  g044(.A(G1gat), .B(G29gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G57gat), .B(G85gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n244_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n249_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n240_), .A2(new_n251_), .A3(new_n243_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT27), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT88), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT22), .B(G169gat), .ZN(new_n257_));
  INV_X1    g056(.A(G176gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT73), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G169gat), .A2(G176gat), .ZN(new_n261_));
  INV_X1    g060(.A(G183gat), .ZN(new_n262_));
  INV_X1    g061(.A(G190gat), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT23), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT23), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n265_), .A2(G183gat), .A3(G190gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n262_), .A2(new_n263_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT73), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n257_), .A2(new_n270_), .A3(new_n258_), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n260_), .A2(new_n261_), .A3(new_n269_), .A4(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n266_), .A2(KEYINPUT72), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT72), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n274_), .A2(new_n265_), .A3(G183gat), .A4(G190gat), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n273_), .A2(new_n264_), .A3(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT25), .B(G183gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT26), .B(G190gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NOR3_X1   g078(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n280_), .B1(new_n282_), .B2(new_n261_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n276_), .A2(new_n279_), .A3(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n272_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(G197gat), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n286_), .A2(G204gat), .ZN(new_n287_));
  INV_X1    g086(.A(G204gat), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n288_), .A2(G197gat), .ZN(new_n289_));
  OAI21_X1  g088(.A(KEYINPUT21), .B1(new_n287_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n288_), .A2(G197gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n286_), .A2(G204gat), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT21), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n291_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G211gat), .B(G218gat), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n290_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n295_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n291_), .A2(new_n292_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n297_), .A2(KEYINPUT21), .A3(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n296_), .A2(new_n299_), .A3(KEYINPUT82), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n296_), .A2(new_n299_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT82), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n285_), .B1(new_n300_), .B2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT20), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n256_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n283_), .A2(new_n279_), .A3(new_n267_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT89), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n276_), .A2(new_n268_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n310_), .A2(new_n261_), .A3(new_n259_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(new_n301_), .ZN(new_n313_));
  AND2_X1   g112(.A1(new_n303_), .A2(new_n300_), .ZN(new_n314_));
  OAI211_X1 g113(.A(KEYINPUT88), .B(KEYINPUT20), .C1(new_n314_), .C2(new_n285_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n306_), .A2(new_n313_), .A3(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G226gat), .A2(G233gat), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n317_), .B(KEYINPUT19), .Z(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT87), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n316_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G8gat), .B(G36gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT18), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(G64gat), .ZN(new_n324_));
  INV_X1    g123(.A(G92gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n314_), .A2(new_n285_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n301_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n309_), .A2(new_n328_), .A3(new_n311_), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n327_), .A2(KEYINPUT20), .A3(new_n318_), .A4(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n321_), .A2(new_n326_), .A3(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n330_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n333_), .B1(new_n320_), .B2(new_n316_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n334_), .A2(new_n326_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n255_), .B1(new_n332_), .B2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n326_), .ZN(new_n337_));
  AND4_X1   g136(.A1(new_n319_), .A2(new_n306_), .A3(new_n313_), .A4(new_n315_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n328_), .A2(new_n311_), .A3(new_n307_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT20), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT94), .ZN(new_n341_));
  AOI22_X1  g140(.A1(new_n340_), .A2(new_n341_), .B1(new_n314_), .B2(new_n285_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n339_), .A2(KEYINPUT94), .A3(KEYINPUT20), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n318_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n337_), .B1(new_n338_), .B2(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n345_), .A2(new_n331_), .A3(KEYINPUT27), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT95), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n345_), .A2(new_n331_), .A3(KEYINPUT95), .A4(KEYINPUT27), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n336_), .A2(new_n348_), .A3(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT83), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT29), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n352_), .B1(new_n222_), .B2(new_n227_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n353_), .A2(new_n328_), .ZN(new_n354_));
  INV_X1    g153(.A(G233gat), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT81), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n356_), .A2(G228gat), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(G228gat), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n355_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n351_), .B1(new_n354_), .B2(new_n361_), .ZN(new_n362_));
  OAI211_X1 g161(.A(KEYINPUT83), .B(new_n360_), .C1(new_n353_), .C2(new_n328_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n228_), .A2(new_n229_), .ZN(new_n365_));
  OAI211_X1 g164(.A(new_n314_), .B(new_n361_), .C1(new_n365_), .C2(new_n352_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n364_), .A2(new_n366_), .ZN(new_n367_));
  XOR2_X1   g166(.A(G78gat), .B(G106gat), .Z(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n364_), .A2(new_n368_), .A3(new_n366_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(KEYINPUT79), .B(KEYINPUT28), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G22gat), .B(G50gat), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n376_), .B1(new_n365_), .B2(new_n352_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n222_), .A2(new_n227_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT78), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n222_), .A2(new_n227_), .A3(KEYINPUT78), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n380_), .A2(new_n352_), .A3(new_n381_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n382_), .A2(new_n375_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n374_), .B1(new_n377_), .B2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n365_), .A2(new_n352_), .A3(new_n376_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n382_), .A2(new_n375_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(new_n386_), .A3(new_n373_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n384_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT80), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT80), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n384_), .A2(new_n390_), .A3(new_n387_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n372_), .A2(new_n389_), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT85), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n301_), .B1(new_n232_), .B2(new_n352_), .ZN(new_n394_));
  AOI21_X1  g193(.A(KEYINPUT83), .B1(new_n394_), .B2(new_n360_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n363_), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n366_), .B(new_n393_), .C1(new_n395_), .C2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n369_), .A2(KEYINPUT84), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n398_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n364_), .A2(new_n393_), .A3(new_n366_), .A4(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  AOI22_X1  g201(.A1(new_n371_), .A2(KEYINPUT85), .B1(new_n384_), .B2(new_n387_), .ZN(new_n403_));
  AND3_X1   g202(.A1(new_n402_), .A2(new_n403_), .A3(KEYINPUT86), .ZN(new_n404_));
  AOI21_X1  g203(.A(KEYINPUT86), .B1(new_n402_), .B2(new_n403_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n392_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G227gat), .A2(G233gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n285_), .B(new_n407_), .ZN(new_n408_));
  XOR2_X1   g207(.A(new_n408_), .B(new_n209_), .Z(new_n409_));
  XOR2_X1   g208(.A(KEYINPUT74), .B(G99gat), .Z(new_n410_));
  XNOR2_X1  g209(.A(KEYINPUT30), .B(G71gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n410_), .B(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G15gat), .B(G43gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT75), .B(KEYINPUT31), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n412_), .B(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n409_), .B(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n406_), .A2(new_n418_), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n417_), .B(new_n392_), .C1(new_n404_), .C2(new_n405_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n350_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n321_), .A2(new_n330_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(new_n337_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n240_), .A2(KEYINPUT33), .A3(new_n251_), .A4(new_n243_), .ZN(new_n424_));
  AND3_X1   g223(.A1(new_n423_), .A2(new_n424_), .A3(new_n331_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n239_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n251_), .B1(new_n237_), .B2(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n427_), .B1(new_n426_), .B2(new_n241_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT93), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT33), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n252_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  AOI211_X1 g230(.A(new_n249_), .B(new_n242_), .C1(new_n237_), .C2(new_n239_), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT93), .B1(new_n432_), .B2(KEYINPUT33), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n425_), .A2(new_n428_), .A3(new_n431_), .A4(new_n433_), .ZN(new_n434_));
  OAI211_X1 g233(.A(KEYINPUT32), .B(new_n326_), .C1(new_n338_), .C2(new_n344_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT32), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n334_), .B1(new_n436_), .B2(new_n337_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n253_), .A2(new_n435_), .A3(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n406_), .B1(new_n434_), .B2(new_n438_), .ZN(new_n439_));
  AOI22_X1  g238(.A1(new_n254_), .A2(new_n421_), .B1(new_n439_), .B2(new_n418_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G230gat), .A2(G233gat), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G57gat), .B(G64gat), .ZN(new_n443_));
  OR2_X1    g242(.A1(G71gat), .A2(G78gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(G71gat), .A2(G78gat), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n443_), .A2(KEYINPUT11), .A3(new_n444_), .A4(new_n445_), .ZN(new_n446_));
  AND2_X1   g245(.A1(G57gat), .A2(G64gat), .ZN(new_n447_));
  NOR2_X1   g246(.A1(G57gat), .A2(G64gat), .ZN(new_n448_));
  OAI21_X1  g247(.A(KEYINPUT11), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n444_), .A2(new_n445_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  OR3_X1    g250(.A1(new_n447_), .A2(new_n448_), .A3(KEYINPUT11), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n446_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT65), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT65), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n446_), .A2(new_n451_), .A3(new_n455_), .A4(new_n452_), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n454_), .A2(new_n456_), .ZN(new_n457_));
  XOR2_X1   g256(.A(G85gat), .B(G92gat), .Z(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(KEYINPUT9), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G99gat), .A2(G106gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT6), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT6), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n462_), .A2(G99gat), .A3(G106gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n461_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(G106gat), .ZN(new_n465_));
  INV_X1    g264(.A(G99gat), .ZN(new_n466_));
  AND2_X1   g265(.A1(new_n466_), .A2(KEYINPUT10), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n466_), .A2(KEYINPUT10), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n465_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(G85gat), .ZN(new_n470_));
  OR3_X1    g269(.A1(new_n470_), .A2(new_n325_), .A3(KEYINPUT9), .ZN(new_n471_));
  AND4_X1   g270(.A1(new_n459_), .A2(new_n464_), .A3(new_n469_), .A4(new_n471_), .ZN(new_n472_));
  AND2_X1   g271(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n473_));
  NOR2_X1   g272(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n474_));
  OAI22_X1  g273(.A1(new_n473_), .A2(new_n474_), .B1(G99gat), .B2(G106gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n476_), .A2(new_n466_), .A3(new_n465_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n475_), .A2(new_n464_), .A3(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(new_n458_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT8), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT8), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n478_), .A2(new_n481_), .A3(new_n458_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n472_), .B1(new_n480_), .B2(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n457_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT66), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n459_), .A2(new_n464_), .A3(new_n469_), .A4(new_n471_), .ZN(new_n486_));
  AND3_X1   g285(.A1(new_n478_), .A2(new_n481_), .A3(new_n458_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n481_), .B1(new_n478_), .B2(new_n458_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n486_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n454_), .A2(new_n456_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  OR2_X1    g290(.A1(new_n491_), .A2(KEYINPUT66), .ZN(new_n492_));
  OAI211_X1 g291(.A(new_n442_), .B(new_n485_), .C1(new_n492_), .C2(new_n484_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT67), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n453_), .A2(KEYINPUT12), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  AND3_X1   g295(.A1(new_n489_), .A2(new_n494_), .A3(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n494_), .B1(new_n489_), .B2(new_n496_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n489_), .A2(new_n490_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT12), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n500_), .B1(new_n491_), .B2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n499_), .A2(new_n441_), .A3(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n493_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G120gat), .B(G148gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT5), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(G176gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(G204gat), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n504_), .A2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n493_), .A2(new_n503_), .A3(new_n508_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n510_), .A2(KEYINPUT68), .A3(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT68), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n504_), .A2(new_n513_), .A3(new_n509_), .ZN(new_n514_));
  AND3_X1   g313(.A1(new_n512_), .A2(KEYINPUT13), .A3(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(KEYINPUT13), .B1(new_n512_), .B2(new_n514_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G15gat), .B(G22gat), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT69), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(G1gat), .ZN(new_n521_));
  INV_X1    g320(.A(G8gat), .ZN(new_n522_));
  OAI21_X1  g321(.A(KEYINPUT14), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT70), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n520_), .A2(new_n524_), .ZN(new_n525_));
  XOR2_X1   g324(.A(G1gat), .B(G8gat), .Z(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G29gat), .B(G36gat), .ZN(new_n528_));
  INV_X1    g327(.A(G43gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(G50gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n528_), .B(G43gat), .ZN(new_n532_));
  INV_X1    g331(.A(G50gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  AND2_X1   g333(.A1(new_n531_), .A2(new_n534_), .ZN(new_n535_));
  OR2_X1    g334(.A1(new_n527_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n527_), .A2(new_n535_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G229gat), .A2(G233gat), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  AND3_X1   g340(.A1(new_n531_), .A2(new_n534_), .A3(KEYINPUT15), .ZN(new_n542_));
  AOI21_X1  g341(.A(KEYINPUT15), .B1(new_n531_), .B2(new_n534_), .ZN(new_n543_));
  OR2_X1    g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n527_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n546_), .A2(new_n539_), .A3(new_n537_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n541_), .A2(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(G113gat), .B(G141gat), .Z(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(G169gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(new_n286_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n548_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n551_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n541_), .A2(new_n547_), .A3(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n552_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n517_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n440_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G231gat), .A2(G233gat), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n545_), .A2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n527_), .A2(G231gat), .A3(G233gat), .ZN(new_n562_));
  AND3_X1   g361(.A1(new_n561_), .A2(new_n562_), .A3(new_n453_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n453_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G127gat), .B(G155gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT16), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(G183gat), .ZN(new_n567_));
  OR2_X1    g366(.A1(new_n567_), .A2(G211gat), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(G211gat), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(KEYINPUT17), .ZN(new_n571_));
  NOR3_X1   g370(.A1(new_n563_), .A2(new_n564_), .A3(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT17), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n568_), .A2(new_n573_), .A3(new_n569_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n571_), .A2(KEYINPUT71), .A3(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n561_), .A2(new_n562_), .A3(new_n457_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n561_), .A2(new_n562_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(new_n490_), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n575_), .A2(new_n576_), .A3(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n571_), .A2(new_n574_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT71), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n572_), .B1(new_n579_), .B2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n544_), .A2(new_n489_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G232gat), .A2(G233gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT34), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n483_), .A2(new_n535_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n584_), .A2(KEYINPUT35), .A3(new_n586_), .A4(new_n587_), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n586_), .A2(KEYINPUT35), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n542_), .A2(new_n543_), .ZN(new_n590_));
  OAI211_X1 g389(.A(new_n587_), .B(new_n589_), .C1(new_n590_), .C2(new_n483_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n586_), .A2(KEYINPUT35), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G190gat), .B(G218gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(G134gat), .ZN(new_n595_));
  INV_X1    g394(.A(G162gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT36), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  AND3_X1   g398(.A1(new_n588_), .A2(new_n593_), .A3(new_n599_), .ZN(new_n600_));
  AOI22_X1  g399(.A1(new_n588_), .A2(new_n593_), .B1(new_n598_), .B2(new_n597_), .ZN(new_n601_));
  OAI21_X1  g400(.A(KEYINPUT37), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n588_), .A2(new_n593_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n597_), .A2(new_n598_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT37), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n588_), .A2(new_n593_), .A3(new_n599_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n605_), .A2(new_n606_), .A3(new_n607_), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n583_), .A2(new_n602_), .A3(new_n608_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n559_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT96), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n610_), .B1(new_n611_), .B2(KEYINPUT38), .ZN(new_n612_));
  NOR3_X1   g411(.A1(new_n612_), .A2(G1gat), .A3(new_n254_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(KEYINPUT38), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(KEYINPUT97), .B1(new_n600_), .B2(new_n601_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT97), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n605_), .A2(new_n617_), .A3(new_n607_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT98), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(KEYINPUT99), .B1(new_n440_), .B2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n434_), .A2(new_n438_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n406_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n623_), .A2(new_n418_), .A3(new_n624_), .ZN(new_n625_));
  AND3_X1   g424(.A1(new_n336_), .A2(new_n348_), .A3(new_n349_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n402_), .A2(new_n403_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT86), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n402_), .A2(new_n403_), .A3(KEYINPUT86), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n417_), .B1(new_n631_), .B2(new_n392_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n420_), .ZN(new_n633_));
  OAI211_X1 g432(.A(new_n626_), .B(new_n254_), .C1(new_n632_), .C2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n625_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT99), .ZN(new_n636_));
  INV_X1    g435(.A(new_n621_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n635_), .A2(new_n636_), .A3(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n622_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n583_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n558_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n639_), .A2(new_n641_), .ZN(new_n642_));
  OAI21_X1  g441(.A(G1gat), .B1(new_n642_), .B2(new_n254_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT100), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n643_), .A2(new_n644_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n615_), .B1(new_n645_), .B2(new_n646_), .ZN(G1324gat));
  AOI21_X1  g446(.A(new_n636_), .B1(new_n635_), .B2(new_n637_), .ZN(new_n648_));
  AOI211_X1 g447(.A(KEYINPUT99), .B(new_n621_), .C1(new_n625_), .C2(new_n634_), .ZN(new_n649_));
  OAI211_X1 g448(.A(new_n350_), .B(new_n641_), .C1(new_n648_), .C2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(KEYINPUT101), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT101), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n639_), .A2(new_n652_), .A3(new_n350_), .A4(new_n641_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n651_), .A2(new_n653_), .A3(G8gat), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(KEYINPUT39), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT39), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n651_), .A2(new_n653_), .A3(new_n656_), .A4(G8gat), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n610_), .A2(new_n522_), .A3(new_n350_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT40), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n658_), .A2(KEYINPUT40), .A3(new_n659_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1325gat));
  INV_X1    g463(.A(G15gat), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n610_), .A2(new_n665_), .A3(new_n417_), .ZN(new_n666_));
  OAI21_X1  g465(.A(G15gat), .B1(new_n642_), .B2(new_n418_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT41), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n667_), .A2(new_n668_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n666_), .B1(new_n669_), .B2(new_n670_), .ZN(G1326gat));
  INV_X1    g470(.A(G22gat), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n610_), .A2(new_n672_), .A3(new_n406_), .ZN(new_n673_));
  OAI21_X1  g472(.A(G22gat), .B1(new_n642_), .B2(new_n624_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n674_), .A2(KEYINPUT42), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n674_), .A2(KEYINPUT42), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n673_), .B1(new_n675_), .B2(new_n676_), .ZN(G1327gat));
  AND2_X1   g476(.A1(new_n602_), .A2(new_n608_), .ZN(new_n678_));
  OAI21_X1  g477(.A(KEYINPUT43), .B1(new_n678_), .B2(KEYINPUT102), .ZN(new_n679_));
  INV_X1    g478(.A(new_n678_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n679_), .B1(new_n635_), .B2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n679_), .ZN(new_n682_));
  AOI211_X1 g481(.A(new_n678_), .B(new_n682_), .C1(new_n625_), .C2(new_n634_), .ZN(new_n683_));
  OAI211_X1 g482(.A(new_n640_), .B(new_n557_), .C1(new_n681_), .C2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(KEYINPUT103), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n684_), .A2(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n682_), .B1(new_n440_), .B2(new_n678_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n635_), .A2(new_n680_), .A3(new_n679_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n691_), .A2(new_n640_), .A3(new_n557_), .A4(new_n686_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n688_), .A2(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(G29gat), .B1(new_n693_), .B2(new_n254_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n619_), .A2(new_n583_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n559_), .A2(new_n695_), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n254_), .A2(G29gat), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n694_), .B1(new_n696_), .B2(new_n697_), .ZN(G1328gat));
  NOR3_X1   g497(.A1(new_n696_), .A2(G36gat), .A3(new_n626_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT45), .Z(new_n700_));
  OAI21_X1  g499(.A(G36gat), .B1(new_n693_), .B2(new_n626_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT46), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n700_), .A2(KEYINPUT46), .A3(new_n701_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1329gat));
  NOR2_X1   g505(.A1(new_n418_), .A2(new_n529_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n688_), .A2(new_n692_), .A3(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(KEYINPUT104), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n529_), .B1(new_n696_), .B2(new_n418_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT104), .ZN(new_n711_));
  NAND4_X1  g510(.A1(new_n688_), .A2(new_n692_), .A3(new_n711_), .A4(new_n707_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n709_), .A2(new_n710_), .A3(new_n712_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g513(.A(G50gat), .B1(new_n693_), .B2(new_n624_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n406_), .A2(new_n533_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n715_), .B1(new_n696_), .B2(new_n716_), .ZN(G1331gat));
  INV_X1    g516(.A(new_n517_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n718_), .B1(new_n622_), .B2(new_n638_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n640_), .A2(new_n555_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT106), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n722_), .B1(new_n253_), .B2(G57gat), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n721_), .A2(new_n722_), .A3(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n635_), .A2(new_n556_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT105), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n726_), .A2(new_n718_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(new_n609_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n729_), .B(new_n253_), .C1(new_n721_), .C2(new_n723_), .ZN(new_n730_));
  INV_X1    g529(.A(G57gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n724_), .B1(new_n730_), .B2(new_n731_), .ZN(G1332gat));
  OR3_X1    g531(.A1(new_n728_), .A2(G64gat), .A3(new_n626_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n719_), .A2(new_n350_), .A3(new_n720_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT48), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n734_), .A2(new_n735_), .A3(G64gat), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n735_), .B1(new_n734_), .B2(G64gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n733_), .B1(new_n737_), .B2(new_n738_), .ZN(G1333gat));
  NAND3_X1  g538(.A1(new_n719_), .A2(new_n417_), .A3(new_n720_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT49), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n740_), .A2(new_n741_), .A3(G71gat), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n741_), .B1(new_n740_), .B2(G71gat), .ZN(new_n744_));
  OR2_X1    g543(.A1(new_n418_), .A2(G71gat), .ZN(new_n745_));
  OAI22_X1  g544(.A1(new_n743_), .A2(new_n744_), .B1(new_n728_), .B2(new_n745_), .ZN(G1334gat));
  NAND3_X1  g545(.A1(new_n719_), .A2(new_n406_), .A3(new_n720_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT50), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n747_), .A2(new_n748_), .A3(G78gat), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n748_), .B1(new_n747_), .B2(G78gat), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n624_), .A2(G78gat), .ZN(new_n752_));
  OAI22_X1  g551(.A1(new_n750_), .A2(new_n751_), .B1(new_n728_), .B2(new_n752_), .ZN(G1335gat));
  INV_X1    g552(.A(KEYINPUT105), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n725_), .B(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n755_), .A2(new_n517_), .A3(new_n695_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n470_), .B1(new_n756_), .B2(new_n254_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT107), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n718_), .A2(new_n583_), .A3(new_n555_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n691_), .A2(new_n759_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n760_), .A2(G85gat), .A3(new_n253_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n758_), .A2(new_n761_), .ZN(G1336gat));
  INV_X1    g561(.A(new_n756_), .ZN(new_n763_));
  AOI21_X1  g562(.A(G92gat), .B1(new_n763_), .B2(new_n350_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n350_), .A2(G92gat), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT108), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n764_), .B1(new_n760_), .B2(new_n766_), .ZN(G1337gat));
  OR2_X1    g566(.A1(new_n467_), .A2(new_n468_), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n727_), .A2(new_n768_), .A3(new_n417_), .A4(new_n695_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT109), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT109), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n763_), .A2(new_n771_), .A3(new_n768_), .A4(new_n417_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n760_), .A2(new_n417_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(G99gat), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n770_), .A2(new_n772_), .A3(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT51), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n770_), .A2(new_n772_), .A3(new_n777_), .A4(new_n774_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n778_), .ZN(G1338gat));
  NAND3_X1  g578(.A1(new_n763_), .A2(new_n465_), .A3(new_n406_), .ZN(new_n780_));
  XOR2_X1   g579(.A(KEYINPUT110), .B(KEYINPUT52), .Z(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n760_), .A2(new_n406_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n782_), .B1(new_n783_), .B2(G106gat), .ZN(new_n784_));
  AOI211_X1 g583(.A(new_n465_), .B(new_n781_), .C1(new_n760_), .C2(new_n406_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n780_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n787_), .B(KEYINPUT112), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n786_), .A2(new_n789_), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n780_), .B(new_n788_), .C1(new_n784_), .C2(new_n785_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(G1339gat));
  OAI211_X1 g591(.A(new_n609_), .B(new_n556_), .C1(new_n515_), .C2(new_n516_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT54), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n793_), .B(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT55), .ZN(new_n796_));
  OAI21_X1  g595(.A(KEYINPUT67), .B1(new_n483_), .B2(new_n495_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n489_), .A2(new_n494_), .A3(new_n496_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n501_), .B1(new_n457_), .B2(new_n483_), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n797_), .B(new_n798_), .C1(new_n799_), .C2(new_n484_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n796_), .B1(new_n800_), .B2(new_n442_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n800_), .A2(new_n442_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n499_), .A2(KEYINPUT55), .A3(new_n502_), .A4(new_n441_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n509_), .B1(new_n803_), .B2(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n806_), .A2(KEYINPUT113), .A3(KEYINPUT56), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT56), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n441_), .B1(new_n499_), .B2(new_n502_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n503_), .B1(new_n809_), .B2(new_n796_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n508_), .B1(new_n810_), .B2(new_n804_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT113), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n808_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n511_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n814_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n807_), .A2(new_n813_), .A3(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n538_), .A2(new_n539_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n546_), .A2(new_n540_), .A3(new_n537_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n817_), .A2(new_n551_), .A3(new_n818_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n819_), .A2(new_n554_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n512_), .A2(new_n820_), .A3(new_n514_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n816_), .A2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n619_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT57), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT58), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n511_), .B1(new_n806_), .B2(KEYINPUT56), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n820_), .B1(new_n811_), .B2(new_n808_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n826_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n814_), .B1(new_n811_), .B2(new_n808_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n806_), .A2(KEYINPUT56), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n830_), .A2(new_n831_), .A3(KEYINPUT58), .A4(new_n820_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n829_), .A2(new_n680_), .A3(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n822_), .A2(KEYINPUT57), .A3(new_n619_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n825_), .A2(new_n833_), .A3(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n795_), .B1(new_n835_), .B2(new_n640_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n350_), .A2(new_n254_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n633_), .ZN(new_n838_));
  OAI21_X1  g637(.A(KEYINPUT59), .B1(new_n836_), .B2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(KEYINPUT114), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n793_), .B(KEYINPUT54), .ZN(new_n841_));
  AOI21_X1  g640(.A(KEYINPUT57), .B1(new_n822_), .B2(new_n619_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n619_), .ZN(new_n843_));
  AOI211_X1 g642(.A(new_n824_), .B(new_n843_), .C1(new_n816_), .C2(new_n821_), .ZN(new_n844_));
  AND3_X1   g643(.A1(new_n829_), .A2(new_n680_), .A3(new_n832_), .ZN(new_n845_));
  NOR3_X1   g644(.A1(new_n842_), .A2(new_n844_), .A3(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n841_), .B1(new_n846_), .B2(new_n583_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n838_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT114), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n849_), .A2(new_n850_), .A3(KEYINPUT59), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n835_), .A2(new_n640_), .ZN(new_n852_));
  AOI21_X1  g651(.A(KEYINPUT59), .B1(new_n852_), .B2(new_n841_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n838_), .B(KEYINPUT115), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(KEYINPUT116), .B1(new_n853_), .B2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT116), .ZN(new_n857_));
  NOR4_X1   g656(.A1(new_n836_), .A2(new_n857_), .A3(KEYINPUT59), .A4(new_n854_), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n840_), .B(new_n851_), .C1(new_n856_), .C2(new_n858_), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n859_), .A2(new_n203_), .A3(new_n556_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n849_), .ZN(new_n861_));
  AOI21_X1  g660(.A(G113gat), .B1(new_n861_), .B2(new_n555_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n860_), .A2(new_n862_), .ZN(G1340gat));
  OAI21_X1  g662(.A(KEYINPUT118), .B1(new_n859_), .B2(new_n718_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(KEYINPUT117), .B(G120gat), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n850_), .B1(new_n849_), .B2(KEYINPUT59), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n867_));
  AOI211_X1 g666(.A(KEYINPUT114), .B(new_n867_), .C1(new_n847_), .C2(new_n848_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n866_), .A2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT118), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n847_), .A2(new_n867_), .A3(new_n855_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n857_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n853_), .A2(KEYINPUT116), .A3(new_n855_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n869_), .A2(new_n870_), .A3(new_n517_), .A4(new_n874_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n864_), .A2(new_n865_), .A3(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n865_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n877_), .B1(new_n718_), .B2(KEYINPUT60), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n861_), .B(new_n878_), .C1(KEYINPUT60), .C2(new_n877_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n876_), .A2(new_n879_), .ZN(G1341gat));
  INV_X1    g679(.A(G127gat), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n881_), .B1(new_n849_), .B2(new_n640_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n583_), .A2(G127gat), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n859_), .B2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(KEYINPUT119), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT119), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n886_), .B(new_n882_), .C1(new_n859_), .C2(new_n883_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n885_), .A2(new_n887_), .ZN(G1342gat));
  AOI21_X1  g687(.A(G134gat), .B1(new_n861_), .B2(new_n621_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(KEYINPUT120), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n869_), .A2(G134gat), .A3(new_n680_), .A4(new_n874_), .ZN(new_n891_));
  AND2_X1   g690(.A1(new_n890_), .A2(new_n891_), .ZN(G1343gat));
  NOR2_X1   g691(.A1(new_n836_), .A2(new_n419_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(new_n837_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n555_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n517_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g698(.A(KEYINPUT121), .ZN(new_n900_));
  NAND4_X1  g699(.A1(new_n893_), .A2(new_n900_), .A3(new_n583_), .A4(new_n837_), .ZN(new_n901_));
  NAND4_X1  g700(.A1(new_n847_), .A2(new_n632_), .A3(new_n583_), .A4(new_n837_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(KEYINPUT121), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n901_), .A2(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(KEYINPUT61), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT61), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n901_), .A2(new_n903_), .A3(new_n906_), .ZN(new_n907_));
  AND3_X1   g706(.A1(new_n905_), .A2(G155gat), .A3(new_n907_), .ZN(new_n908_));
  AOI21_X1  g707(.A(G155gat), .B1(new_n905_), .B2(new_n907_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n908_), .A2(new_n909_), .ZN(G1346gat));
  OAI21_X1  g709(.A(new_n596_), .B1(new_n894_), .B2(new_n637_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n680_), .A2(G162gat), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n911_), .B1(new_n894_), .B2(new_n912_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(KEYINPUT122), .ZN(G1347gat));
  NOR2_X1   g713(.A1(new_n836_), .A2(new_n420_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n626_), .A2(new_n253_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(new_n917_));
  OAI21_X1  g716(.A(G169gat), .B1(new_n917_), .B2(new_n556_), .ZN(new_n918_));
  NAND4_X1  g717(.A1(new_n915_), .A2(new_n257_), .A3(new_n555_), .A4(new_n916_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(new_n920_));
  MUX2_X1   g719(.A(new_n918_), .B(new_n920_), .S(KEYINPUT62), .Z(G1348gat));
  NOR2_X1   g720(.A1(new_n917_), .A2(new_n718_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n258_), .A2(KEYINPUT123), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  XOR2_X1   g723(.A(KEYINPUT123), .B(G176gat), .Z(new_n925_));
  AOI21_X1  g724(.A(new_n924_), .B1(new_n922_), .B2(new_n925_), .ZN(G1349gat));
  NOR2_X1   g725(.A1(new_n917_), .A2(new_n640_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(new_n277_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n928_), .B1(new_n262_), .B2(new_n927_), .ZN(G1350gat));
  OAI21_X1  g728(.A(G190gat), .B1(new_n917_), .B2(new_n678_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n621_), .A2(new_n278_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(KEYINPUT124), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n930_), .B1(new_n917_), .B2(new_n932_), .ZN(G1351gat));
  NAND3_X1  g732(.A1(new_n893_), .A2(KEYINPUT125), .A3(new_n916_), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n847_), .A2(new_n632_), .A3(new_n916_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT125), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n934_), .A2(new_n937_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n938_), .A2(new_n555_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n939_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g739(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n941_));
  XNOR2_X1  g740(.A(KEYINPUT126), .B(G204gat), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n938_), .A2(new_n517_), .ZN(new_n943_));
  MUX2_X1   g742(.A(new_n941_), .B(new_n942_), .S(new_n943_), .Z(G1353gat));
  OR2_X1    g743(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n945_));
  NAND2_X1  g744(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n946_));
  AND4_X1   g745(.A1(new_n583_), .A2(new_n938_), .A3(new_n945_), .A4(new_n946_), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n945_), .B1(new_n938_), .B2(new_n583_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n947_), .A2(new_n948_), .ZN(G1354gat));
  INV_X1    g748(.A(G218gat), .ZN(new_n950_));
  AOI211_X1 g749(.A(new_n950_), .B(new_n678_), .C1(new_n934_), .C2(new_n937_), .ZN(new_n951_));
  AOI21_X1  g750(.A(KEYINPUT127), .B1(new_n938_), .B2(new_n621_), .ZN(new_n952_));
  INV_X1    g751(.A(KEYINPUT127), .ZN(new_n953_));
  AOI211_X1 g752(.A(new_n953_), .B(new_n637_), .C1(new_n934_), .C2(new_n937_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n952_), .A2(new_n954_), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n951_), .B1(new_n955_), .B2(new_n950_), .ZN(G1355gat));
endmodule


