//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 1 1 1 1 1 1 0 0 1 0 1 0 1 1 0 0 0 0 1 0 1 1 0 1 0 0 1 1 1 0 0 0 1 0 0 0 0 1 1 0 1 0 0 1 0 0 1 1 0 1 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n837_, new_n838_, new_n839_, new_n841_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n858_, new_n859_, new_n860_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_,
    new_n877_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n948_, new_n949_, new_n951_, new_n952_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n959_, new_n961_,
    new_n962_, new_n964_, new_n965_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n986_, new_n987_, new_n988_,
    new_n989_, new_n990_, new_n991_, new_n992_, new_n994_, new_n995_,
    new_n996_, new_n997_, new_n999_, new_n1000_, new_n1002_, new_n1003_,
    new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1010_, new_n1011_,
    new_n1012_, new_n1013_, new_n1015_, new_n1016_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G99gat), .A2(G106gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT7), .ZN(new_n205_));
  NAND3_X1  g004(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  AOI21_X1  g006(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT67), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n208_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT67), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n210_), .A2(new_n211_), .A3(new_n206_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n205_), .A2(new_n209_), .A3(new_n212_), .ZN(new_n213_));
  AND2_X1   g012(.A1(G85gat), .A2(G92gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G85gat), .A2(G92gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n213_), .A2(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n207_), .A2(new_n208_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n205_), .A2(new_n218_), .ZN(new_n219_));
  NOR3_X1   g018(.A1(new_n214_), .A2(new_n215_), .A3(KEYINPUT8), .ZN(new_n220_));
  AOI22_X1  g019(.A1(new_n217_), .A2(KEYINPUT8), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT10), .B(G99gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n218_), .B1(G106gat), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT65), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT9), .B1(new_n214_), .B2(new_n215_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G85gat), .A2(G92gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT9), .ZN(new_n228_));
  AOI21_X1  g027(.A(KEYINPUT64), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n226_), .A2(new_n229_), .ZN(new_n230_));
  AND4_X1   g029(.A1(KEYINPUT64), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n225_), .B1(new_n230_), .B2(new_n232_), .ZN(new_n233_));
  AOI211_X1 g032(.A(KEYINPUT65), .B(new_n231_), .C1(new_n226_), .C2(new_n229_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n224_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(KEYINPUT66), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n237_));
  OAI211_X1 g036(.A(new_n237_), .B(new_n224_), .C1(new_n233_), .C2(new_n234_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n221_), .B1(new_n236_), .B2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G57gat), .B(G64gat), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n240_), .A2(KEYINPUT11), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n240_), .A2(KEYINPUT11), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G71gat), .B(G78gat), .ZN(new_n243_));
  OR3_X1    g042(.A1(new_n241_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n240_), .A2(new_n243_), .A3(KEYINPUT11), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n203_), .B1(new_n239_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT12), .ZN(new_n248_));
  INV_X1    g047(.A(new_n221_), .ZN(new_n249_));
  INV_X1    g048(.A(G85gat), .ZN(new_n250_));
  INV_X1    g049(.A(G92gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n228_), .B1(new_n252_), .B2(new_n227_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT64), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n254_), .B1(new_n214_), .B2(KEYINPUT9), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n232_), .B1(new_n253_), .B2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT65), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n230_), .A2(new_n225_), .A3(new_n232_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n237_), .B1(new_n259_), .B2(new_n224_), .ZN(new_n260_));
  AOI211_X1 g059(.A(KEYINPUT66), .B(new_n223_), .C1(new_n257_), .C2(new_n258_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n249_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n246_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n248_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  NOR3_X1   g063(.A1(new_n239_), .A2(KEYINPUT12), .A3(new_n246_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n247_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT68), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  OAI211_X1 g067(.A(new_n249_), .B(new_n246_), .C1(new_n260_), .C2(new_n261_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n239_), .A2(new_n246_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n203_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n262_), .A2(new_n248_), .A3(new_n263_), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT12), .B1(new_n239_), .B2(new_n246_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n275_), .A2(KEYINPUT68), .A3(new_n247_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G120gat), .B(G148gat), .ZN(new_n277_));
  INV_X1    g076(.A(G204gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  XOR2_X1   g078(.A(KEYINPUT5), .B(G176gat), .Z(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n268_), .A2(new_n272_), .A3(new_n276_), .A4(new_n281_), .ZN(new_n282_));
  AND3_X1   g081(.A1(new_n268_), .A2(new_n272_), .A3(new_n276_), .ZN(new_n283_));
  XOR2_X1   g082(.A(new_n281_), .B(KEYINPUT69), .Z(new_n284_));
  OAI21_X1  g083(.A(new_n282_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(KEYINPUT13), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT13), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n287_), .B(new_n282_), .C1(new_n283_), .C2(new_n284_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(G8gat), .ZN(new_n290_));
  INV_X1    g089(.A(G1gat), .ZN(new_n291_));
  XOR2_X1   g090(.A(KEYINPUT74), .B(G1gat), .Z(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT14), .B1(new_n292_), .B2(new_n290_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(KEYINPUT75), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT14), .ZN(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT74), .B(G1gat), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n295_), .B1(new_n296_), .B2(G8gat), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT75), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n294_), .A2(new_n299_), .ZN(new_n300_));
  XOR2_X1   g099(.A(G15gat), .B(G22gat), .Z(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n291_), .B1(new_n300_), .B2(new_n302_), .ZN(new_n303_));
  AOI211_X1 g102(.A(G1gat), .B(new_n301_), .C1(new_n294_), .C2(new_n299_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n290_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n299_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n297_), .A2(new_n298_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n302_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(G1gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n300_), .A2(new_n291_), .A3(new_n302_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n309_), .A2(G8gat), .A3(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n305_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G231gat), .A2(G233gat), .ZN(new_n313_));
  XOR2_X1   g112(.A(new_n313_), .B(KEYINPUT76), .Z(new_n314_));
  XOR2_X1   g113(.A(new_n246_), .B(new_n314_), .Z(new_n315_));
  XNOR2_X1  g114(.A(new_n312_), .B(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT17), .ZN(new_n317_));
  XNOR2_X1  g116(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G127gat), .B(G155gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G183gat), .B(G211gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  OR3_X1    g121(.A1(new_n316_), .A2(new_n317_), .A3(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(KEYINPUT17), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n316_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n323_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G190gat), .B(G218gat), .ZN(new_n328_));
  INV_X1    g127(.A(G134gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT72), .ZN(new_n331_));
  INV_X1    g130(.A(G162gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT36), .ZN(new_n334_));
  INV_X1    g133(.A(G36gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(G29gat), .ZN(new_n336_));
  INV_X1    g135(.A(G29gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(G36gat), .ZN(new_n338_));
  INV_X1    g137(.A(G43gat), .ZN(new_n339_));
  AND3_X1   g138(.A1(new_n336_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n339_), .B1(new_n336_), .B2(new_n338_), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT70), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n336_), .A2(new_n338_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(G43gat), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT70), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n336_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n344_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n347_));
  AND3_X1   g146(.A1(new_n342_), .A2(new_n347_), .A3(G50gat), .ZN(new_n348_));
  AOI21_X1  g147(.A(G50gat), .B1(new_n342_), .B2(new_n347_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT15), .ZN(new_n350_));
  NOR3_X1   g149(.A1(new_n348_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n342_), .A2(new_n347_), .ZN(new_n352_));
  INV_X1    g151(.A(G50gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n342_), .A2(new_n347_), .A3(G50gat), .ZN(new_n355_));
  AOI21_X1  g154(.A(KEYINPUT15), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n351_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT35), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G232gat), .A2(G233gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT34), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  AOI22_X1  g160(.A1(new_n357_), .A2(new_n262_), .B1(new_n358_), .B2(new_n361_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n348_), .A2(new_n349_), .ZN(new_n363_));
  NOR3_X1   g162(.A1(new_n262_), .A2(KEYINPUT71), .A3(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT71), .ZN(new_n365_));
  INV_X1    g164(.A(new_n363_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n365_), .B1(new_n239_), .B2(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n362_), .B1(new_n364_), .B2(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n361_), .A2(new_n358_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n369_), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n362_), .B(new_n371_), .C1(new_n364_), .C2(new_n367_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n334_), .B1(new_n370_), .B2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n370_), .A2(KEYINPUT73), .A3(new_n372_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n333_), .A2(KEYINPUT36), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n370_), .A2(KEYINPUT73), .A3(new_n372_), .A4(new_n375_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n373_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n379_), .A2(KEYINPUT37), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT37), .ZN(new_n381_));
  AOI211_X1 g180(.A(new_n381_), .B(new_n373_), .C1(new_n377_), .C2(new_n378_), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n289_), .B(new_n327_), .C1(new_n380_), .C2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G155gat), .A2(G162gat), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(G155gat), .A2(G162gat), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(G141gat), .ZN(new_n388_));
  INV_X1    g187(.A(G148gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT87), .ZN(new_n391_));
  NOR3_X1   g190(.A1(new_n390_), .A2(new_n391_), .A3(KEYINPUT3), .ZN(new_n392_));
  NOR3_X1   g191(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n393_), .A2(KEYINPUT87), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n392_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G141gat), .A2(G148gat), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT2), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n390_), .A2(KEYINPUT3), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT2), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n396_), .A2(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n398_), .A2(new_n399_), .A3(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n387_), .B1(new_n395_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT1), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n386_), .B1(new_n385_), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n384_), .A2(KEYINPUT1), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT86), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(KEYINPUT86), .B1(new_n384_), .B2(KEYINPUT1), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n405_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n390_), .A2(new_n396_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n410_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n403_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT4), .ZN(new_n415_));
  INV_X1    g214(.A(G120gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(G113gat), .ZN(new_n417_));
  INV_X1    g216(.A(G113gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(G120gat), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT85), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n417_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n420_), .B1(new_n417_), .B2(new_n419_), .ZN(new_n423_));
  OAI21_X1  g222(.A(G127gat), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n417_), .A2(new_n419_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(KEYINPUT85), .ZN(new_n426_));
  INV_X1    g225(.A(G127gat), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n426_), .A2(new_n427_), .A3(new_n421_), .ZN(new_n428_));
  AND3_X1   g227(.A1(new_n424_), .A2(new_n428_), .A3(G134gat), .ZN(new_n429_));
  AOI21_X1  g228(.A(G134gat), .B1(new_n424_), .B2(new_n428_), .ZN(new_n430_));
  OAI211_X1 g229(.A(new_n414_), .B(new_n415_), .C1(new_n429_), .C2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT97), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n414_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n434_));
  AOI22_X1  g233(.A1(new_n397_), .A2(KEYINPUT2), .B1(new_n390_), .B2(KEYINPUT3), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n435_), .B(new_n401_), .C1(new_n394_), .C2(new_n392_), .ZN(new_n436_));
  AOI22_X1  g235(.A1(new_n436_), .A2(new_n387_), .B1(new_n410_), .B2(new_n412_), .ZN(new_n437_));
  NOR3_X1   g236(.A1(new_n422_), .A2(new_n423_), .A3(G127gat), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n427_), .B1(new_n426_), .B2(new_n421_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n329_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n424_), .A2(new_n428_), .A3(G134gat), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n437_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n434_), .A2(KEYINPUT4), .A3(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G225gat), .A2(G233gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n440_), .A2(new_n441_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n445_), .A2(KEYINPUT97), .A3(new_n415_), .A4(new_n414_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n433_), .A2(new_n443_), .A3(new_n444_), .A4(new_n446_), .ZN(new_n447_));
  OR2_X1    g246(.A1(new_n447_), .A2(KEYINPUT100), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(KEYINPUT100), .ZN(new_n449_));
  INV_X1    g248(.A(new_n444_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n434_), .A2(new_n450_), .A3(new_n442_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G1gat), .B(G29gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n452_), .B(KEYINPUT0), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(G57gat), .ZN(new_n454_));
  OR2_X1    g253(.A1(new_n452_), .A2(KEYINPUT0), .ZN(new_n455_));
  INV_X1    g254(.A(G57gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n452_), .A2(KEYINPUT0), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n455_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  AND3_X1   g257(.A1(new_n454_), .A2(new_n458_), .A3(G85gat), .ZN(new_n459_));
  AOI21_X1  g258(.A(G85gat), .B1(new_n454_), .B2(new_n458_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  AND3_X1   g260(.A1(new_n451_), .A2(KEYINPUT99), .A3(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(KEYINPUT99), .B1(new_n451_), .B2(new_n461_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n448_), .A2(new_n449_), .A3(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G226gat), .A2(G233gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(KEYINPUT19), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT20), .ZN(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT25), .B(G183gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(KEYINPUT26), .B(G190gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  OR2_X1    g271(.A1(G169gat), .A2(G176gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G169gat), .A2(G176gat), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n473_), .A2(KEYINPUT24), .A3(new_n474_), .ZN(new_n475_));
  OR2_X1    g274(.A1(new_n473_), .A2(KEYINPUT24), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n472_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G183gat), .A2(G190gat), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT83), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(KEYINPUT83), .A2(G183gat), .A3(G190gat), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n480_), .A2(KEYINPUT23), .A3(new_n481_), .ZN(new_n482_));
  OR2_X1    g281(.A1(KEYINPUT82), .A2(KEYINPUT23), .ZN(new_n483_));
  NAND2_X1  g282(.A1(KEYINPUT82), .A2(KEYINPUT23), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n482_), .B1(new_n478_), .B2(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(KEYINPUT23), .B1(new_n480_), .B2(new_n481_), .ZN(new_n487_));
  AOI22_X1  g286(.A1(new_n483_), .A2(new_n484_), .B1(G183gat), .B2(G190gat), .ZN(new_n488_));
  OAI22_X1  g287(.A1(new_n487_), .A2(new_n488_), .B1(G183gat), .B2(G190gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT22), .B(G169gat), .ZN(new_n490_));
  INV_X1    g289(.A(G176gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n492_), .A2(new_n474_), .ZN(new_n493_));
  AOI22_X1  g292(.A1(new_n477_), .A2(new_n486_), .B1(new_n489_), .B2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G197gat), .B(G204gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(KEYINPUT90), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT21), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G211gat), .B(G218gat), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n496_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  XOR2_X1   g298(.A(G211gat), .B(G218gat), .Z(new_n500_));
  AOI21_X1  g299(.A(new_n500_), .B1(KEYINPUT90), .B2(new_n495_), .ZN(new_n501_));
  XOR2_X1   g300(.A(G197gat), .B(G204gat), .Z(new_n502_));
  OAI21_X1  g301(.A(KEYINPUT21), .B1(new_n502_), .B2(new_n498_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n499_), .B1(new_n501_), .B2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n469_), .B1(new_n494_), .B2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(KEYINPUT91), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT91), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n508_), .B(new_n499_), .C1(new_n501_), .C2(new_n503_), .ZN(new_n509_));
  AND2_X1   g308(.A1(new_n507_), .A2(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n476_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT80), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n470_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT25), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n512_), .B1(new_n514_), .B2(G183gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n471_), .A2(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n475_), .B1(new_n513_), .B2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT81), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n511_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  OAI211_X1 g318(.A(KEYINPUT81), .B(new_n475_), .C1(new_n513_), .C2(new_n516_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n486_), .B1(G183gat), .B2(G190gat), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT84), .ZN(new_n522_));
  AOI21_X1  g321(.A(G176gat), .B1(new_n522_), .B2(KEYINPUT22), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(G169gat), .ZN(new_n524_));
  AOI22_X1  g323(.A1(new_n519_), .A2(new_n520_), .B1(new_n521_), .B2(new_n524_), .ZN(new_n525_));
  OAI211_X1 g324(.A(new_n468_), .B(new_n506_), .C1(new_n510_), .C2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT94), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n519_), .A2(new_n520_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n521_), .A2(new_n524_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n507_), .A2(new_n509_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT94), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n532_), .A2(new_n533_), .A3(new_n468_), .A4(new_n506_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n477_), .A2(new_n486_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n489_), .A2(new_n493_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n469_), .B1(new_n537_), .B2(new_n504_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n538_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(new_n467_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G64gat), .B(G92gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G8gat), .B(G36gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT96), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n543_), .B(new_n545_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n527_), .A2(new_n534_), .A3(new_n540_), .A4(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n527_), .A2(new_n534_), .A3(new_n540_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n546_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  AND3_X1   g349(.A1(new_n465_), .A2(new_n547_), .A3(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT98), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n552_), .A2(KEYINPUT33), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n450_), .B1(new_n434_), .B2(new_n442_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n433_), .A2(new_n443_), .A3(new_n446_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n555_), .B1(new_n556_), .B2(new_n450_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n461_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n554_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  NOR3_X1   g359(.A1(new_n557_), .A2(new_n461_), .A3(new_n553_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n551_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n557_), .A2(new_n461_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT102), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n557_), .A2(KEYINPUT102), .A3(new_n461_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n558_), .A2(new_n559_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n566_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n546_), .A2(KEYINPUT32), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n548_), .A2(new_n571_), .ZN(new_n572_));
  AOI22_X1  g371(.A1(new_n528_), .A2(new_n529_), .B1(new_n507_), .B2(new_n509_), .ZN(new_n573_));
  OAI21_X1  g372(.A(KEYINPUT20), .B1(new_n537_), .B2(new_n504_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n467_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(KEYINPUT20), .B1(new_n494_), .B2(new_n505_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n576_), .B1(new_n510_), .B2(new_n525_), .ZN(new_n577_));
  AOI22_X1  g376(.A1(new_n575_), .A2(KEYINPUT101), .B1(new_n577_), .B2(new_n468_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n468_), .B1(new_n532_), .B2(new_n506_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT101), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n570_), .B1(new_n578_), .B2(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n572_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n569_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n563_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G228gat), .A2(G233gat), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n586_), .B(KEYINPUT89), .Z(new_n587_));
  INV_X1    g386(.A(new_n387_), .ZN(new_n588_));
  AND3_X1   g387(.A1(new_n398_), .A2(new_n399_), .A3(new_n401_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n393_), .B(KEYINPUT87), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n588_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n406_), .B(new_n407_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n411_), .B1(new_n592_), .B2(new_n405_), .ZN(new_n593_));
  OAI21_X1  g392(.A(KEYINPUT29), .B1(new_n591_), .B2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n531_), .A2(new_n587_), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT92), .ZN(new_n596_));
  AOI211_X1 g395(.A(new_n596_), .B(new_n587_), .C1(new_n594_), .C2(new_n504_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT29), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n504_), .B1(new_n437_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n587_), .ZN(new_n600_));
  AOI21_X1  g399(.A(KEYINPUT92), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n595_), .B1(new_n597_), .B2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G78gat), .B(G106gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT93), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n606_), .B1(new_n414_), .B2(KEYINPUT29), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G22gat), .B(G50gat), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n606_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n437_), .A2(new_n598_), .A3(new_n610_), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n607_), .A2(new_n609_), .A3(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n609_), .B1(new_n607_), .B2(new_n611_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n604_), .ZN(new_n615_));
  OAI211_X1 g414(.A(new_n615_), .B(new_n595_), .C1(new_n597_), .C2(new_n601_), .ZN(new_n616_));
  AND3_X1   g415(.A1(new_n605_), .A2(new_n614_), .A3(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n614_), .B1(new_n605_), .B2(new_n616_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT31), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n445_), .A2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n440_), .A2(KEYINPUT31), .A3(new_n441_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(G227gat), .A2(G233gat), .ZN(new_n623_));
  AND3_X1   g422(.A1(new_n621_), .A2(new_n622_), .A3(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n623_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G15gat), .B(G43gat), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  AND3_X1   g428(.A1(new_n528_), .A2(KEYINPUT30), .A3(new_n529_), .ZN(new_n630_));
  AOI21_X1  g429(.A(KEYINPUT30), .B1(new_n528_), .B2(new_n529_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n629_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT30), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n530_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n525_), .A2(KEYINPUT30), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n634_), .A2(new_n635_), .A3(new_n628_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(G71gat), .B(G99gat), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  AND3_X1   g437(.A1(new_n632_), .A2(new_n636_), .A3(new_n638_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n638_), .B1(new_n632_), .B2(new_n636_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n627_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n630_), .A2(new_n631_), .A3(new_n629_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n628_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n637_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n632_), .A2(new_n636_), .A3(new_n638_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n644_), .A2(new_n626_), .A3(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n641_), .A2(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n619_), .A2(new_n647_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n639_), .A2(new_n640_), .A3(new_n627_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n626_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n650_));
  OAI22_X1  g449(.A1(new_n649_), .A2(new_n650_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n614_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n599_), .A2(new_n600_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(new_n596_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n599_), .A2(KEYINPUT92), .A3(new_n600_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n615_), .B1(new_n656_), .B2(new_n595_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n616_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n652_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n605_), .A2(new_n614_), .A3(new_n616_), .ZN(new_n660_));
  NAND4_X1  g459(.A1(new_n641_), .A2(new_n659_), .A3(new_n646_), .A4(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n569_), .B1(new_n651_), .B2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n547_), .A2(KEYINPUT27), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n546_), .B1(new_n578_), .B2(new_n581_), .ZN(new_n664_));
  OAI21_X1  g463(.A(KEYINPUT103), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  OAI211_X1 g464(.A(new_n538_), .B(new_n468_), .C1(new_n530_), .C2(new_n531_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n666_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n575_), .A2(KEYINPUT101), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n549_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT103), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n669_), .A2(new_n670_), .A3(KEYINPUT27), .A4(new_n547_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT27), .ZN(new_n672_));
  INV_X1    g471(.A(new_n547_), .ZN(new_n673_));
  AOI22_X1  g472(.A1(new_n526_), .A2(KEYINPUT94), .B1(new_n539_), .B2(new_n467_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n546_), .B1(new_n674_), .B2(new_n534_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n672_), .B1(new_n673_), .B2(new_n675_), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n665_), .A2(new_n671_), .A3(new_n676_), .ZN(new_n677_));
  AOI22_X1  g476(.A1(new_n585_), .A2(new_n648_), .B1(new_n662_), .B2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(G229gat), .A2(G233gat), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n305_), .A2(new_n311_), .A3(new_n363_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n363_), .B1(new_n305_), .B2(new_n311_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n680_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n312_), .A2(new_n366_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n357_), .A2(new_n311_), .A3(new_n305_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n684_), .A2(new_n679_), .A3(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n683_), .A2(new_n686_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(G113gat), .B(G141gat), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(G169gat), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n689_), .B(G197gat), .Z(new_n690_));
  NAND3_X1  g489(.A1(new_n687_), .A2(KEYINPUT78), .A3(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n690_), .B1(new_n687_), .B2(KEYINPUT78), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n692_), .A2(new_n693_), .A3(KEYINPUT79), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT79), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n687_), .A2(KEYINPUT78), .ZN(new_n696_));
  INV_X1    g495(.A(new_n690_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n695_), .B1(new_n698_), .B2(new_n691_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n694_), .A2(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(KEYINPUT104), .B1(new_n678_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n569_), .ZN(new_n702_));
  AND4_X1   g501(.A1(new_n660_), .A2(new_n641_), .A3(new_n659_), .A4(new_n646_), .ZN(new_n703_));
  AOI22_X1  g502(.A1(new_n646_), .A2(new_n641_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n702_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n665_), .A2(new_n671_), .A3(new_n676_), .ZN(new_n706_));
  AOI22_X1  g505(.A1(new_n551_), .A2(new_n562_), .B1(new_n569_), .B2(new_n583_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n648_), .ZN(new_n708_));
  OAI22_X1  g507(.A1(new_n705_), .A2(new_n706_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n700_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT104), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n709_), .A2(new_n710_), .A3(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n383_), .B1(new_n701_), .B2(new_n712_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n569_), .B(KEYINPUT105), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n713_), .A2(new_n292_), .A3(new_n715_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT38), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n709_), .A2(new_n379_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT106), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n692_), .A2(new_n693_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n289_), .A2(new_n720_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n721_), .A2(new_n326_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n719_), .A2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT107), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n723_), .B(new_n724_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n725_), .A2(new_n569_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n717_), .B1(new_n726_), .B2(new_n291_), .ZN(G1324gat));
  NAND3_X1  g526(.A1(new_n719_), .A2(new_n706_), .A3(new_n722_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT108), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n728_), .A2(new_n729_), .A3(G8gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n728_), .B2(G8gat), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT39), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n730_), .A2(new_n731_), .A3(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n732_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n713_), .A2(new_n290_), .A3(new_n706_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT40), .ZN(new_n737_));
  OR3_X1    g536(.A1(new_n733_), .A2(new_n736_), .A3(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n737_), .B1(new_n733_), .B2(new_n736_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(G1325gat));
  INV_X1    g539(.A(G15gat), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n713_), .A2(new_n741_), .A3(new_n647_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n725_), .A2(new_n647_), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n743_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n744_));
  AOI21_X1  g543(.A(KEYINPUT41), .B1(new_n743_), .B2(G15gat), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n742_), .B1(new_n744_), .B2(new_n745_), .ZN(G1326gat));
  INV_X1    g545(.A(G22gat), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n713_), .A2(new_n747_), .A3(new_n619_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT42), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n725_), .A2(new_n619_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n750_), .B2(G22gat), .ZN(new_n751_));
  AOI211_X1 g550(.A(KEYINPUT42), .B(new_n747_), .C1(new_n725_), .C2(new_n619_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n748_), .B1(new_n751_), .B2(new_n752_), .ZN(G1327gat));
  NAND2_X1  g552(.A1(new_n377_), .A2(new_n378_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n373_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n756_), .A2(new_n326_), .A3(KEYINPUT110), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT110), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n758_), .B1(new_n379_), .B2(new_n327_), .ZN(new_n759_));
  AOI22_X1  g558(.A1(new_n757_), .A2(new_n759_), .B1(new_n286_), .B2(new_n288_), .ZN(new_n760_));
  NOR3_X1   g559(.A1(new_n678_), .A2(KEYINPUT104), .A3(new_n700_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n711_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n762_));
  OAI211_X1 g561(.A(KEYINPUT111), .B(new_n760_), .C1(new_n761_), .C2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n701_), .A2(new_n712_), .ZN(new_n765_));
  AOI21_X1  g564(.A(KEYINPUT111), .B1(new_n765_), .B2(new_n760_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n764_), .A2(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(G29gat), .B1(new_n767_), .B2(new_n569_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n289_), .A2(new_n326_), .A3(new_n720_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n756_), .A2(new_n381_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n379_), .A2(KEYINPUT37), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n770_), .A2(new_n771_), .A3(KEYINPUT109), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n771_), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n772_), .B(KEYINPUT43), .C1(new_n773_), .C2(new_n678_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n380_), .A2(new_n382_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT43), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n775_), .B(new_n709_), .C1(KEYINPUT109), .C2(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n769_), .B1(new_n774_), .B2(new_n777_), .ZN(new_n778_));
  AOI211_X1 g577(.A(new_n337_), .B(new_n714_), .C1(new_n778_), .C2(KEYINPUT44), .ZN(new_n779_));
  INV_X1    g578(.A(new_n778_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT44), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n768_), .B1(new_n779_), .B2(new_n782_), .ZN(G1328gat));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT113), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n677_), .A2(G36gat), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n785_), .B1(new_n767_), .B2(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n760_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT111), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n790_), .A2(new_n763_), .A3(new_n786_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n791_), .A2(KEYINPUT113), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n784_), .B1(new_n787_), .B2(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n767_), .A2(new_n785_), .A3(new_n786_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n791_), .A2(KEYINPUT113), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n794_), .A2(KEYINPUT45), .A3(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n677_), .B1(new_n778_), .B2(KEYINPUT44), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n335_), .B1(new_n782_), .B2(new_n797_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n798_), .A2(KEYINPUT112), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT112), .ZN(new_n800_));
  AOI211_X1 g599(.A(new_n800_), .B(new_n335_), .C1(new_n782_), .C2(new_n797_), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n793_), .B(new_n796_), .C1(new_n799_), .C2(new_n801_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(KEYINPUT114), .A2(KEYINPUT46), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n798_), .B(KEYINPUT112), .ZN(new_n805_));
  INV_X1    g604(.A(new_n803_), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n805_), .A2(new_n806_), .A3(new_n796_), .A4(new_n793_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n804_), .A2(new_n807_), .ZN(G1329gat));
  INV_X1    g607(.A(KEYINPUT47), .ZN(new_n809_));
  INV_X1    g608(.A(new_n767_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n647_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n339_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT115), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n778_), .A2(KEYINPUT44), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n782_), .A2(G43gat), .A3(new_n647_), .A4(new_n814_), .ZN(new_n815_));
  AND3_X1   g614(.A1(new_n812_), .A2(new_n813_), .A3(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n813_), .B1(new_n812_), .B2(new_n815_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n809_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n812_), .A2(new_n815_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT115), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n812_), .A2(new_n813_), .A3(new_n815_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n820_), .A2(KEYINPUT47), .A3(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n818_), .A2(new_n822_), .ZN(G1330gat));
  NAND3_X1  g622(.A1(new_n782_), .A2(new_n619_), .A3(new_n814_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(G50gat), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n619_), .A2(new_n353_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n826_), .B(KEYINPUT116), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n825_), .B1(new_n810_), .B2(new_n827_), .ZN(G1331gat));
  INV_X1    g627(.A(new_n289_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n719_), .A2(new_n327_), .A3(new_n829_), .A4(new_n700_), .ZN(new_n830_));
  OAI21_X1  g629(.A(G57gat), .B1(new_n830_), .B2(new_n702_), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n678_), .A2(new_n720_), .A3(new_n289_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n326_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n715_), .A2(new_n456_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n831_), .B1(new_n834_), .B2(new_n835_), .ZN(G1332gat));
  OAI21_X1  g635(.A(G64gat), .B1(new_n830_), .B2(new_n677_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(KEYINPUT48), .ZN(new_n838_));
  OR2_X1    g637(.A1(new_n677_), .A2(G64gat), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n838_), .B1(new_n834_), .B2(new_n839_), .ZN(G1333gat));
  OAI21_X1  g639(.A(G71gat), .B1(new_n830_), .B2(new_n811_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(KEYINPUT49), .ZN(new_n842_));
  OR2_X1    g641(.A1(new_n811_), .A2(G71gat), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n834_), .B2(new_n843_), .ZN(G1334gat));
  INV_X1    g643(.A(new_n619_), .ZN(new_n845_));
  OAI21_X1  g644(.A(G78gat), .B1(new_n830_), .B2(new_n845_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(KEYINPUT50), .ZN(new_n847_));
  OR2_X1    g646(.A1(new_n845_), .A2(G78gat), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n847_), .B1(new_n834_), .B2(new_n848_), .ZN(G1335gat));
  NAND2_X1  g648(.A1(new_n774_), .A2(new_n777_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n720_), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n850_), .A2(new_n326_), .A3(new_n851_), .A4(new_n829_), .ZN(new_n852_));
  OAI21_X1  g651(.A(G85gat), .B1(new_n852_), .B2(new_n702_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n757_), .A2(new_n759_), .ZN(new_n854_));
  AND2_X1   g653(.A1(new_n832_), .A2(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n855_), .A2(new_n250_), .A3(new_n715_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n853_), .A2(new_n856_), .ZN(G1336gat));
  AOI21_X1  g656(.A(G92gat), .B1(new_n855_), .B2(new_n706_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(KEYINPUT117), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n852_), .A2(new_n251_), .A3(new_n677_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n859_), .A2(new_n860_), .ZN(G1337gat));
  NOR2_X1   g660(.A1(new_n811_), .A2(new_n222_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n855_), .A2(new_n862_), .ZN(new_n863_));
  XOR2_X1   g662(.A(new_n863_), .B(KEYINPUT118), .Z(new_n864_));
  OAI21_X1  g663(.A(G99gat), .B1(new_n852_), .B2(new_n811_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g666(.A(G106gat), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n855_), .A2(new_n868_), .A3(new_n619_), .ZN(new_n869_));
  OR2_X1    g668(.A1(new_n852_), .A2(new_n845_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT52), .ZN(new_n871_));
  AND3_X1   g670(.A1(new_n870_), .A2(new_n871_), .A3(G106gat), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n871_), .B1(new_n870_), .B2(G106gat), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n869_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(KEYINPUT53), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT53), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n876_), .B(new_n869_), .C1(new_n872_), .C2(new_n873_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n875_), .A2(new_n877_), .ZN(G1339gat));
  OAI21_X1  g677(.A(KEYINPUT54), .B1(new_n383_), .B2(new_n710_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT54), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n833_), .A2(new_n880_), .A3(new_n289_), .A4(new_n700_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n687_), .A2(new_n690_), .ZN(new_n884_));
  AND3_X1   g683(.A1(new_n684_), .A2(new_n680_), .A3(new_n685_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n305_), .A2(new_n311_), .A3(new_n363_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n680_), .B1(new_n684_), .B2(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n697_), .B1(new_n885_), .B2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n884_), .A2(new_n888_), .ZN(new_n889_));
  AND2_X1   g688(.A1(new_n889_), .A2(new_n282_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT55), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n268_), .A2(new_n891_), .A3(new_n276_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n275_), .A2(new_n269_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n269_), .A2(new_n202_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n894_), .B1(new_n274_), .B2(new_n273_), .ZN(new_n895_));
  AOI22_X1  g694(.A1(new_n893_), .A2(new_n203_), .B1(new_n895_), .B2(KEYINPUT55), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n892_), .A2(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n284_), .ZN(new_n898_));
  AOI21_X1  g697(.A(KEYINPUT56), .B1(new_n897_), .B2(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT56), .ZN(new_n900_));
  AOI211_X1 g699(.A(new_n900_), .B(new_n284_), .C1(new_n892_), .C2(new_n896_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n890_), .B1(new_n899_), .B2(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT58), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  OAI211_X1 g703(.A(KEYINPUT58), .B(new_n890_), .C1(new_n899_), .C2(new_n901_), .ZN(new_n905_));
  AND3_X1   g704(.A1(new_n904_), .A2(new_n775_), .A3(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n906_), .ZN(new_n907_));
  AND3_X1   g706(.A1(new_n698_), .A2(new_n691_), .A3(new_n282_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n908_), .B1(new_n899_), .B2(new_n901_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT119), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  OAI211_X1 g710(.A(new_n908_), .B(KEYINPUT119), .C1(new_n899_), .C2(new_n901_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n285_), .A2(new_n889_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n911_), .A2(new_n912_), .A3(new_n913_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n914_), .A2(KEYINPUT57), .A3(new_n379_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n913_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n916_), .B1(new_n909_), .B2(new_n910_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n756_), .B1(new_n917_), .B2(new_n912_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n919_));
  OAI211_X1 g718(.A(new_n907_), .B(new_n915_), .C1(new_n918_), .C2(new_n919_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n883_), .B1(new_n920_), .B2(new_n326_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n921_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT59), .ZN(new_n923_));
  NOR3_X1   g722(.A1(new_n714_), .A2(new_n706_), .A3(new_n651_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n923_), .B1(new_n924_), .B2(KEYINPUT122), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n925_), .B1(KEYINPUT122), .B2(new_n924_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n922_), .A2(new_n926_), .ZN(new_n927_));
  INV_X1    g726(.A(new_n924_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n906_), .B1(new_n918_), .B2(KEYINPUT57), .ZN(new_n929_));
  OAI21_X1  g728(.A(KEYINPUT121), .B1(new_n918_), .B2(new_n919_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n929_), .A2(new_n930_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n914_), .A2(new_n379_), .ZN(new_n932_));
  INV_X1    g731(.A(new_n919_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n934_), .A2(KEYINPUT121), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n326_), .B1(new_n931_), .B2(new_n935_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n928_), .B1(new_n936_), .B2(new_n882_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n927_), .B1(new_n937_), .B2(new_n923_), .ZN(new_n938_));
  OAI21_X1  g737(.A(G113gat), .B1(new_n938_), .B2(new_n700_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n937_), .A2(new_n418_), .A3(new_n720_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n939_), .A2(new_n940_), .ZN(G1340gat));
  XNOR2_X1  g740(.A(KEYINPUT123), .B(G120gat), .ZN(new_n942_));
  INV_X1    g741(.A(new_n942_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n943_), .B1(new_n938_), .B2(new_n289_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n942_), .B1(new_n289_), .B2(KEYINPUT60), .ZN(new_n945_));
  OAI211_X1 g744(.A(new_n937_), .B(new_n945_), .C1(KEYINPUT60), .C2(new_n942_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n944_), .A2(new_n946_), .ZN(G1341gat));
  OAI21_X1  g746(.A(G127gat), .B1(new_n938_), .B2(new_n326_), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n937_), .A2(new_n427_), .A3(new_n327_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n948_), .A2(new_n949_), .ZN(G1342gat));
  OAI21_X1  g749(.A(G134gat), .B1(new_n938_), .B2(new_n773_), .ZN(new_n951_));
  NAND3_X1  g750(.A1(new_n937_), .A2(new_n329_), .A3(new_n756_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n951_), .A2(new_n952_), .ZN(G1343gat));
  NAND2_X1  g752(.A1(new_n936_), .A2(new_n882_), .ZN(new_n954_));
  NOR3_X1   g753(.A1(new_n714_), .A2(new_n706_), .A3(new_n661_), .ZN(new_n955_));
  XNOR2_X1  g754(.A(new_n955_), .B(KEYINPUT124), .ZN(new_n956_));
  NAND3_X1  g755(.A1(new_n954_), .A2(new_n720_), .A3(new_n956_), .ZN(new_n957_));
  XNOR2_X1  g756(.A(new_n957_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g757(.A1(new_n954_), .A2(new_n829_), .A3(new_n956_), .ZN(new_n959_));
  XNOR2_X1  g758(.A(new_n959_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g759(.A1(new_n954_), .A2(new_n327_), .A3(new_n956_), .ZN(new_n961_));
  XNOR2_X1  g760(.A(KEYINPUT61), .B(G155gat), .ZN(new_n962_));
  XNOR2_X1  g761(.A(new_n961_), .B(new_n962_), .ZN(G1346gat));
  NAND4_X1  g762(.A1(new_n954_), .A2(new_n332_), .A3(new_n756_), .A4(new_n956_), .ZN(new_n964_));
  AND3_X1   g763(.A1(new_n954_), .A2(new_n775_), .A3(new_n956_), .ZN(new_n965_));
  OAI21_X1  g764(.A(new_n964_), .B1(new_n965_), .B2(new_n332_), .ZN(G1347gat));
  NOR2_X1   g765(.A1(new_n677_), .A2(new_n811_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n967_), .A2(new_n714_), .ZN(new_n968_));
  NOR2_X1   g767(.A1(new_n968_), .A2(new_n851_), .ZN(new_n969_));
  NAND4_X1  g768(.A1(new_n922_), .A2(new_n490_), .A3(new_n845_), .A4(new_n969_), .ZN(new_n970_));
  INV_X1    g769(.A(KEYINPUT62), .ZN(new_n971_));
  OR3_X1    g770(.A1(new_n968_), .A2(KEYINPUT125), .A3(new_n851_), .ZN(new_n972_));
  OAI21_X1  g771(.A(KEYINPUT125), .B1(new_n968_), .B2(new_n851_), .ZN(new_n973_));
  NAND3_X1  g772(.A1(new_n972_), .A2(new_n845_), .A3(new_n973_), .ZN(new_n974_));
  OAI211_X1 g773(.A(new_n971_), .B(G169gat), .C1(new_n921_), .C2(new_n974_), .ZN(new_n975_));
  INV_X1    g774(.A(new_n975_), .ZN(new_n976_));
  INV_X1    g775(.A(new_n974_), .ZN(new_n977_));
  AOI21_X1  g776(.A(new_n327_), .B1(new_n929_), .B2(new_n934_), .ZN(new_n978_));
  OAI21_X1  g777(.A(new_n977_), .B1(new_n978_), .B2(new_n883_), .ZN(new_n979_));
  AOI21_X1  g778(.A(new_n971_), .B1(new_n979_), .B2(G169gat), .ZN(new_n980_));
  OAI21_X1  g779(.A(new_n970_), .B1(new_n976_), .B2(new_n980_), .ZN(new_n981_));
  INV_X1    g780(.A(KEYINPUT126), .ZN(new_n982_));
  NAND2_X1  g781(.A1(new_n981_), .A2(new_n982_), .ZN(new_n983_));
  OAI211_X1 g782(.A(KEYINPUT126), .B(new_n970_), .C1(new_n976_), .C2(new_n980_), .ZN(new_n984_));
  NAND2_X1  g783(.A1(new_n983_), .A2(new_n984_), .ZN(G1348gat));
  OR3_X1    g784(.A1(new_n921_), .A2(new_n619_), .A3(new_n968_), .ZN(new_n986_));
  OAI211_X1 g785(.A(KEYINPUT127), .B(new_n491_), .C1(new_n986_), .C2(new_n289_), .ZN(new_n987_));
  INV_X1    g786(.A(KEYINPUT127), .ZN(new_n988_));
  NOR4_X1   g787(.A1(new_n921_), .A2(new_n619_), .A3(new_n289_), .A4(new_n968_), .ZN(new_n989_));
  OAI21_X1  g788(.A(new_n988_), .B1(new_n989_), .B2(G176gat), .ZN(new_n990_));
  AOI21_X1  g789(.A(new_n619_), .B1(new_n936_), .B2(new_n882_), .ZN(new_n991_));
  NOR3_X1   g790(.A1(new_n968_), .A2(new_n491_), .A3(new_n289_), .ZN(new_n992_));
  AOI22_X1  g791(.A1(new_n987_), .A2(new_n990_), .B1(new_n991_), .B2(new_n992_), .ZN(G1349gat));
  NOR2_X1   g792(.A1(new_n968_), .A2(new_n326_), .ZN(new_n994_));
  AOI21_X1  g793(.A(G183gat), .B1(new_n991_), .B2(new_n994_), .ZN(new_n995_));
  NOR2_X1   g794(.A1(new_n921_), .A2(new_n619_), .ZN(new_n996_));
  NOR3_X1   g795(.A1(new_n968_), .A2(new_n470_), .A3(new_n326_), .ZN(new_n997_));
  AOI21_X1  g796(.A(new_n995_), .B1(new_n996_), .B2(new_n997_), .ZN(G1350gat));
  OAI21_X1  g797(.A(G190gat), .B1(new_n986_), .B2(new_n773_), .ZN(new_n999_));
  NAND2_X1  g798(.A1(new_n756_), .A2(new_n471_), .ZN(new_n1000_));
  OAI21_X1  g799(.A(new_n999_), .B1(new_n986_), .B2(new_n1000_), .ZN(G1351gat));
  NOR3_X1   g800(.A1(new_n677_), .A2(new_n569_), .A3(new_n661_), .ZN(new_n1002_));
  NAND3_X1  g801(.A1(new_n954_), .A2(new_n720_), .A3(new_n1002_), .ZN(new_n1003_));
  XNOR2_X1  g802(.A(new_n1003_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g803(.A1(new_n954_), .A2(new_n1002_), .ZN(new_n1005_));
  INV_X1    g804(.A(new_n1005_), .ZN(new_n1006_));
  AOI21_X1  g805(.A(G204gat), .B1(new_n1006_), .B2(new_n829_), .ZN(new_n1007_));
  NOR3_X1   g806(.A1(new_n1005_), .A2(new_n278_), .A3(new_n289_), .ZN(new_n1008_));
  NOR2_X1   g807(.A1(new_n1007_), .A2(new_n1008_), .ZN(G1353gat));
  XNOR2_X1  g808(.A(KEYINPUT63), .B(G211gat), .ZN(new_n1010_));
  NOR3_X1   g809(.A1(new_n1005_), .A2(new_n326_), .A3(new_n1010_), .ZN(new_n1011_));
  NAND2_X1  g810(.A1(new_n1006_), .A2(new_n327_), .ZN(new_n1012_));
  NOR2_X1   g811(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1013_));
  AOI21_X1  g812(.A(new_n1011_), .B1(new_n1012_), .B2(new_n1013_), .ZN(G1354gat));
  OR3_X1    g813(.A1(new_n1005_), .A2(G218gat), .A3(new_n379_), .ZN(new_n1015_));
  OAI21_X1  g814(.A(G218gat), .B1(new_n1005_), .B2(new_n773_), .ZN(new_n1016_));
  NAND2_X1  g815(.A1(new_n1015_), .A2(new_n1016_), .ZN(G1355gat));
endmodule


