//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 1 1 1 1 1 1 0 1 1 0 1 1 1 0 0 1 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 0 1 1 0 1 1 0 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n754_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n769_, new_n770_, new_n771_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n778_, new_n779_, new_n780_, new_n781_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n790_,
    new_n791_, new_n793_, new_n794_, new_n795_, new_n796_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_, new_n902_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n909_, new_n911_, new_n912_, new_n913_,
    new_n915_, new_n916_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n937_, new_n938_, new_n939_, new_n941_, new_n942_,
    new_n944_, new_n945_, new_n947_, new_n948_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n956_, new_n957_;
  XOR2_X1   g000(.A(G57gat), .B(G64gat), .Z(new_n202_));
  INV_X1    g001(.A(KEYINPUT11), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  OR2_X1    g003(.A1(G71gat), .A2(G78gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G71gat), .A2(G78gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT67), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n202_), .A2(new_n203_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT6), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n211_), .B(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT9), .ZN(new_n214_));
  INV_X1    g013(.A(G85gat), .ZN(new_n215_));
  INV_X1    g014(.A(G92gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n214_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  XOR2_X1   g016(.A(G85gat), .B(G92gat), .Z(new_n218_));
  OAI21_X1  g017(.A(new_n217_), .B1(new_n218_), .B2(new_n214_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT64), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT64), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n221_), .B(new_n217_), .C1(new_n218_), .C2(new_n214_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n213_), .B1(new_n220_), .B2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT10), .B(G99gat), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n223_), .B1(G106gat), .B2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT8), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n211_), .B(KEYINPUT6), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT65), .B(KEYINPUT66), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n228_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n213_), .A2(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(G99gat), .A2(G106gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT7), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n229_), .A2(new_n231_), .A3(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n226_), .B1(new_n234_), .B2(new_n218_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n218_), .A2(new_n226_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n236_), .B1(new_n233_), .B2(new_n227_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n225_), .B1(new_n235_), .B2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n210_), .B(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G230gat), .A2(G233gat), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n235_), .A2(new_n237_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n224_), .A2(G106gat), .ZN(new_n244_));
  AOI211_X1 g043(.A(new_n213_), .B(new_n244_), .C1(new_n220_), .C2(new_n222_), .ZN(new_n245_));
  OAI211_X1 g044(.A(new_n242_), .B(KEYINPUT12), .C1(new_n243_), .C2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT12), .ZN(new_n247_));
  OAI211_X1 g046(.A(new_n225_), .B(new_n247_), .C1(new_n235_), .C2(new_n237_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n209_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n208_), .B(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n249_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n210_), .A2(new_n246_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n252_), .A2(new_n240_), .A3(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT69), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT69), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n252_), .A2(new_n256_), .A3(new_n240_), .A4(new_n253_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n241_), .B1(new_n255_), .B2(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G120gat), .B(G148gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G176gat), .B(G204gat), .ZN(new_n262_));
  XOR2_X1   g061(.A(new_n261_), .B(new_n262_), .Z(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  OR2_X1    g063(.A1(new_n258_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n258_), .A2(new_n264_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT71), .B(KEYINPUT13), .ZN(new_n268_));
  OR2_X1    g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT71), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n267_), .B1(new_n270_), .B2(KEYINPUT13), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT81), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G29gat), .B(G36gat), .ZN(new_n275_));
  INV_X1    g074(.A(G43gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(G50gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n275_), .B(G43gat), .ZN(new_n279_));
  INV_X1    g078(.A(G50gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n278_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT80), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n278_), .A2(new_n281_), .A3(KEYINPUT80), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT78), .ZN(new_n287_));
  XOR2_X1   g086(.A(G1gat), .B(G8gat), .Z(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G15gat), .B(G22gat), .ZN(new_n290_));
  INV_X1    g089(.A(G1gat), .ZN(new_n291_));
  INV_X1    g090(.A(G8gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT14), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n290_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n289_), .B(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT77), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n294_), .B(new_n288_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n298_), .A2(KEYINPUT77), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n287_), .B1(new_n297_), .B2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n295_), .A2(new_n296_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n298_), .A2(KEYINPUT77), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n301_), .A2(KEYINPUT78), .A3(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n286_), .A2(new_n300_), .A3(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n286_), .B1(new_n303_), .B2(new_n300_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n274_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n300_), .A2(new_n303_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n308_), .A2(new_n285_), .A3(new_n284_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n309_), .A2(KEYINPUT81), .A3(new_n304_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G229gat), .A2(G233gat), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n307_), .A2(new_n310_), .A3(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G113gat), .B(G141gat), .ZN(new_n314_));
  INV_X1    g113(.A(G169gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(G197gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(KEYINPUT82), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n308_), .ZN(new_n321_));
  XOR2_X1   g120(.A(new_n282_), .B(KEYINPUT15), .Z(new_n322_));
  AOI21_X1  g121(.A(new_n306_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(new_n311_), .ZN(new_n324_));
  AND3_X1   g123(.A1(new_n313_), .A2(new_n320_), .A3(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n320_), .B1(new_n313_), .B2(new_n324_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n273_), .A2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G78gat), .B(G106gat), .ZN(new_n330_));
  XOR2_X1   g129(.A(new_n330_), .B(KEYINPUT91), .Z(new_n331_));
  NAND2_X1  g130(.A1(G228gat), .A2(G233gat), .ZN(new_n332_));
  XOR2_X1   g131(.A(new_n332_), .B(KEYINPUT92), .Z(new_n333_));
  INV_X1    g132(.A(KEYINPUT29), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT90), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G155gat), .A2(G162gat), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT3), .ZN(new_n338_));
  INV_X1    g137(.A(G141gat), .ZN(new_n339_));
  INV_X1    g138(.A(G148gat), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n338_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G141gat), .A2(G148gat), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT2), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n345_));
  OAI21_X1  g144(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n341_), .A2(new_n344_), .A3(new_n345_), .A4(new_n346_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(G155gat), .A2(G162gat), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n347_), .A2(new_n349_), .ZN(new_n350_));
  XOR2_X1   g149(.A(G141gat), .B(G148gat), .Z(new_n351_));
  OR2_X1    g150(.A1(new_n348_), .A2(KEYINPUT1), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n337_), .B1(new_n350_), .B2(new_n353_), .ZN(new_n354_));
  OR3_X1    g153(.A1(new_n336_), .A2(KEYINPUT89), .A3(KEYINPUT1), .ZN(new_n355_));
  OAI21_X1  g154(.A(KEYINPUT89), .B1(new_n336_), .B2(KEYINPUT1), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n355_), .A2(new_n351_), .A3(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n335_), .B1(new_n354_), .B2(new_n358_), .ZN(new_n359_));
  AOI22_X1  g158(.A1(new_n347_), .A2(new_n349_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n360_));
  OAI211_X1 g159(.A(KEYINPUT90), .B(new_n357_), .C1(new_n360_), .C2(new_n337_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n334_), .B1(new_n359_), .B2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(G211gat), .ZN(new_n363_));
  INV_X1    g162(.A(G218gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G211gat), .A2(G218gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT94), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n365_), .A2(KEYINPUT94), .A3(new_n366_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G197gat), .B(G204gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(KEYINPUT93), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT21), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT21), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n372_), .A2(KEYINPUT93), .A3(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n371_), .A2(new_n374_), .A3(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT95), .ZN(new_n378_));
  OR2_X1    g177(.A1(new_n372_), .A2(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n375_), .B1(new_n372_), .B2(new_n378_), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n379_), .A2(new_n380_), .A3(new_n369_), .A4(new_n370_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n377_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n333_), .B1(new_n362_), .B2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n359_), .A2(new_n334_), .A3(new_n361_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n346_), .ZN(new_n386_));
  NOR3_X1   g185(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n345_), .ZN(new_n389_));
  AOI21_X1  g188(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n348_), .B1(new_n388_), .B2(new_n391_), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n351_), .A2(new_n352_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n336_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(new_n357_), .ZN(new_n395_));
  XOR2_X1   g194(.A(KEYINPUT96), .B(KEYINPUT29), .Z(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n333_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n397_), .A2(new_n382_), .A3(new_n398_), .ZN(new_n399_));
  AND3_X1   g198(.A1(new_n384_), .A2(new_n385_), .A3(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n385_), .B1(new_n384_), .B2(new_n399_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n331_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n385_), .ZN(new_n403_));
  AOI21_X1  g202(.A(KEYINPUT90), .B1(new_n394_), .B2(new_n357_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n361_), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT29), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n398_), .B1(new_n406_), .B2(new_n382_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n399_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n403_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n384_), .A2(new_n385_), .A3(new_n399_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n331_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n409_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n402_), .A2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G22gat), .B(G50gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT28), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n413_), .A2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n402_), .A2(new_n412_), .A3(new_n415_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  XOR2_X1   g218(.A(G71gat), .B(G99gat), .Z(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(KEYINPUT30), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G227gat), .A2(G233gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G169gat), .A2(G176gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(KEYINPUT22), .B(G169gat), .ZN(new_n425_));
  INV_X1    g224(.A(G176gat), .ZN(new_n426_));
  AOI21_X1  g225(.A(KEYINPUT85), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  AND2_X1   g226(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n428_));
  NOR2_X1   g227(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n429_));
  OAI211_X1 g228(.A(KEYINPUT85), .B(new_n426_), .C1(new_n428_), .C2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n424_), .B1(new_n427_), .B2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT87), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G183gat), .A2(G190gat), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT84), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(KEYINPUT84), .A2(G183gat), .A3(G190gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(KEYINPUT86), .B1(new_n434_), .B2(KEYINPUT23), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT86), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT23), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n440_), .A2(new_n441_), .A3(G183gat), .A4(G190gat), .ZN(new_n442_));
  AOI22_X1  g241(.A1(new_n438_), .A2(KEYINPUT23), .B1(new_n439_), .B2(new_n442_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(G183gat), .A2(G190gat), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n433_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n439_), .A2(new_n442_), .ZN(new_n446_));
  AND3_X1   g245(.A1(KEYINPUT84), .A2(G183gat), .A3(G190gat), .ZN(new_n447_));
  AOI21_X1  g246(.A(KEYINPUT84), .B1(G183gat), .B2(G190gat), .ZN(new_n448_));
  OAI21_X1  g247(.A(KEYINPUT23), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n446_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n444_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n450_), .A2(KEYINPUT87), .A3(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n432_), .B1(new_n445_), .B2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n434_), .A2(KEYINPUT23), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n454_), .B1(new_n438_), .B2(KEYINPUT23), .ZN(new_n455_));
  XNOR2_X1  g254(.A(KEYINPUT25), .B(G183gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(KEYINPUT26), .B(G190gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(KEYINPUT83), .B1(G169gat), .B2(G176gat), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NOR3_X1   g259(.A1(KEYINPUT83), .A2(G169gat), .A3(G176gat), .ZN(new_n461_));
  OAI211_X1 g260(.A(KEYINPUT24), .B(new_n424_), .C1(new_n460_), .C2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT83), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n463_), .A2(new_n315_), .A3(new_n426_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT24), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n464_), .A2(new_n465_), .A3(new_n459_), .ZN(new_n466_));
  AND4_X1   g265(.A1(new_n455_), .A2(new_n458_), .A3(new_n462_), .A4(new_n466_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n453_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(G120gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G127gat), .B(G134gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(G113gat), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n470_), .A2(G113gat), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n469_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  OR2_X1    g273(.A1(new_n470_), .A2(G113gat), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n475_), .A2(G120gat), .A3(new_n471_), .ZN(new_n476_));
  AND2_X1   g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n468_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n474_), .A2(new_n476_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n479_), .B1(new_n453_), .B2(new_n467_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G15gat), .B(G43gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT31), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n478_), .A2(new_n480_), .A3(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n483_), .B1(new_n478_), .B2(new_n480_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n423_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NOR3_X1   g287(.A1(new_n485_), .A2(new_n486_), .A3(new_n423_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n419_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT101), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G1gat), .B(G29gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(G85gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT0), .ZN(new_n495_));
  INV_X1    g294(.A(G57gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G225gat), .A2(G233gat), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT4), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n479_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n477_), .A2(new_n394_), .A3(new_n357_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n500_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n477_), .B1(new_n359_), .B2(new_n361_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n504_), .A2(KEYINPUT4), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n499_), .B1(new_n503_), .B2(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n501_), .A2(new_n498_), .A3(new_n502_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n497_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n395_), .A2(new_n479_), .ZN(new_n509_));
  OAI21_X1  g308(.A(KEYINPUT4), .B1(new_n504_), .B2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n501_), .A2(new_n500_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n498_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n507_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n497_), .ZN(new_n514_));
  NOR3_X1   g313(.A1(new_n512_), .A2(new_n513_), .A3(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n492_), .B1(new_n508_), .B2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n506_), .A2(new_n507_), .A3(new_n497_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n514_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n517_), .A2(new_n518_), .A3(KEYINPUT101), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G8gat), .B(G36gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT18), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(G64gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(new_n216_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G226gat), .A2(G233gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT19), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT20), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n528_), .B1(new_n468_), .B2(new_n383_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n465_), .A2(new_n315_), .A3(new_n426_), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n450_), .A2(new_n530_), .A3(new_n458_), .A4(new_n462_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT97), .ZN(new_n532_));
  AOI22_X1  g331(.A1(new_n464_), .A2(new_n459_), .B1(G169gat), .B2(G176gat), .ZN(new_n533_));
  AOI22_X1  g332(.A1(new_n533_), .A2(KEYINPUT24), .B1(new_n456_), .B2(new_n457_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT97), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n534_), .A2(new_n535_), .A3(new_n530_), .A4(new_n450_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n532_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n455_), .A2(new_n451_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n425_), .A2(new_n426_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n538_), .A2(new_n539_), .A3(new_n424_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n537_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(new_n382_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n527_), .B1(new_n529_), .B2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n537_), .A2(new_n383_), .A3(new_n540_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n382_), .B1(new_n453_), .B2(new_n467_), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n544_), .A2(new_n545_), .A3(KEYINPUT20), .A4(new_n527_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n524_), .B1(new_n543_), .B2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n445_), .A2(new_n452_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n432_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n467_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n551_), .A2(new_n383_), .A3(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT20), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n383_), .B1(new_n537_), .B2(new_n540_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n526_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n556_), .A2(new_n523_), .A3(new_n546_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n548_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT27), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT100), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n540_), .A2(new_n381_), .A3(new_n377_), .A4(new_n531_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n561_), .B1(new_n562_), .B2(KEYINPUT20), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n383_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n562_), .A2(new_n561_), .A3(KEYINPUT20), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n527_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  NOR3_X1   g366(.A1(new_n554_), .A2(new_n526_), .A3(new_n555_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n524_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n569_), .A2(KEYINPUT27), .A3(new_n557_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n516_), .A2(new_n519_), .A3(new_n560_), .A4(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(KEYINPUT103), .B1(new_n491_), .B2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n490_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n573_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n574_));
  AND2_X1   g373(.A1(new_n516_), .A2(new_n519_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT103), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n560_), .A2(new_n570_), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n574_), .A2(new_n575_), .A3(new_n576_), .A4(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n572_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT88), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n580_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n489_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n582_), .A2(KEYINPUT88), .A3(new_n487_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  AND3_X1   g383(.A1(new_n402_), .A2(new_n412_), .A3(new_n415_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n415_), .B1(new_n402_), .B2(new_n412_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n584_), .B1(new_n571_), .B2(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n499_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n589_));
  NOR3_X1   g388(.A1(new_n504_), .A2(new_n498_), .A3(new_n509_), .ZN(new_n590_));
  NOR3_X1   g389(.A1(new_n589_), .A2(new_n590_), .A3(new_n497_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n558_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT98), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n593_), .B1(new_n515_), .B2(KEYINPUT33), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT33), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n517_), .A2(KEYINPUT98), .A3(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n515_), .A2(KEYINPUT33), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n592_), .A2(new_n594_), .A3(new_n596_), .A4(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n517_), .A2(new_n518_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n567_), .A2(new_n568_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n523_), .A2(KEYINPUT32), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT99), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n556_), .A2(new_n602_), .A3(new_n546_), .ZN(new_n603_));
  AND3_X1   g402(.A1(new_n600_), .A2(new_n601_), .A3(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n543_), .A2(new_n547_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n601_), .B1(new_n605_), .B2(KEYINPUT99), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n599_), .B1(new_n604_), .B2(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n598_), .A2(new_n607_), .A3(new_n419_), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n588_), .A2(KEYINPUT102), .A3(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(KEYINPUT102), .B1(new_n588_), .B2(new_n608_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n579_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(G231gat), .ZN(new_n612_));
  INV_X1    g411(.A(G233gat), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n210_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n251_), .A2(new_n614_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n321_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n617_), .A2(new_n616_), .A3(new_n321_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n619_), .A2(new_n242_), .A3(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n620_), .ZN(new_n622_));
  OAI21_X1  g421(.A(KEYINPUT68), .B1(new_n622_), .B2(new_n618_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G127gat), .B(G155gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT16), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(G183gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(new_n363_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n628_), .A2(KEYINPUT17), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n621_), .A2(new_n623_), .A3(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT79), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT79), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n621_), .A2(new_n623_), .A3(new_n632_), .A4(new_n629_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n633_), .ZN(new_n634_));
  NOR3_X1   g433(.A1(new_n622_), .A2(new_n629_), .A3(new_n618_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n635_), .B1(KEYINPUT17), .B2(new_n628_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n634_), .A2(new_n636_), .ZN(new_n637_));
  AND3_X1   g436(.A1(new_n329_), .A2(new_n611_), .A3(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT37), .ZN(new_n639_));
  XNOR2_X1  g438(.A(G190gat), .B(G218gat), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(G134gat), .ZN(new_n641_));
  INV_X1    g440(.A(G162gat), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n641_), .B(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT36), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n643_), .A2(new_n644_), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n238_), .A2(new_n282_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(G232gat), .A2(G233gat), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n649_), .B(KEYINPUT72), .Z(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT34), .ZN(new_n651_));
  XOR2_X1   g450(.A(KEYINPUT73), .B(KEYINPUT35), .Z(new_n652_));
  AND2_X1   g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  OR2_X1    g452(.A1(new_n653_), .A2(KEYINPUT75), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(KEYINPUT75), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n648_), .A2(new_n654_), .A3(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(KEYINPUT76), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n322_), .A2(new_n238_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(KEYINPUT74), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT76), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n648_), .A2(new_n661_), .A3(new_n654_), .A4(new_n655_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT74), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n658_), .A2(new_n663_), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n657_), .A2(new_n660_), .A3(new_n662_), .A4(new_n664_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n651_), .A2(new_n652_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  OR3_X1    g466(.A1(new_n656_), .A2(new_n666_), .A3(new_n659_), .ZN(new_n668_));
  AOI211_X1 g467(.A(new_n646_), .B(new_n647_), .C1(new_n667_), .C2(new_n668_), .ZN(new_n669_));
  NAND4_X1  g468(.A1(new_n667_), .A2(new_n644_), .A3(new_n643_), .A4(new_n668_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n639_), .B1(new_n669_), .B2(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n647_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(new_n645_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n674_), .A2(KEYINPUT37), .A3(new_n670_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n672_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n638_), .A2(new_n677_), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n678_), .A2(G1gat), .A3(new_n575_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n679_), .A2(KEYINPUT38), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT105), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(KEYINPUT38), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT104), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n669_), .A2(new_n671_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n638_), .A2(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(G1gat), .B1(new_n686_), .B2(new_n575_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n681_), .A2(new_n683_), .A3(new_n687_), .ZN(G1324gat));
  INV_X1    g487(.A(KEYINPUT39), .ZN(new_n689_));
  INV_X1    g488(.A(new_n577_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n638_), .A2(new_n690_), .A3(new_n685_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n689_), .B1(new_n691_), .B2(G8gat), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n691_), .A2(new_n689_), .A3(G8gat), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n690_), .A2(new_n292_), .ZN(new_n695_));
  OAI22_X1  g494(.A1(new_n692_), .A2(new_n694_), .B1(new_n678_), .B2(new_n695_), .ZN(new_n696_));
  XOR2_X1   g495(.A(new_n696_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g496(.A(new_n584_), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n678_), .A2(G15gat), .A3(new_n698_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT106), .Z(new_n700_));
  OAI21_X1  g499(.A(G15gat), .B1(new_n686_), .B2(new_n698_), .ZN(new_n701_));
  XOR2_X1   g500(.A(new_n701_), .B(KEYINPUT41), .Z(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n702_), .ZN(G1326gat));
  OAI21_X1  g502(.A(G22gat), .B1(new_n686_), .B2(new_n419_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT42), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n419_), .A2(G22gat), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n705_), .B1(new_n678_), .B2(new_n706_), .ZN(G1327gat));
  NOR2_X1   g506(.A1(new_n685_), .A2(new_n637_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n329_), .A2(new_n611_), .A3(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n575_), .ZN(new_n711_));
  AOI21_X1  g510(.A(G29gat), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT43), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n611_), .A2(new_n713_), .A3(new_n676_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT107), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n611_), .A2(new_n676_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(KEYINPUT43), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n611_), .A2(KEYINPUT107), .A3(new_n713_), .A4(new_n676_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n716_), .A2(new_n718_), .A3(new_n719_), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n273_), .A2(new_n328_), .A3(new_n637_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT44), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n724_), .A2(G29gat), .A3(new_n711_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n720_), .A2(KEYINPUT44), .A3(new_n721_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n712_), .B1(new_n725_), .B2(new_n726_), .ZN(G1328gat));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n690_), .ZN(new_n728_));
  AOI21_X1  g527(.A(KEYINPUT44), .B1(new_n720_), .B2(new_n721_), .ZN(new_n729_));
  OAI21_X1  g528(.A(G36gat), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(G36gat), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n329_), .A2(new_n731_), .A3(new_n611_), .A4(new_n708_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n732_), .A2(new_n577_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT45), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n733_), .B(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(KEYINPUT108), .B1(new_n730_), .B2(new_n735_), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n736_), .A2(KEYINPUT109), .A3(KEYINPUT46), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n736_), .A2(KEYINPUT109), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT46), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n730_), .A2(new_n735_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n740_), .B2(KEYINPUT109), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n737_), .B1(new_n738_), .B2(new_n741_), .ZN(G1329gat));
  OAI21_X1  g541(.A(new_n276_), .B1(new_n709_), .B2(new_n698_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT111), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n724_), .A2(G43gat), .A3(new_n490_), .A4(new_n726_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT110), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n745_), .A2(new_n746_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n744_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT47), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT47), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n751_), .B(new_n744_), .C1(new_n747_), .C2(new_n748_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(G1330gat));
  AND3_X1   g552(.A1(new_n724_), .A2(new_n587_), .A3(new_n726_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n587_), .A2(new_n280_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT112), .ZN(new_n756_));
  OAI22_X1  g555(.A1(new_n754_), .A2(new_n280_), .B1(new_n709_), .B2(new_n756_), .ZN(G1331gat));
  AND2_X1   g556(.A1(new_n273_), .A2(new_n611_), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n758_), .A2(new_n328_), .A3(new_n637_), .A4(new_n685_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n759_), .A2(new_n496_), .A3(new_n575_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n634_), .A2(new_n328_), .A3(new_n636_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n676_), .A2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n758_), .A2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  OR2_X1    g563(.A1(new_n764_), .A2(KEYINPUT113), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(KEYINPUT113), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n765_), .A2(new_n711_), .A3(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n760_), .B1(new_n767_), .B2(new_n496_), .ZN(G1332gat));
  OAI21_X1  g567(.A(G64gat), .B1(new_n759_), .B2(new_n577_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT48), .ZN(new_n770_));
  OR2_X1    g569(.A1(new_n577_), .A2(G64gat), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n770_), .B1(new_n763_), .B2(new_n771_), .ZN(G1333gat));
  OAI21_X1  g571(.A(G71gat), .B1(new_n759_), .B2(new_n698_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT49), .ZN(new_n774_));
  OR2_X1    g573(.A1(new_n698_), .A2(G71gat), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n774_), .B1(new_n763_), .B2(new_n775_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT114), .ZN(G1334gat));
  OAI21_X1  g576(.A(G78gat), .B1(new_n759_), .B2(new_n419_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT50), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n419_), .A2(G78gat), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT115), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n779_), .B1(new_n763_), .B2(new_n781_), .ZN(G1335gat));
  NOR2_X1   g581(.A1(new_n637_), .A2(new_n327_), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n758_), .A2(new_n684_), .A3(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(G85gat), .B1(new_n784_), .B2(new_n711_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n720_), .A2(new_n273_), .A3(new_n783_), .ZN(new_n786_));
  XOR2_X1   g585(.A(new_n786_), .B(KEYINPUT116), .Z(new_n787_));
  AND2_X1   g586(.A1(new_n787_), .A2(new_n711_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n785_), .B1(new_n788_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g588(.A(G92gat), .B1(new_n784_), .B2(new_n690_), .ZN(new_n790_));
  AND2_X1   g589(.A1(new_n787_), .A2(new_n690_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n791_), .B2(G92gat), .ZN(G1337gat));
  OAI21_X1  g591(.A(G99gat), .B1(new_n786_), .B2(new_n698_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n224_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n784_), .A2(new_n794_), .A3(new_n490_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n793_), .A2(new_n795_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g596(.A(G106gat), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n784_), .A2(new_n798_), .A3(new_n587_), .ZN(new_n799_));
  OR2_X1    g598(.A1(new_n786_), .A2(new_n419_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT52), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n800_), .A2(new_n801_), .A3(G106gat), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n801_), .B1(new_n800_), .B2(G106gat), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n799_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(KEYINPUT53), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n806_), .B(new_n799_), .C1(new_n802_), .C2(new_n803_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n805_), .A2(new_n807_), .ZN(G1339gat));
  NAND2_X1  g607(.A1(new_n762_), .A2(new_n272_), .ZN(new_n809_));
  AOI21_X1  g608(.A(KEYINPUT117), .B1(new_n809_), .B2(KEYINPUT54), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT117), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n812_));
  AOI211_X1 g611(.A(new_n811_), .B(new_n812_), .C1(new_n762_), .C2(new_n272_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n809_), .A2(KEYINPUT54), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n810_), .A2(new_n813_), .A3(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n637_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n312_), .B1(new_n307_), .B2(new_n310_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n323_), .A2(new_n311_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n318_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n318_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n313_), .A2(new_n820_), .A3(new_n324_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n819_), .A2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n822_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(KEYINPUT55), .B1(new_n255_), .B2(new_n257_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n252_), .A2(new_n253_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n240_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n828_), .B1(new_n829_), .B2(new_n254_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n263_), .B1(new_n825_), .B2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT56), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT118), .ZN(new_n834_));
  OAI211_X1 g633(.A(KEYINPUT56), .B(new_n263_), .C1(new_n825_), .C2(new_n830_), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n833_), .A2(new_n834_), .A3(new_n835_), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n327_), .B(new_n266_), .C1(new_n835_), .C2(new_n834_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n824_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n838_), .A2(KEYINPUT57), .A3(new_n685_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT120), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n838_), .A2(KEYINPUT120), .A3(KEYINPUT57), .A4(new_n685_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n327_), .A2(new_n266_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n835_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n845_), .B1(new_n846_), .B2(KEYINPUT118), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n833_), .A2(new_n834_), .A3(new_n835_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n823_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n844_), .B1(new_n849_), .B2(new_n684_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(KEYINPUT119), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT119), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n852_), .B(new_n844_), .C1(new_n849_), .C2(new_n684_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n833_), .A2(new_n835_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n822_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n855_), .A2(new_n266_), .A3(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT58), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n855_), .A2(KEYINPUT58), .A3(new_n266_), .A4(new_n856_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n859_), .A2(new_n676_), .A3(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n843_), .A2(new_n854_), .A3(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n815_), .B1(new_n816_), .B2(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n711_), .A2(new_n574_), .A3(new_n577_), .ZN(new_n864_));
  OAI21_X1  g663(.A(KEYINPUT121), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n862_), .A2(new_n816_), .ZN(new_n866_));
  OR3_X1    g665(.A1(new_n810_), .A2(new_n813_), .A3(new_n814_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n864_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT121), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n865_), .A2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n327_), .ZN(new_n872_));
  INV_X1    g671(.A(G113gat), .ZN(new_n873_));
  OAI21_X1  g672(.A(KEYINPUT59), .B1(new_n863_), .B2(new_n864_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n864_), .A2(KEYINPUT59), .ZN(new_n875_));
  INV_X1    g674(.A(new_n861_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n876_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n637_), .B1(new_n877_), .B2(new_n850_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n875_), .B1(new_n878_), .B2(new_n815_), .ZN(new_n879_));
  AND2_X1   g678(.A1(new_n874_), .A2(new_n879_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(KEYINPUT122), .B(G113gat), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n327_), .A2(new_n881_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(KEYINPUT123), .ZN(new_n883_));
  AOI22_X1  g682(.A1(new_n872_), .A2(new_n873_), .B1(new_n880_), .B2(new_n883_), .ZN(G1340gat));
  INV_X1    g683(.A(KEYINPUT59), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n273_), .B(new_n879_), .C1(new_n868_), .C2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(KEYINPUT124), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT124), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n874_), .A2(new_n888_), .A3(new_n273_), .A4(new_n879_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n887_), .A2(new_n889_), .A3(G120gat), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n469_), .B1(new_n272_), .B2(KEYINPUT60), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n871_), .B(new_n891_), .C1(KEYINPUT60), .C2(new_n469_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n890_), .A2(new_n892_), .ZN(G1341gat));
  AOI21_X1  g692(.A(G127gat), .B1(new_n871_), .B2(new_n637_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT125), .ZN(new_n895_));
  OR2_X1    g694(.A1(new_n895_), .A2(G127gat), .ZN(new_n896_));
  OAI21_X1  g695(.A(G127gat), .B1(new_n816_), .B2(new_n895_), .ZN(new_n897_));
  AND4_X1   g696(.A1(new_n874_), .A2(new_n879_), .A3(new_n896_), .A4(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n894_), .A2(new_n898_), .ZN(G1342gat));
  NAND2_X1  g698(.A1(new_n871_), .A2(new_n684_), .ZN(new_n900_));
  INV_X1    g699(.A(G134gat), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n677_), .A2(new_n901_), .ZN(new_n902_));
  AOI22_X1  g701(.A1(new_n900_), .A2(new_n901_), .B1(new_n880_), .B2(new_n902_), .ZN(G1343gat));
  NAND2_X1  g702(.A1(new_n866_), .A2(new_n867_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n904_), .A2(new_n587_), .A3(new_n698_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n711_), .A2(new_n577_), .ZN(new_n906_));
  NOR3_X1   g705(.A1(new_n905_), .A2(new_n328_), .A3(new_n906_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(new_n339_), .ZN(G1344gat));
  NOR3_X1   g707(.A1(new_n905_), .A2(new_n272_), .A3(new_n906_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(new_n340_), .ZN(G1345gat));
  NOR3_X1   g709(.A1(new_n905_), .A2(new_n816_), .A3(new_n906_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(KEYINPUT61), .B(G155gat), .ZN(new_n912_));
  INV_X1    g711(.A(new_n912_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n911_), .B(new_n913_), .ZN(G1346gat));
  NOR2_X1   g713(.A1(new_n905_), .A2(new_n906_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(new_n684_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n677_), .A2(new_n642_), .ZN(new_n917_));
  AOI22_X1  g716(.A1(new_n916_), .A2(new_n642_), .B1(new_n915_), .B2(new_n917_), .ZN(G1347gat));
  OR2_X1    g717(.A1(new_n878_), .A2(new_n815_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n711_), .A2(new_n577_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n920_), .A2(new_n419_), .A3(new_n584_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n921_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n919_), .A2(new_n327_), .A3(new_n922_), .ZN(new_n923_));
  XOR2_X1   g722(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n924_));
  INV_X1    g723(.A(new_n924_), .ZN(new_n925_));
  AND3_X1   g724(.A1(new_n923_), .A2(G169gat), .A3(new_n925_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n925_), .B1(new_n923_), .B2(G169gat), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n919_), .A2(new_n922_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n327_), .A2(new_n425_), .ZN(new_n929_));
  XOR2_X1   g728(.A(new_n929_), .B(KEYINPUT127), .Z(new_n930_));
  OAI22_X1  g729(.A1(new_n926_), .A2(new_n927_), .B1(new_n928_), .B2(new_n930_), .ZN(G1348gat));
  INV_X1    g730(.A(new_n928_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n932_), .A2(new_n426_), .A3(new_n273_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n273_), .A2(new_n922_), .ZN(new_n934_));
  OAI21_X1  g733(.A(G176gat), .B1(new_n863_), .B2(new_n934_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n933_), .A2(new_n935_), .ZN(G1349gat));
  NOR3_X1   g735(.A1(new_n928_), .A2(new_n456_), .A3(new_n816_), .ZN(new_n937_));
  INV_X1    g736(.A(G183gat), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n815_), .A2(new_n637_), .A3(new_n922_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n937_), .B1(new_n938_), .B2(new_n939_), .ZN(G1350gat));
  OAI21_X1  g739(.A(G190gat), .B1(new_n928_), .B2(new_n677_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n684_), .A2(new_n457_), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n941_), .B1(new_n928_), .B2(new_n942_), .ZN(G1351gat));
  INV_X1    g742(.A(new_n920_), .ZN(new_n944_));
  NOR3_X1   g743(.A1(new_n905_), .A2(new_n328_), .A3(new_n944_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(new_n945_), .B(new_n317_), .ZN(G1352gat));
  NOR3_X1   g745(.A1(new_n905_), .A2(new_n272_), .A3(new_n944_), .ZN(new_n947_));
  INV_X1    g746(.A(G204gat), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n947_), .B(new_n948_), .ZN(G1353gat));
  XNOR2_X1  g748(.A(KEYINPUT63), .B(G211gat), .ZN(new_n950_));
  NOR4_X1   g749(.A1(new_n905_), .A2(new_n816_), .A3(new_n944_), .A4(new_n950_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n905_), .A2(new_n944_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n952_), .A2(new_n637_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n951_), .B1(new_n953_), .B2(new_n954_), .ZN(G1354gat));
  NAND2_X1  g754(.A1(new_n952_), .A2(new_n684_), .ZN(new_n956_));
  NOR2_X1   g755(.A1(new_n677_), .A2(new_n364_), .ZN(new_n957_));
  AOI22_X1  g756(.A1(new_n956_), .A2(new_n364_), .B1(new_n952_), .B2(new_n957_), .ZN(G1355gat));
endmodule


