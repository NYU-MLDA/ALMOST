//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 0 1 1 0 1 0 0 1 0 1 0 1 1 0 0 1 1 1 0 0 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 1 0 1 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n671_,
    new_n672_, new_n673_, new_n675_, new_n676_, new_n677_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n779_, new_n780_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n886_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_, new_n923_,
    new_n924_, new_n925_, new_n927_, new_n928_, new_n929_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n936_, new_n937_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_;
  INV_X1    g000(.A(KEYINPUT38), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G1gat), .B(G8gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT78), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT79), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT14), .ZN(new_n208_));
  INV_X1    g007(.A(G1gat), .ZN(new_n209_));
  INV_X1    g008(.A(G8gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(G15gat), .ZN(new_n212_));
  INV_X1    g011(.A(G22gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G15gat), .A2(G22gat), .ZN(new_n215_));
  OAI22_X1  g014(.A1(new_n208_), .A2(new_n211_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n207_), .A2(new_n216_), .ZN(new_n217_));
  OR2_X1    g016(.A1(new_n205_), .A2(new_n206_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n216_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n205_), .A2(new_n206_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n217_), .A2(new_n221_), .ZN(new_n222_));
  XOR2_X1   g021(.A(G29gat), .B(G36gat), .Z(new_n223_));
  XOR2_X1   g022(.A(G43gat), .B(G50gat), .Z(new_n224_));
  XOR2_X1   g023(.A(new_n223_), .B(new_n224_), .Z(new_n225_));
  NAND2_X1  g024(.A1(new_n222_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n225_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n217_), .A2(new_n221_), .A3(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(KEYINPUT82), .A3(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G229gat), .A2(G233gat), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT82), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n222_), .A2(new_n232_), .A3(new_n225_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n229_), .A2(new_n231_), .A3(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT75), .B(KEYINPUT15), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n225_), .B(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n222_), .A2(new_n236_), .ZN(new_n237_));
  NAND4_X1  g036(.A1(new_n237_), .A2(KEYINPUT83), .A3(new_n228_), .A4(new_n230_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n237_), .A2(new_n230_), .A3(new_n228_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT83), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n234_), .A2(new_n238_), .A3(new_n241_), .ZN(new_n242_));
  XOR2_X1   g041(.A(G113gat), .B(G141gat), .Z(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT84), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G169gat), .B(G197gat), .ZN(new_n245_));
  XOR2_X1   g044(.A(new_n244_), .B(new_n245_), .Z(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n242_), .A2(new_n247_), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n234_), .A2(new_n241_), .A3(new_n238_), .A4(new_n246_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT24), .ZN(new_n252_));
  NOR2_X1   g051(.A1(G169gat), .A2(G176gat), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT86), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n253_), .B(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT25), .B(G183gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT26), .B(G190gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT85), .ZN(new_n259_));
  AOI22_X1  g058(.A1(new_n252_), .A2(new_n255_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT23), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n261_), .B1(G183gat), .B2(G190gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G183gat), .A2(G190gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT87), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n262_), .B1(new_n264_), .B2(new_n261_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n256_), .A2(new_n257_), .A3(KEYINPUT85), .ZN(new_n267_));
  INV_X1    g066(.A(new_n255_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n252_), .B1(G169gat), .B2(G176gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n260_), .A2(new_n266_), .A3(new_n267_), .A4(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n272_), .B1(new_n264_), .B2(KEYINPUT23), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n273_), .B1(G183gat), .B2(G190gat), .ZN(new_n274_));
  NOR2_X1   g073(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(G169gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n274_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n271_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT30), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n271_), .A2(new_n277_), .A3(KEYINPUT30), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  OR2_X1    g081(.A1(new_n282_), .A2(KEYINPUT89), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(KEYINPUT89), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G227gat), .A2(G233gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(G15gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT88), .B(G43gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  XOR2_X1   g088(.A(G71gat), .B(G99gat), .Z(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n285_), .A2(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n282_), .A2(KEYINPUT89), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n294_), .A2(new_n292_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  XOR2_X1   g095(.A(G127gat), .B(G134gat), .Z(new_n297_));
  XOR2_X1   g096(.A(G113gat), .B(G120gat), .Z(new_n298_));
  XOR2_X1   g097(.A(new_n297_), .B(new_n298_), .Z(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT31), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n293_), .A2(new_n296_), .A3(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n300_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n291_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n302_), .B1(new_n303_), .B2(new_n295_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n301_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT20), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G169gat), .A2(G176gat), .ZN(new_n308_));
  NOR2_X1   g107(.A1(G183gat), .A2(G190gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT22), .B(G169gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT100), .ZN(new_n311_));
  OAI221_X1 g110(.A(new_n308_), .B1(new_n265_), .B2(new_n309_), .C1(G176gat), .C2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n269_), .A2(KEYINPUT99), .ZN(new_n313_));
  OR2_X1    g112(.A1(new_n269_), .A2(KEYINPUT99), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n268_), .A2(new_n313_), .A3(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n253_), .A2(new_n252_), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n315_), .A2(new_n273_), .A3(new_n258_), .A4(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n312_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT21), .ZN(new_n319_));
  XOR2_X1   g118(.A(KEYINPUT92), .B(G197gat), .Z(new_n320_));
  INV_X1    g119(.A(KEYINPUT93), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n320_), .A2(new_n321_), .A3(G204gat), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(G197gat), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT93), .B1(new_n324_), .B2(G204gat), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n325_), .B1(new_n320_), .B2(G204gat), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n319_), .B1(new_n323_), .B2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G211gat), .B(G218gat), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(G204gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n320_), .A2(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n319_), .B1(G197gat), .B2(G204gat), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n329_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n327_), .A2(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n323_), .A2(new_n326_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n329_), .A2(KEYINPUT94), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT94), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n319_), .B1(new_n328_), .B2(new_n337_), .ZN(new_n338_));
  AND2_X1   g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n335_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n334_), .A2(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n307_), .B1(new_n318_), .B2(new_n341_), .ZN(new_n342_));
  AOI22_X1  g141(.A1(new_n327_), .A2(new_n333_), .B1(new_n335_), .B2(new_n339_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n343_), .A2(new_n271_), .A3(new_n277_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n342_), .A2(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT98), .B(KEYINPUT19), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G226gat), .A2(G233gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n345_), .A2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n343_), .A2(new_n317_), .A3(new_n312_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n341_), .A2(new_n278_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n348_), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n350_), .A2(new_n351_), .A3(KEYINPUT20), .A4(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n349_), .A2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G8gat), .B(G36gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT18), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G64gat), .B(G92gat), .ZN(new_n357_));
  XOR2_X1   g156(.A(new_n356_), .B(new_n357_), .Z(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n354_), .A2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n349_), .A2(new_n358_), .A3(new_n353_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT27), .ZN(new_n362_));
  AND3_X1   g161(.A1(new_n360_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT102), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n350_), .A2(new_n351_), .A3(KEYINPUT20), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(new_n348_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n342_), .A2(new_n352_), .A3(new_n344_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n364_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(KEYINPUT102), .B1(new_n365_), .B2(new_n348_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n359_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT105), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n361_), .A2(new_n371_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n349_), .A2(KEYINPUT105), .A3(new_n358_), .A4(new_n353_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n370_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n363_), .B1(new_n374_), .B2(KEYINPUT27), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G155gat), .B(G162gat), .ZN(new_n376_));
  NAND3_X1  g175(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT90), .ZN(new_n378_));
  INV_X1    g177(.A(G141gat), .ZN(new_n379_));
  INV_X1    g178(.A(G148gat), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n379_), .A2(new_n380_), .A3(KEYINPUT3), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT3), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n382_), .B1(G141gat), .B2(G148gat), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT2), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G141gat), .A2(G148gat), .ZN(new_n385_));
  AOI22_X1  g184(.A1(new_n381_), .A2(new_n383_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n376_), .B1(new_n378_), .B2(new_n386_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n376_), .A2(KEYINPUT1), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n379_), .A2(new_n380_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n389_), .A2(new_n390_), .A3(new_n385_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n388_), .A2(new_n391_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n387_), .A2(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(new_n299_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(KEYINPUT4), .ZN(new_n395_));
  INV_X1    g194(.A(new_n393_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(new_n299_), .ZN(new_n397_));
  OR2_X1    g196(.A1(new_n397_), .A2(KEYINPUT4), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G225gat), .A2(G233gat), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n395_), .A2(new_n398_), .A3(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G1gat), .B(G29gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(G85gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT0), .B(G57gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n299_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(new_n393_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n397_), .A2(new_n408_), .A3(new_n399_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT101), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT101), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n394_), .A2(new_n411_), .A3(new_n399_), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n401_), .A2(new_n406_), .A3(new_n410_), .A4(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(KEYINPUT103), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n401_), .A2(new_n410_), .A3(new_n412_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(new_n405_), .ZN(new_n416_));
  AND2_X1   g215(.A1(new_n410_), .A2(new_n412_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT103), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n417_), .A2(new_n418_), .A3(new_n406_), .A4(new_n401_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n414_), .A2(new_n416_), .A3(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT104), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n396_), .A2(KEYINPUT29), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G228gat), .A2(G233gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(KEYINPUT95), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n424_), .A2(KEYINPUT95), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  AOI22_X1  g226(.A1(new_n341_), .A2(new_n423_), .B1(new_n425_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G78gat), .B(G106gat), .ZN(new_n430_));
  XOR2_X1   g229(.A(new_n430_), .B(KEYINPUT96), .Z(new_n431_));
  NAND3_X1  g230(.A1(new_n341_), .A2(new_n423_), .A3(new_n427_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n429_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n431_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n432_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n434_), .B1(new_n435_), .B2(new_n428_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT29), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n393_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT28), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n438_), .B(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G22gat), .B(G50gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n438_), .B(KEYINPUT28), .ZN(new_n443_));
  INV_X1    g242(.A(new_n441_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n433_), .A2(new_n436_), .A3(new_n442_), .A4(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT97), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n429_), .A2(new_n447_), .A3(new_n431_), .A4(new_n432_), .ZN(new_n448_));
  AND3_X1   g247(.A1(new_n442_), .A2(new_n445_), .A3(KEYINPUT91), .ZN(new_n449_));
  AOI21_X1  g248(.A(KEYINPUT91), .B1(new_n442_), .B2(new_n445_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n448_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  AND3_X1   g250(.A1(new_n433_), .A2(new_n436_), .A3(KEYINPUT97), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n446_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n414_), .A2(new_n416_), .A3(new_n419_), .A4(KEYINPUT104), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n422_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n375_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n358_), .A2(KEYINPUT32), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n458_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n349_), .A2(new_n457_), .A3(new_n353_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n420_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  AND3_X1   g260(.A1(new_n395_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n394_), .A2(new_n400_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n405_), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT33), .B1(new_n462_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(new_n413_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n417_), .A2(KEYINPUT33), .A3(new_n406_), .A4(new_n401_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n466_), .A2(new_n360_), .A3(new_n467_), .A4(new_n361_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n453_), .B1(new_n461_), .B2(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n306_), .B1(new_n456_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n374_), .A2(KEYINPUT27), .ZN(new_n471_));
  INV_X1    g270(.A(new_n363_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n422_), .A2(new_n454_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n453_), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n473_), .A2(new_n475_), .A3(new_n476_), .A4(new_n305_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n251_), .B1(new_n470_), .B2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(G64gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(G57gat), .ZN(new_n480_));
  INV_X1    g279(.A(G57gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(G64gat), .ZN(new_n482_));
  AND3_X1   g281(.A1(new_n480_), .A2(new_n482_), .A3(KEYINPUT69), .ZN(new_n483_));
  AOI21_X1  g282(.A(KEYINPUT69), .B1(new_n480_), .B2(new_n482_), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT11), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n480_), .A2(new_n482_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT69), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT11), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n480_), .A2(new_n482_), .A3(KEYINPUT69), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n488_), .A2(new_n489_), .A3(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G71gat), .B(G78gat), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n485_), .A2(new_n491_), .A3(new_n493_), .ZN(new_n494_));
  OAI211_X1 g293(.A(KEYINPUT11), .B(new_n492_), .C1(new_n483_), .C2(new_n484_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  XOR2_X1   g296(.A(KEYINPUT10), .B(G99gat), .Z(new_n498_));
  AND2_X1   g297(.A1(KEYINPUT64), .A2(G106gat), .ZN(new_n499_));
  NOR2_X1   g298(.A1(KEYINPUT64), .A2(G106gat), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  AND2_X1   g300(.A1(G85gat), .A2(G92gat), .ZN(new_n502_));
  NOR2_X1   g301(.A1(G85gat), .A2(G92gat), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  AOI22_X1  g303(.A1(new_n498_), .A2(new_n501_), .B1(new_n504_), .B2(KEYINPUT9), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G99gat), .A2(G106gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(KEYINPUT6), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT6), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n508_), .A2(G99gat), .A3(G106gat), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT9), .ZN(new_n510_));
  AOI22_X1  g309(.A1(new_n507_), .A2(new_n509_), .B1(new_n502_), .B2(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(KEYINPUT65), .B1(new_n505_), .B2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(G85gat), .ZN(new_n513_));
  INV_X1    g312(.A(G92gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G85gat), .A2(G92gat), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n515_), .A2(KEYINPUT9), .A3(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(KEYINPUT10), .B(G99gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(KEYINPUT64), .B(G106gat), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n517_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n508_), .B1(G99gat), .B2(G106gat), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n506_), .A2(KEYINPUT6), .ZN(new_n522_));
  OAI22_X1  g321(.A1(new_n521_), .A2(new_n522_), .B1(KEYINPUT9), .B2(new_n516_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT65), .ZN(new_n524_));
  NOR3_X1   g323(.A1(new_n520_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  OAI22_X1  g324(.A1(KEYINPUT66), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n526_));
  NOR2_X1   g325(.A1(G99gat), .A2(G106gat), .ZN(new_n527_));
  NOR2_X1   g326(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  OAI211_X1 g328(.A(new_n526_), .B(new_n529_), .C1(new_n521_), .C2(new_n522_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT8), .ZN(new_n531_));
  NOR3_X1   g330(.A1(new_n502_), .A2(new_n503_), .A3(KEYINPUT67), .ZN(new_n532_));
  AND3_X1   g331(.A1(new_n530_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n531_), .B1(new_n530_), .B2(new_n532_), .ZN(new_n534_));
  OAI22_X1  g333(.A1(new_n512_), .A2(new_n525_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n497_), .A2(new_n535_), .A3(KEYINPUT12), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G230gat), .A2(G233gat), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n521_), .A2(new_n522_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n529_), .A2(new_n526_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n532_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(KEYINPUT8), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n530_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n524_), .B1(new_n520_), .B2(new_n523_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n498_), .A2(new_n501_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n546_), .A2(KEYINPUT65), .A3(new_n511_), .A4(new_n517_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n545_), .A2(new_n547_), .ZN(new_n548_));
  AND3_X1   g347(.A1(new_n544_), .A2(KEYINPUT68), .A3(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(KEYINPUT68), .B1(new_n544_), .B2(new_n548_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT70), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n494_), .A2(new_n552_), .A3(new_n495_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n552_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n538_), .B1(new_n551_), .B2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT68), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n535_), .A2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n544_), .A2(KEYINPUT68), .A3(new_n548_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n496_), .A2(KEYINPUT70), .ZN(new_n561_));
  AOI22_X1  g360(.A1(new_n559_), .A2(new_n560_), .B1(new_n561_), .B2(new_n553_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT72), .ZN(new_n563_));
  NOR3_X1   g362(.A1(new_n562_), .A2(new_n563_), .A3(KEYINPUT12), .ZN(new_n564_));
  OAI22_X1  g363(.A1(new_n549_), .A2(new_n550_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT12), .ZN(new_n566_));
  AOI21_X1  g365(.A(KEYINPUT72), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  OAI211_X1 g366(.A(new_n536_), .B(new_n557_), .C1(new_n564_), .C2(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(G120gat), .B(G148gat), .Z(new_n569_));
  XNOR2_X1  g368(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G176gat), .B(G204gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n565_), .B(KEYINPUT71), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n551_), .A2(new_n556_), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  OAI211_X1 g375(.A(new_n568_), .B(new_n573_), .C1(new_n576_), .C2(new_n537_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n573_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n568_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n537_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n578_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT74), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n577_), .A2(new_n581_), .A3(new_n582_), .ZN(new_n583_));
  OAI211_X1 g382(.A(KEYINPUT74), .B(new_n578_), .C1(new_n579_), .C2(new_n580_), .ZN(new_n584_));
  AOI21_X1  g383(.A(KEYINPUT13), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n583_), .A2(KEYINPUT13), .A3(new_n584_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G231gat), .A2(G233gat), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n589_), .B(KEYINPUT80), .Z(new_n590_));
  XNOR2_X1  g389(.A(new_n222_), .B(new_n590_), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n591_), .A2(new_n556_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n556_), .ZN(new_n593_));
  XOR2_X1   g392(.A(G127gat), .B(G155gat), .Z(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT16), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G183gat), .B(G211gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT17), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n592_), .A2(new_n593_), .A3(new_n598_), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n591_), .A2(KEYINPUT81), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n591_), .A2(KEYINPUT81), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n600_), .A2(new_n497_), .A3(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT17), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n597_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n497_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n599_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(KEYINPUT76), .A2(KEYINPUT37), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n608_), .B(KEYINPUT77), .Z(new_n609_));
  XNOR2_X1  g408(.A(G190gat), .B(G218gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G134gat), .B(G162gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n612_), .B(KEYINPUT36), .Z(new_n613_));
  NAND2_X1  g412(.A1(new_n551_), .A2(new_n227_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(G232gat), .A2(G233gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT34), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT35), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  AOI22_X1  g419(.A1(new_n236_), .A2(new_n535_), .B1(new_n618_), .B2(new_n617_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n614_), .A2(new_n620_), .A3(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n620_), .B1(new_n614_), .B2(new_n621_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n613_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n624_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n612_), .A2(KEYINPUT36), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n626_), .A2(new_n627_), .A3(new_n622_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n625_), .A2(new_n628_), .ZN(new_n629_));
  OR2_X1    g428(.A1(KEYINPUT76), .A2(KEYINPUT37), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n609_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n629_), .A2(new_n630_), .A3(new_n609_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n607_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n478_), .A2(new_n588_), .A3(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT106), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n635_), .B(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n474_), .A2(new_n209_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n202_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n635_), .B(KEYINPUT106), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n640_), .A2(KEYINPUT38), .A3(new_n209_), .A4(new_n474_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n588_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n642_), .A2(new_n251_), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n461_), .A2(new_n468_), .ZN(new_n644_));
  OAI22_X1  g443(.A1(new_n644_), .A2(new_n453_), .B1(new_n375_), .B2(new_n455_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n375_), .A2(new_n453_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n306_), .A2(new_n474_), .ZN(new_n647_));
  AOI22_X1  g446(.A1(new_n645_), .A2(new_n306_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n629_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n607_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n643_), .A2(new_n650_), .A3(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(G1gat), .B1(new_n652_), .B2(new_n475_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n639_), .A2(new_n641_), .A3(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT107), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n639_), .A2(new_n641_), .A3(KEYINPUT107), .A4(new_n653_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(G1324gat));
  NAND3_X1  g457(.A1(new_n640_), .A2(new_n210_), .A3(new_n375_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT39), .ZN(new_n660_));
  INV_X1    g459(.A(new_n652_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(new_n375_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n660_), .B1(new_n662_), .B2(G8gat), .ZN(new_n663_));
  AOI211_X1 g462(.A(KEYINPUT39), .B(new_n210_), .C1(new_n661_), .C2(new_n375_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n659_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(new_n668_));
  OAI211_X1 g467(.A(new_n659_), .B(new_n666_), .C1(new_n663_), .C2(new_n664_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(G1325gat));
  OAI21_X1  g469(.A(G15gat), .B1(new_n652_), .B2(new_n306_), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n671_), .B(KEYINPUT41), .Z(new_n672_));
  NAND3_X1  g471(.A1(new_n640_), .A2(new_n212_), .A3(new_n305_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1326gat));
  OAI21_X1  g473(.A(G22gat), .B1(new_n652_), .B2(new_n476_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT42), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n640_), .A2(new_n213_), .A3(new_n453_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(G1327gat));
  NOR2_X1   g477(.A1(new_n651_), .A2(new_n629_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n588_), .A2(new_n679_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n680_), .A2(new_n478_), .ZN(new_n681_));
  AOI21_X1  g480(.A(G29gat), .B1(new_n681_), .B2(new_n474_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n588_), .A2(new_n250_), .A3(new_n607_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT43), .ZN(new_n685_));
  INV_X1    g484(.A(new_n455_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n469_), .B1(new_n473_), .B2(new_n686_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n477_), .B1(new_n687_), .B2(new_n305_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT109), .ZN(new_n689_));
  INV_X1    g488(.A(new_n633_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n689_), .B1(new_n690_), .B2(new_n631_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n632_), .A2(KEYINPUT109), .A3(new_n633_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n685_), .B1(new_n688_), .B2(new_n693_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n690_), .A2(new_n631_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(new_n685_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n648_), .A2(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n684_), .B1(new_n694_), .B2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT110), .ZN(new_n701_));
  AOI21_X1  g500(.A(KEYINPUT44), .B1(new_n698_), .B2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n693_), .ZN(new_n703_));
  OAI21_X1  g502(.A(KEYINPUT43), .B1(new_n648_), .B2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n688_), .A2(new_n685_), .A3(new_n695_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n683_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(KEYINPUT110), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n700_), .B1(new_n702_), .B2(new_n707_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n474_), .A2(G29gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n682_), .B1(new_n708_), .B2(new_n709_), .ZN(G1328gat));
  INV_X1    g509(.A(KEYINPUT111), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT46), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n706_), .A2(KEYINPUT44), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n699_), .B1(new_n706_), .B2(KEYINPUT110), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n698_), .A2(new_n701_), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n375_), .B(new_n715_), .C1(new_n716_), .C2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(G36gat), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n473_), .A2(G36gat), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n478_), .A2(new_n588_), .A3(new_n679_), .A4(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(KEYINPUT45), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT45), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n680_), .A2(new_n723_), .A3(new_n478_), .A4(new_n720_), .ZN(new_n724_));
  AOI22_X1  g523(.A1(new_n722_), .A2(new_n724_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n714_), .B1(new_n719_), .B2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n725_), .ZN(new_n727_));
  AOI211_X1 g526(.A(new_n713_), .B(new_n727_), .C1(new_n718_), .C2(G36gat), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n726_), .A2(new_n728_), .ZN(G1329gat));
  INV_X1    g528(.A(KEYINPUT47), .ZN(new_n730_));
  INV_X1    g529(.A(G43gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n731_), .B1(new_n708_), .B2(new_n305_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n681_), .A2(new_n731_), .A3(new_n305_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n730_), .B1(new_n732_), .B2(new_n734_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n715_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n736_));
  OAI21_X1  g535(.A(G43gat), .B1(new_n736_), .B2(new_n306_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n737_), .A2(KEYINPUT47), .A3(new_n733_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n735_), .A2(new_n738_), .ZN(G1330gat));
  AOI21_X1  g538(.A(G50gat), .B1(new_n681_), .B2(new_n453_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n453_), .A2(G50gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n708_), .B2(new_n741_), .ZN(G1331gat));
  NOR3_X1   g541(.A1(new_n648_), .A2(new_n588_), .A3(new_n250_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n743_), .A2(new_n634_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n744_), .A2(new_n481_), .A3(new_n474_), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n650_), .A2(new_n251_), .A3(new_n642_), .A4(new_n651_), .ZN(new_n746_));
  OAI21_X1  g545(.A(G57gat), .B1(new_n746_), .B2(new_n475_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n747_), .ZN(G1332gat));
  OAI21_X1  g547(.A(G64gat), .B1(new_n746_), .B2(new_n473_), .ZN(new_n749_));
  XOR2_X1   g548(.A(KEYINPUT112), .B(KEYINPUT48), .Z(new_n750_));
  XNOR2_X1  g549(.A(new_n749_), .B(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n744_), .A2(new_n479_), .A3(new_n375_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(G1333gat));
  OAI21_X1  g552(.A(G71gat), .B1(new_n746_), .B2(new_n306_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(KEYINPUT113), .B(KEYINPUT49), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n754_), .B(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(G71gat), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n744_), .A2(new_n757_), .A3(new_n305_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(G1334gat));
  INV_X1    g558(.A(G78gat), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n744_), .A2(new_n760_), .A3(new_n453_), .ZN(new_n761_));
  OR2_X1    g560(.A1(new_n746_), .A2(new_n476_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT50), .ZN(new_n763_));
  AND3_X1   g562(.A1(new_n762_), .A2(new_n763_), .A3(G78gat), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n762_), .B2(G78gat), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n761_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT114), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT114), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n768_), .B(new_n761_), .C1(new_n764_), .C2(new_n765_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(G1335gat));
  NAND2_X1  g569(.A1(new_n704_), .A2(new_n705_), .ZN(new_n771_));
  NOR3_X1   g570(.A1(new_n588_), .A2(new_n250_), .A3(new_n651_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(G85gat), .B1(new_n773_), .B2(new_n475_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n743_), .A2(new_n679_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n776_), .A2(new_n513_), .A3(new_n474_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n774_), .A2(new_n777_), .ZN(G1336gat));
  OAI21_X1  g577(.A(G92gat), .B1(new_n773_), .B2(new_n473_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n776_), .A2(new_n514_), .A3(new_n375_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(G1337gat));
  NAND3_X1  g580(.A1(new_n776_), .A2(new_n305_), .A3(new_n498_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n771_), .A2(new_n305_), .A3(new_n772_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT115), .ZN(new_n784_));
  AND3_X1   g583(.A1(new_n783_), .A2(new_n784_), .A3(G99gat), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n784_), .B1(new_n783_), .B2(G99gat), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n782_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT51), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n788_), .A2(KEYINPUT116), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n787_), .B(new_n789_), .ZN(G1338gat));
  NAND3_X1  g589(.A1(new_n776_), .A2(new_n453_), .A3(new_n501_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n771_), .A2(new_n453_), .A3(new_n772_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n793_));
  AND3_X1   g592(.A1(new_n792_), .A2(new_n793_), .A3(G106gat), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n793_), .B1(new_n792_), .B2(G106gat), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n791_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g596(.A(new_n587_), .ZN(new_n798_));
  OAI211_X1 g597(.A(new_n634_), .B(new_n251_), .C1(new_n798_), .C2(new_n585_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT54), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n799_), .B(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n229_), .A2(new_n230_), .A3(new_n233_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n237_), .A2(new_n231_), .A3(new_n228_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n802_), .A2(KEYINPUT117), .A3(new_n247_), .A4(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n249_), .A2(new_n804_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n803_), .A2(new_n247_), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT117), .B1(new_n806_), .B2(new_n802_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n805_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n577_), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n536_), .B(new_n575_), .C1(new_n564_), .C2(new_n567_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n538_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n568_), .A2(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n563_), .B1(new_n562_), .B2(KEYINPUT12), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n565_), .A2(KEYINPUT72), .A3(new_n566_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n816_), .A2(KEYINPUT55), .A3(new_n536_), .A4(new_n557_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n811_), .A2(new_n813_), .A3(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n578_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT56), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n818_), .A2(KEYINPUT56), .A3(new_n578_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n809_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n695_), .B1(new_n823_), .B2(KEYINPUT58), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n808_), .A2(new_n577_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n822_), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT56), .B1(new_n818_), .B2(new_n578_), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n825_), .B(KEYINPUT58), .C1(new_n826_), .C2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(KEYINPUT118), .B1(new_n824_), .B2(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n825_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT58), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT118), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n833_), .A2(new_n834_), .A3(new_n695_), .A4(new_n828_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n250_), .A2(new_n577_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n836_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n837_));
  AND3_X1   g636(.A1(new_n583_), .A2(new_n584_), .A3(new_n808_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n629_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT57), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  OAI211_X1 g640(.A(KEYINPUT57), .B(new_n629_), .C1(new_n837_), .C2(new_n838_), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n830_), .A2(new_n835_), .A3(new_n841_), .A4(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n801_), .B1(new_n843_), .B2(new_n607_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n475_), .A2(new_n306_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n646_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n844_), .A2(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(G113gat), .B1(new_n847_), .B2(new_n250_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT59), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n846_), .B1(KEYINPUT119), .B2(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n850_), .B1(KEYINPUT119), .B2(new_n846_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n841_), .A2(new_n842_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n833_), .A2(new_n695_), .A3(new_n828_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n651_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n851_), .B1(new_n854_), .B2(new_n801_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n855_), .B1(new_n847_), .B2(new_n849_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n250_), .A2(G113gat), .ZN(new_n858_));
  XOR2_X1   g657(.A(new_n858_), .B(KEYINPUT120), .Z(new_n859_));
  AOI21_X1  g658(.A(new_n848_), .B1(new_n857_), .B2(new_n859_), .ZN(G1340gat));
  OAI21_X1  g659(.A(G120gat), .B1(new_n856_), .B2(new_n588_), .ZN(new_n861_));
  OR2_X1    g660(.A1(new_n844_), .A2(new_n846_), .ZN(new_n862_));
  INV_X1    g661(.A(G120gat), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n863_), .B1(new_n588_), .B2(KEYINPUT60), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n864_), .B1(KEYINPUT60), .B2(new_n863_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n861_), .B1(new_n862_), .B2(new_n865_), .ZN(G1341gat));
  AOI21_X1  g665(.A(G127gat), .B1(new_n847_), .B2(new_n651_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n651_), .A2(G127gat), .ZN(new_n868_));
  XOR2_X1   g667(.A(new_n868_), .B(KEYINPUT121), .Z(new_n869_));
  AOI21_X1  g668(.A(new_n867_), .B1(new_n857_), .B2(new_n869_), .ZN(G1342gat));
  INV_X1    g669(.A(KEYINPUT122), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n844_), .A2(new_n629_), .A3(new_n846_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n871_), .B1(new_n872_), .B2(G134gat), .ZN(new_n873_));
  INV_X1    g672(.A(G134gat), .ZN(new_n874_));
  OAI211_X1 g673(.A(KEYINPUT122), .B(new_n874_), .C1(new_n862_), .C2(new_n629_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n695_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n876_), .A2(new_n874_), .ZN(new_n877_));
  AOI22_X1  g676(.A1(new_n873_), .A2(new_n875_), .B1(new_n857_), .B2(new_n877_), .ZN(G1343gat));
  NOR2_X1   g677(.A1(new_n305_), .A2(new_n476_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n879_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n843_), .A2(new_n607_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n801_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n880_), .B1(new_n881_), .B2(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(new_n250_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n642_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g686(.A(KEYINPUT61), .B(G155gat), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n881_), .A2(new_n882_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n880_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n889_), .A2(new_n651_), .A3(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(KEYINPUT123), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT123), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n883_), .A2(new_n893_), .A3(new_n651_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n888_), .B1(new_n892_), .B2(new_n894_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n893_), .B1(new_n883_), .B2(new_n651_), .ZN(new_n896_));
  NOR4_X1   g695(.A1(new_n844_), .A2(KEYINPUT123), .A3(new_n607_), .A4(new_n880_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n888_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n896_), .A2(new_n897_), .A3(new_n898_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n895_), .A2(new_n899_), .ZN(G1346gat));
  AOI21_X1  g699(.A(G162gat), .B1(new_n883_), .B2(new_n649_), .ZN(new_n901_));
  AND2_X1   g700(.A1(new_n693_), .A2(G162gat), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n901_), .B1(new_n883_), .B2(new_n902_), .ZN(G1347gat));
  NOR2_X1   g702(.A1(new_n854_), .A2(new_n801_), .ZN(new_n904_));
  NOR3_X1   g703(.A1(new_n473_), .A2(new_n306_), .A3(new_n474_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(new_n476_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n904_), .A2(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n311_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n907_), .A2(new_n908_), .A3(new_n250_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n905_), .A2(new_n250_), .ZN(new_n911_));
  XOR2_X1   g710(.A(new_n911_), .B(KEYINPUT124), .Z(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(new_n476_), .ZN(new_n913_));
  OR2_X1    g712(.A1(new_n904_), .A2(new_n913_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n910_), .B1(new_n914_), .B2(G169gat), .ZN(new_n915_));
  OAI211_X1 g714(.A(G169gat), .B(new_n910_), .C1(new_n904_), .C2(new_n913_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n916_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n909_), .B1(new_n915_), .B2(new_n917_), .ZN(G1348gat));
  AOI21_X1  g717(.A(G176gat), .B1(new_n907_), .B2(new_n642_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n844_), .A2(new_n906_), .ZN(new_n920_));
  AND2_X1   g719(.A1(new_n642_), .A2(G176gat), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n919_), .B1(new_n920_), .B2(new_n921_), .ZN(G1349gat));
  AOI21_X1  g721(.A(G183gat), .B1(new_n920_), .B2(new_n651_), .ZN(new_n923_));
  OR2_X1    g722(.A1(new_n607_), .A2(new_n256_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n924_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n923_), .B1(new_n907_), .B2(new_n925_), .ZN(G1350gat));
  NAND3_X1  g725(.A1(new_n907_), .A2(new_n257_), .A3(new_n649_), .ZN(new_n927_));
  NOR3_X1   g726(.A1(new_n904_), .A2(new_n876_), .A3(new_n906_), .ZN(new_n928_));
  INV_X1    g727(.A(G190gat), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n927_), .B1(new_n928_), .B2(new_n929_), .ZN(G1351gat));
  NOR3_X1   g729(.A1(new_n473_), .A2(new_n455_), .A3(new_n305_), .ZN(new_n931_));
  INV_X1    g730(.A(new_n931_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n844_), .A2(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(new_n250_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n934_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g734(.A1(new_n933_), .A2(new_n642_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n330_), .A2(KEYINPUT126), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n936_), .B(new_n937_), .ZN(G1353gat));
  NAND2_X1  g737(.A1(new_n889_), .A2(new_n931_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n940_));
  AND2_X1   g739(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n941_));
  NOR4_X1   g740(.A1(new_n939_), .A2(new_n607_), .A3(new_n940_), .A4(new_n941_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n933_), .A2(new_n651_), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n942_), .B1(new_n943_), .B2(new_n940_), .ZN(G1354gat));
  OAI21_X1  g743(.A(G218gat), .B1(new_n939_), .B2(new_n876_), .ZN(new_n945_));
  NOR4_X1   g744(.A1(new_n844_), .A2(G218gat), .A3(new_n629_), .A4(new_n932_), .ZN(new_n946_));
  INV_X1    g745(.A(new_n946_), .ZN(new_n947_));
  INV_X1    g746(.A(KEYINPUT127), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n945_), .A2(new_n947_), .A3(new_n948_), .ZN(new_n949_));
  INV_X1    g748(.A(G218gat), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n950_), .B1(new_n933_), .B2(new_n695_), .ZN(new_n951_));
  OAI21_X1  g750(.A(KEYINPUT127), .B1(new_n951_), .B2(new_n946_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n949_), .A2(new_n952_), .ZN(G1355gat));
endmodule


