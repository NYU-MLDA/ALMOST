//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 1 0 1 0 0 0 0 1 1 0 1 1 0 1 0 1 1 0 0 1 0 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 1 0 0 0 1 0 0 0 1 0 1 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n677_, new_n678_,
    new_n679_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n687_, new_n688_, new_n689_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n702_, new_n703_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n797_, new_n798_, new_n799_, new_n800_, new_n802_,
    new_n803_, new_n804_, new_n806_, new_n807_, new_n808_, new_n810_,
    new_n811_, new_n813_, new_n814_, new_n816_, new_n817_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n830_, new_n831_, new_n832_,
    new_n834_, new_n836_, new_n837_, new_n839_, new_n840_, new_n842_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n849_, new_n850_,
    new_n851_, new_n852_;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202_));
  INV_X1    g001(.A(G1gat), .ZN(new_n203_));
  INV_X1    g002(.A(G8gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT14), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n202_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G1gat), .B(G8gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT73), .B(KEYINPUT74), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  XOR2_X1   g009(.A(G29gat), .B(G36gat), .Z(new_n211_));
  XOR2_X1   g010(.A(G43gat), .B(G50gat), .Z(new_n212_));
  XNOR2_X1  g011(.A(new_n211_), .B(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n213_), .B(KEYINPUT15), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n210_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT75), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n215_), .B(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n213_), .ZN(new_n218_));
  OR2_X1    g017(.A1(new_n210_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G229gat), .A2(G233gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n217_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n210_), .B(new_n218_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n220_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  AND2_X1   g023(.A1(new_n221_), .A2(new_n224_), .ZN(new_n225_));
  XOR2_X1   g024(.A(G113gat), .B(G141gat), .Z(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT76), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G169gat), .B(G197gat), .ZN(new_n228_));
  XOR2_X1   g027(.A(new_n227_), .B(new_n228_), .Z(new_n229_));
  NOR2_X1   g028(.A1(new_n225_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT77), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n231_), .B1(new_n225_), .B2(new_n229_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n225_), .A2(new_n231_), .A3(new_n229_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n230_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT79), .ZN(new_n236_));
  INV_X1    g035(.A(G169gat), .ZN(new_n237_));
  INV_X1    g036(.A(G176gat), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n236_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(KEYINPUT79), .B1(G169gat), .B2(G176gat), .ZN(new_n240_));
  AOI21_X1  g039(.A(KEYINPUT24), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G183gat), .A2(G190gat), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT23), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT80), .B1(new_n241_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT24), .ZN(new_n246_));
  INV_X1    g045(.A(new_n240_), .ZN(new_n247_));
  NOR3_X1   g046(.A1(KEYINPUT79), .A2(G169gat), .A3(G176gat), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n246_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT80), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n242_), .B(KEYINPUT23), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n249_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G169gat), .A2(G176gat), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n239_), .A2(KEYINPUT24), .A3(new_n253_), .A4(new_n240_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(KEYINPUT25), .B(G183gat), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT78), .ZN(new_n256_));
  INV_X1    g055(.A(G190gat), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n256_), .B1(new_n257_), .B2(KEYINPUT26), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT26), .B(G190gat), .ZN(new_n259_));
  OAI211_X1 g058(.A(new_n255_), .B(new_n258_), .C1(new_n259_), .C2(new_n256_), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n245_), .A2(new_n252_), .A3(new_n254_), .A4(new_n260_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(G183gat), .A2(G190gat), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n262_), .B1(new_n243_), .B2(new_n242_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT22), .B(G169gat), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT81), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(KEYINPUT82), .B(G176gat), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n267_), .B1(new_n237_), .B2(KEYINPUT22), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n265_), .B(new_n253_), .C1(new_n268_), .C2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n261_), .A2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G71gat), .B(G99gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(G43gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n273_), .B(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G227gat), .A2(G233gat), .ZN(new_n277_));
  INV_X1    g076(.A(G15gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT30), .ZN(new_n280_));
  XOR2_X1   g079(.A(new_n276_), .B(new_n280_), .Z(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT85), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT86), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G127gat), .B(G134gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G113gat), .B(G120gat), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT83), .ZN(new_n287_));
  OAI21_X1  g086(.A(KEYINPUT84), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  XOR2_X1   g087(.A(G127gat), .B(G134gat), .Z(new_n289_));
  XOR2_X1   g088(.A(G113gat), .B(G120gat), .Z(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT84), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n291_), .A2(KEYINPUT83), .A3(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n288_), .A2(new_n293_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n289_), .A2(new_n290_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n288_), .A2(new_n293_), .A3(new_n295_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT31), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n300_), .B1(new_n281_), .B2(KEYINPUT85), .ZN(new_n301_));
  OR2_X1    g100(.A1(new_n283_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n283_), .A2(new_n301_), .ZN(new_n303_));
  AND2_X1   g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  XOR2_X1   g103(.A(G1gat), .B(G29gat), .Z(new_n305_));
  XNOR2_X1  g104(.A(G57gat), .B(G85gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G225gat), .A2(G233gat), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G155gat), .A2(G162gat), .ZN(new_n312_));
  NOR2_X1   g111(.A1(G155gat), .A2(G162gat), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(G141gat), .A2(G148gat), .ZN(new_n315_));
  XOR2_X1   g114(.A(new_n315_), .B(KEYINPUT3), .Z(new_n316_));
  NAND2_X1  g115(.A1(G141gat), .A2(G148gat), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n317_), .B(KEYINPUT2), .Z(new_n318_));
  OAI211_X1 g117(.A(new_n312_), .B(new_n314_), .C1(new_n316_), .C2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n317_), .ZN(new_n320_));
  OR2_X1    g119(.A1(new_n320_), .A2(new_n315_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n312_), .B1(new_n313_), .B2(KEYINPUT1), .ZN(new_n322_));
  OR2_X1    g121(.A1(new_n322_), .A2(KEYINPUT87), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n312_), .A2(KEYINPUT1), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n324_), .B1(new_n322_), .B2(KEYINPUT87), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n321_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n326_), .A2(KEYINPUT88), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT88), .ZN(new_n328_));
  AOI211_X1 g127(.A(new_n328_), .B(new_n321_), .C1(new_n323_), .C2(new_n325_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n319_), .B1(new_n327_), .B2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(new_n299_), .ZN(new_n331_));
  OAI221_X1 g130(.A(new_n319_), .B1(new_n295_), .B2(new_n286_), .C1(new_n327_), .C2(new_n329_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n311_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(KEYINPUT4), .B1(new_n330_), .B2(new_n299_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n331_), .A2(new_n332_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n334_), .B1(new_n335_), .B2(KEYINPUT4), .ZN(new_n336_));
  AOI211_X1 g135(.A(new_n309_), .B(new_n333_), .C1(new_n336_), .C2(new_n311_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n309_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n335_), .A2(KEYINPUT4), .ZN(new_n339_));
  INV_X1    g138(.A(new_n334_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n339_), .A2(new_n311_), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n333_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n338_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n337_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G78gat), .B(G106gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(KEYINPUT90), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(G211gat), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n348_), .A2(G218gat), .ZN(new_n349_));
  INV_X1    g148(.A(G218gat), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n350_), .A2(G211gat), .ZN(new_n351_));
  OAI21_X1  g150(.A(KEYINPUT89), .B1(new_n349_), .B2(new_n351_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(G197gat), .A2(G204gat), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G197gat), .A2(G204gat), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n354_), .A2(KEYINPUT21), .A3(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT21), .ZN(new_n357_));
  INV_X1    g156(.A(new_n355_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n357_), .B1(new_n358_), .B2(new_n353_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n350_), .A2(G211gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n348_), .A2(G218gat), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT89), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n360_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n352_), .A2(new_n356_), .A3(new_n359_), .A4(new_n363_), .ZN(new_n364_));
  NOR3_X1   g163(.A1(new_n358_), .A2(new_n353_), .A3(new_n357_), .ZN(new_n365_));
  AND3_X1   g164(.A1(new_n360_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n362_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n365_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  AND2_X1   g167(.A1(new_n364_), .A2(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n369_), .B1(new_n330_), .B2(KEYINPUT29), .ZN(new_n370_));
  INV_X1    g169(.A(G228gat), .ZN(new_n371_));
  INV_X1    g170(.A(G233gat), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n370_), .A2(new_n374_), .ZN(new_n375_));
  AOI211_X1 g174(.A(new_n369_), .B(new_n373_), .C1(new_n330_), .C2(KEYINPUT29), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n347_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT91), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  OR2_X1    g178(.A1(new_n330_), .A2(KEYINPUT29), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G22gat), .B(G50gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT28), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n380_), .B(new_n382_), .ZN(new_n383_));
  OR2_X1    g182(.A1(new_n370_), .A2(new_n374_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n370_), .A2(new_n374_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n384_), .A2(new_n346_), .A3(new_n385_), .ZN(new_n386_));
  AOI22_X1  g185(.A1(new_n379_), .A2(new_n383_), .B1(new_n386_), .B2(new_n377_), .ZN(new_n387_));
  AND4_X1   g186(.A1(KEYINPUT91), .A2(new_n386_), .A3(new_n377_), .A4(new_n383_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n344_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n241_), .A2(new_n244_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n259_), .A2(new_n255_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n390_), .A2(new_n254_), .A3(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n266_), .A2(new_n269_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n253_), .B(KEYINPUT93), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(KEYINPUT94), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT94), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n393_), .A2(new_n394_), .A3(new_n397_), .ZN(new_n398_));
  AND2_X1   g197(.A1(new_n396_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n265_), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n369_), .B(new_n392_), .C1(new_n399_), .C2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n369_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n273_), .A2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n401_), .A2(KEYINPUT20), .A3(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G226gat), .A2(G233gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(KEYINPUT19), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n404_), .A2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n261_), .A2(new_n369_), .A3(new_n272_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(KEYINPUT20), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT92), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n400_), .B1(new_n396_), .B2(new_n398_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n392_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n402_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT92), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n408_), .A2(new_n414_), .A3(KEYINPUT20), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n410_), .A2(new_n413_), .A3(new_n415_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n407_), .B1(new_n416_), .B2(new_n406_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G8gat), .B(G36gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(KEYINPUT18), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G64gat), .B(G92gat), .ZN(new_n420_));
  XOR2_X1   g219(.A(new_n419_), .B(new_n420_), .Z(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n417_), .A2(KEYINPUT101), .A3(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(KEYINPUT101), .B1(new_n417_), .B2(new_n422_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n406_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n401_), .A2(KEYINPUT20), .A3(new_n403_), .A4(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT96), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n427_), .B(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT95), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n415_), .A2(new_n413_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n414_), .B1(new_n408_), .B2(KEYINPUT20), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n430_), .B(new_n406_), .C1(new_n431_), .C2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n430_), .B1(new_n416_), .B2(new_n406_), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n429_), .B(new_n421_), .C1(new_n434_), .C2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT27), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n425_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT97), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n436_), .A2(new_n439_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n406_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT95), .ZN(new_n442_));
  OR2_X1    g241(.A1(new_n427_), .A2(new_n428_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n427_), .A2(new_n428_), .ZN(new_n444_));
  AOI22_X1  g243(.A1(new_n442_), .A2(new_n433_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n445_), .A2(KEYINPUT97), .A3(new_n421_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT98), .ZN(new_n447_));
  NOR3_X1   g246(.A1(new_n445_), .A2(new_n447_), .A3(new_n421_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n429_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n449_));
  AOI21_X1  g248(.A(KEYINPUT98), .B1(new_n449_), .B2(new_n422_), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n440_), .B(new_n446_), .C1(new_n448_), .C2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT27), .ZN(new_n452_));
  AOI211_X1 g251(.A(new_n389_), .B(new_n438_), .C1(new_n451_), .C2(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n387_), .A2(new_n388_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT33), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n343_), .A2(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n333_), .B1(new_n336_), .B2(new_n311_), .ZN(new_n458_));
  OAI21_X1  g257(.A(KEYINPUT33), .B1(new_n458_), .B2(new_n338_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n331_), .A2(new_n311_), .A3(new_n332_), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n460_), .A2(new_n338_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n461_), .B1(new_n336_), .B2(new_n311_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT100), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT100), .ZN(new_n464_));
  OAI211_X1 g263(.A(new_n461_), .B(new_n464_), .C1(new_n336_), .C2(new_n311_), .ZN(new_n465_));
  AOI22_X1  g264(.A1(new_n457_), .A2(new_n459_), .B1(new_n463_), .B2(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n447_), .B1(new_n445_), .B2(new_n421_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n449_), .A2(KEYINPUT98), .A3(new_n422_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n466_), .A2(new_n469_), .A3(new_n440_), .A4(new_n446_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n344_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n417_), .A2(KEYINPUT32), .A3(new_n421_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT32), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n445_), .B1(new_n473_), .B2(new_n422_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n471_), .A2(new_n472_), .A3(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n455_), .B1(new_n470_), .B2(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n304_), .B1(new_n453_), .B2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n302_), .A2(new_n303_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n438_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n478_), .A2(new_n479_), .A3(new_n344_), .A4(new_n454_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n235_), .B1(new_n477_), .B2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G57gat), .B(G64gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT11), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT65), .ZN(new_n484_));
  XOR2_X1   g283(.A(G71gat), .B(G78gat), .Z(new_n485_));
  OAI21_X1  g284(.A(new_n485_), .B1(KEYINPUT11), .B2(new_n482_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n484_), .B(new_n486_), .ZN(new_n487_));
  XOR2_X1   g286(.A(KEYINPUT10), .B(G99gat), .Z(new_n488_));
  INV_X1    g287(.A(G106gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(G85gat), .B(G92gat), .Z(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT9), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G99gat), .A2(G106gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(KEYINPUT6), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT6), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n495_), .A2(G99gat), .A3(G106gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(G85gat), .ZN(new_n498_));
  INV_X1    g297(.A(G92gat), .ZN(new_n499_));
  OR3_X1    g298(.A1(new_n498_), .A2(new_n499_), .A3(KEYINPUT9), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n490_), .A2(new_n492_), .A3(new_n497_), .A4(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT8), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT64), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n497_), .A2(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(G99gat), .A2(G106gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT7), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n494_), .A2(new_n496_), .A3(KEYINPUT64), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n504_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n502_), .B1(new_n508_), .B2(new_n491_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n491_), .A2(new_n502_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n510_), .B1(new_n497_), .B2(new_n506_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n501_), .B1(new_n509_), .B2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n487_), .A2(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n487_), .A2(new_n512_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT12), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n513_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G230gat), .A2(G233gat), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT66), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n512_), .A2(new_n518_), .ZN(new_n519_));
  OAI211_X1 g318(.A(KEYINPUT66), .B(new_n501_), .C1(new_n509_), .C2(new_n511_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n519_), .A2(KEYINPUT12), .A3(new_n487_), .A4(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n516_), .A2(new_n517_), .A3(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n513_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n523_), .A2(new_n514_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n522_), .B1(new_n517_), .B2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G176gat), .B(G204gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT68), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G120gat), .B(G148gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  XOR2_X1   g330(.A(new_n525_), .B(new_n531_), .Z(new_n532_));
  INV_X1    g331(.A(KEYINPUT13), .ZN(new_n533_));
  OR2_X1    g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n532_), .A2(new_n533_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT37), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G232gat), .A2(G233gat), .ZN(new_n538_));
  XOR2_X1   g337(.A(new_n538_), .B(KEYINPUT34), .Z(new_n539_));
  INV_X1    g338(.A(KEYINPUT35), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT70), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n542_), .B1(new_n512_), .B2(new_n218_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n539_), .A2(new_n540_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n519_), .A2(new_n214_), .A3(new_n520_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n543_), .B1(new_n546_), .B2(KEYINPUT69), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT69), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n519_), .A2(new_n549_), .A3(new_n214_), .A4(new_n520_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(KEYINPUT71), .B1(new_n551_), .B2(new_n544_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT71), .ZN(new_n553_));
  INV_X1    g352(.A(new_n544_), .ZN(new_n554_));
  AOI211_X1 g353(.A(new_n553_), .B(new_n554_), .C1(new_n548_), .C2(new_n550_), .ZN(new_n555_));
  OAI211_X1 g354(.A(KEYINPUT72), .B(new_n547_), .C1(new_n552_), .C2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT36), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G190gat), .B(G218gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G134gat), .B(G162gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n556_), .A2(new_n557_), .A3(new_n561_), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n560_), .B(new_n547_), .C1(new_n552_), .C2(new_n555_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n557_), .B1(new_n556_), .B2(new_n561_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n537_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n565_), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n567_), .A2(KEYINPUT37), .A3(new_n563_), .A4(new_n562_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n566_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G231gat), .A2(G233gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n210_), .B(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(new_n487_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G127gat), .B(G155gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT16), .ZN(new_n575_));
  XOR2_X1   g374(.A(G183gat), .B(G211gat), .Z(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT17), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n577_), .A2(new_n578_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n573_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n582_), .B1(new_n580_), .B2(new_n573_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n570_), .A2(new_n583_), .ZN(new_n584_));
  AND3_X1   g383(.A1(new_n481_), .A2(new_n536_), .A3(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n585_), .A2(new_n203_), .A3(new_n471_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT38), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n564_), .A2(new_n565_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n590_), .B1(new_n477_), .B2(new_n480_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n235_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n583_), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n591_), .A2(new_n592_), .A3(new_n536_), .A4(new_n593_), .ZN(new_n594_));
  OAI21_X1  g393(.A(G1gat), .B1(new_n594_), .B2(new_n344_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n586_), .A2(new_n587_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n588_), .A2(new_n595_), .A3(new_n596_), .ZN(G1324gat));
  OAI21_X1  g396(.A(G8gat), .B1(new_n594_), .B2(new_n479_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT39), .ZN(new_n599_));
  INV_X1    g398(.A(new_n479_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n585_), .A2(new_n204_), .A3(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n602_), .B(KEYINPUT40), .Z(G1325gat));
  NAND3_X1  g402(.A1(new_n585_), .A2(new_n278_), .A3(new_n478_), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n604_), .B(KEYINPUT102), .Z(new_n605_));
  OAI21_X1  g404(.A(G15gat), .B1(new_n594_), .B2(new_n304_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(KEYINPUT41), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n606_), .A2(KEYINPUT41), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n605_), .A2(new_n607_), .A3(new_n608_), .ZN(G1326gat));
  OAI21_X1  g408(.A(G22gat), .B1(new_n594_), .B2(new_n454_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT42), .ZN(new_n611_));
  INV_X1    g410(.A(G22gat), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n585_), .A2(new_n612_), .A3(new_n455_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n613_), .ZN(G1327gat));
  NOR2_X1   g413(.A1(new_n589_), .A2(new_n593_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(new_n536_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n481_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(G29gat), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n619_), .A2(new_n620_), .A3(new_n471_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT104), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n536_), .A2(new_n592_), .A3(new_n583_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT103), .ZN(new_n625_));
  AOI221_X4 g424(.A(new_n569_), .B1(new_n625_), .B2(KEYINPUT43), .C1(new_n477_), .C2(new_n480_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n566_), .A2(new_n568_), .A3(KEYINPUT103), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(KEYINPUT43), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n477_), .A2(new_n480_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n628_), .B1(new_n629_), .B2(new_n570_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n624_), .B1(new_n626_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT44), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  OAI211_X1 g432(.A(KEYINPUT44), .B(new_n624_), .C1(new_n626_), .C2(new_n630_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(new_n471_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n622_), .B1(new_n637_), .B2(G29gat), .ZN(new_n638_));
  AOI211_X1 g437(.A(KEYINPUT104), .B(new_n620_), .C1(new_n636_), .C2(new_n471_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n621_), .B1(new_n638_), .B2(new_n639_), .ZN(G1328gat));
  NOR3_X1   g439(.A1(new_n618_), .A2(G36gat), .A3(new_n479_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT107), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n642_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT45), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT106), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT105), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n633_), .A2(new_n648_), .A3(new_n600_), .A4(new_n634_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n649_), .A2(G36gat), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n633_), .A2(new_n600_), .A3(new_n634_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(KEYINPUT105), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n647_), .B1(new_n650_), .B2(new_n652_), .ZN(new_n653_));
  AND4_X1   g452(.A1(new_n647_), .A2(new_n652_), .A3(G36gat), .A4(new_n649_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n646_), .B1(new_n653_), .B2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT46), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  OAI211_X1 g456(.A(KEYINPUT46), .B(new_n646_), .C1(new_n653_), .C2(new_n654_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(G1329gat));
  NAND2_X1  g458(.A1(new_n478_), .A2(G43gat), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n618_), .A2(new_n304_), .ZN(new_n661_));
  OAI22_X1  g460(.A1(new_n635_), .A2(new_n660_), .B1(G43gat), .B2(new_n661_), .ZN(new_n662_));
  XOR2_X1   g461(.A(KEYINPUT108), .B(KEYINPUT47), .Z(new_n663_));
  XNOR2_X1  g462(.A(new_n662_), .B(new_n663_), .ZN(G1330gat));
  AOI21_X1  g463(.A(G50gat), .B1(new_n619_), .B2(new_n455_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n455_), .A2(G50gat), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n665_), .B1(new_n636_), .B2(new_n666_), .ZN(G1331gat));
  NOR2_X1   g466(.A1(new_n536_), .A2(new_n592_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n591_), .A2(new_n593_), .A3(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(G57gat), .ZN(new_n670_));
  NOR3_X1   g469(.A1(new_n669_), .A2(new_n670_), .A3(new_n344_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n629_), .A2(new_n668_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(new_n584_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n344_), .B1(new_n673_), .B2(KEYINPUT109), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n674_), .B1(KEYINPUT109), .B2(new_n673_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n671_), .B1(new_n675_), .B2(new_n670_), .ZN(G1332gat));
  OAI21_X1  g475(.A(G64gat), .B1(new_n669_), .B2(new_n479_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT48), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n479_), .A2(G64gat), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n678_), .B1(new_n673_), .B2(new_n679_), .ZN(G1333gat));
  OAI21_X1  g479(.A(G71gat), .B1(new_n669_), .B2(new_n304_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT49), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n304_), .A2(G71gat), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT110), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n682_), .B1(new_n673_), .B2(new_n684_), .ZN(new_n685_));
  XOR2_X1   g484(.A(new_n685_), .B(KEYINPUT111), .Z(G1334gat));
  OAI21_X1  g485(.A(G78gat), .B1(new_n669_), .B2(new_n454_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT50), .ZN(new_n688_));
  OR2_X1    g487(.A1(new_n454_), .A2(G78gat), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n688_), .B1(new_n673_), .B2(new_n689_), .ZN(G1335gat));
  NAND2_X1  g489(.A1(new_n629_), .A2(new_n570_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n628_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n629_), .A2(new_n570_), .A3(new_n628_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  AND3_X1   g494(.A1(new_n695_), .A2(new_n583_), .A3(new_n668_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(G85gat), .B1(new_n697_), .B2(new_n344_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n672_), .A2(new_n615_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n471_), .A2(new_n498_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n698_), .B1(new_n699_), .B2(new_n700_), .ZN(G1336gat));
  OAI21_X1  g500(.A(G92gat), .B1(new_n697_), .B2(new_n479_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n600_), .A2(new_n499_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n702_), .B1(new_n699_), .B2(new_n703_), .ZN(G1337gat));
  NAND2_X1  g503(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n478_), .A2(new_n488_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n705_), .B1(new_n699_), .B2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n696_), .A2(new_n478_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n707_), .B1(new_n708_), .B2(G99gat), .ZN(new_n709_));
  NOR2_X1   g508(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n709_), .B(new_n710_), .ZN(G1338gat));
  NAND2_X1  g510(.A1(new_n696_), .A2(new_n455_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(G106gat), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n713_), .A2(KEYINPUT113), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT52), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT113), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n716_), .B1(new_n712_), .B2(G106gat), .ZN(new_n717_));
  NOR3_X1   g516(.A1(new_n714_), .A2(new_n715_), .A3(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n455_), .A2(new_n489_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n699_), .A2(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n720_), .B1(new_n717_), .B2(new_n715_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  OAI21_X1  g521(.A(KEYINPUT53), .B1(new_n718_), .B2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT53), .ZN(new_n724_));
  OR2_X1    g523(.A1(new_n717_), .A2(new_n715_), .ZN(new_n725_));
  OAI211_X1 g524(.A(new_n724_), .B(new_n721_), .C1(new_n725_), .C2(new_n714_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n723_), .A2(new_n726_), .ZN(G1339gat));
  NAND4_X1  g526(.A1(new_n479_), .A2(new_n471_), .A3(new_n478_), .A4(new_n454_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n229_), .B1(new_n222_), .B2(new_n220_), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n729_), .A2(KEYINPUT115), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(KEYINPUT115), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n217_), .A2(new_n219_), .A3(new_n223_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n730_), .A2(new_n731_), .A3(new_n732_), .ZN(new_n733_));
  AND3_X1   g532(.A1(new_n225_), .A2(new_n231_), .A3(new_n229_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n733_), .B1(new_n734_), .B2(new_n232_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n735_), .A2(new_n532_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n525_), .A2(new_n531_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n235_), .A2(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n517_), .B1(new_n516_), .B2(new_n521_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT114), .ZN(new_n740_));
  OR2_X1    g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT55), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n522_), .A2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n522_), .A2(new_n742_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n739_), .A2(new_n740_), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n741_), .A2(new_n743_), .A3(new_n744_), .A4(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(new_n531_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT56), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n746_), .A2(KEYINPUT56), .A3(new_n531_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n736_), .B1(new_n738_), .B2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT57), .ZN(new_n753_));
  OR3_X1    g552(.A1(new_n752_), .A2(new_n753_), .A3(new_n590_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT116), .ZN(new_n755_));
  INV_X1    g554(.A(new_n751_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n737_), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n757_), .B(new_n733_), .C1(new_n734_), .C2(new_n232_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n755_), .B1(new_n756_), .B2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(KEYINPUT58), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT58), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n755_), .B(new_n761_), .C1(new_n756_), .C2(new_n758_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n760_), .A2(new_n570_), .A3(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n753_), .B1(new_n752_), .B2(new_n590_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n754_), .A2(new_n763_), .A3(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(new_n583_), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n569_), .A2(new_n235_), .A3(new_n536_), .A4(new_n593_), .ZN(new_n767_));
  OR2_X1    g566(.A1(new_n767_), .A2(KEYINPUT54), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(KEYINPUT54), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n728_), .B1(new_n766_), .B2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(G113gat), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n771_), .A2(new_n772_), .A3(new_n592_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n766_), .A2(new_n770_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n728_), .A2(KEYINPUT119), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n728_), .A2(KEYINPUT119), .ZN(new_n776_));
  XOR2_X1   g575(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n777_));
  NOR3_X1   g576(.A1(new_n775_), .A2(new_n776_), .A3(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n774_), .A2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT59), .ZN(new_n781_));
  OAI21_X1  g580(.A(KEYINPUT117), .B1(new_n771_), .B2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT117), .ZN(new_n783_));
  AOI22_X1  g582(.A1(new_n765_), .A2(new_n583_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n783_), .B(KEYINPUT59), .C1(new_n784_), .C2(new_n728_), .ZN(new_n785_));
  AOI211_X1 g584(.A(KEYINPUT120), .B(new_n780_), .C1(new_n782_), .C2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT120), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n782_), .A2(new_n785_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n787_), .B1(new_n788_), .B2(new_n779_), .ZN(new_n789_));
  NOR3_X1   g588(.A1(new_n786_), .A2(new_n789_), .A3(new_n235_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n773_), .B1(new_n790_), .B2(new_n772_), .ZN(G1340gat));
  INV_X1    g590(.A(G120gat), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n792_), .B1(new_n536_), .B2(KEYINPUT60), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n771_), .B(new_n793_), .C1(KEYINPUT60), .C2(new_n792_), .ZN(new_n794_));
  AOI211_X1 g593(.A(new_n536_), .B(new_n780_), .C1(new_n782_), .C2(new_n785_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n794_), .B1(new_n795_), .B2(new_n792_), .ZN(G1341gat));
  AOI21_X1  g595(.A(G127gat), .B1(new_n771_), .B2(new_n593_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n786_), .A2(new_n789_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n593_), .A2(G127gat), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n799_), .B(KEYINPUT121), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n797_), .B1(new_n798_), .B2(new_n800_), .ZN(G1342gat));
  AOI21_X1  g600(.A(G134gat), .B1(new_n771_), .B2(new_n590_), .ZN(new_n802_));
  XOR2_X1   g601(.A(new_n802_), .B(KEYINPUT122), .Z(new_n803_));
  AND2_X1   g602(.A1(new_n570_), .A2(G134gat), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n803_), .B1(new_n798_), .B2(new_n804_), .ZN(G1343gat));
  NOR4_X1   g604(.A1(new_n600_), .A2(new_n478_), .A3(new_n344_), .A4(new_n454_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n774_), .A2(new_n806_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n807_), .A2(new_n235_), .ZN(new_n808_));
  XOR2_X1   g607(.A(new_n808_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g608(.A1(new_n807_), .A2(new_n536_), .ZN(new_n810_));
  XOR2_X1   g609(.A(KEYINPUT123), .B(G148gat), .Z(new_n811_));
  XNOR2_X1  g610(.A(new_n810_), .B(new_n811_), .ZN(G1345gat));
  NOR2_X1   g611(.A1(new_n807_), .A2(new_n583_), .ZN(new_n813_));
  XOR2_X1   g612(.A(KEYINPUT61), .B(G155gat), .Z(new_n814_));
  XNOR2_X1  g613(.A(new_n813_), .B(new_n814_), .ZN(G1346gat));
  OAI21_X1  g614(.A(G162gat), .B1(new_n807_), .B2(new_n569_), .ZN(new_n816_));
  OR2_X1    g615(.A1(new_n589_), .A2(G162gat), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n816_), .B1(new_n807_), .B2(new_n817_), .ZN(G1347gat));
  NOR3_X1   g617(.A1(new_n304_), .A2(new_n479_), .A3(new_n471_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n819_), .B(KEYINPUT124), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n592_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(KEYINPUT125), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n784_), .A2(new_n455_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n237_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  XOR2_X1   g623(.A(new_n824_), .B(KEYINPUT62), .Z(new_n825_));
  NAND2_X1  g624(.A1(new_n823_), .A2(new_n820_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n827_), .A2(new_n266_), .A3(new_n592_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n825_), .A2(new_n828_), .ZN(G1348gat));
  INV_X1    g628(.A(new_n536_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n827_), .A2(new_n830_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n831_), .A2(new_n238_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n832_), .B1(new_n269_), .B2(new_n831_), .ZN(G1349gat));
  NOR2_X1   g632(.A1(new_n826_), .A2(new_n583_), .ZN(new_n834_));
  MUX2_X1   g633(.A(G183gat), .B(new_n255_), .S(new_n834_), .Z(G1350gat));
  OAI21_X1  g634(.A(G190gat), .B1(new_n826_), .B2(new_n569_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n590_), .A2(new_n259_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n836_), .B1(new_n826_), .B2(new_n837_), .ZN(G1351gat));
  NOR4_X1   g637(.A1(new_n784_), .A2(new_n389_), .A3(new_n479_), .A4(new_n478_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n592_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g640(.A1(new_n839_), .A2(new_n830_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g642(.A1(new_n839_), .A2(new_n593_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n845_));
  AND2_X1   g644(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n846_));
  NOR3_X1   g645(.A1(new_n844_), .A2(new_n845_), .A3(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n847_), .B1(new_n844_), .B2(new_n845_), .ZN(G1354gat));
  XNOR2_X1  g647(.A(KEYINPUT126), .B(G218gat), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n839_), .A2(new_n570_), .A3(new_n849_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n839_), .A2(new_n590_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n850_), .B1(new_n851_), .B2(new_n849_), .ZN(new_n852_));
  XOR2_X1   g651(.A(new_n852_), .B(KEYINPUT127), .Z(G1355gat));
endmodule


