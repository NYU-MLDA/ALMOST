//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 1 0 1 1 0 0 0 0 0 1 0 0 1 0 1 0 1 1 0 1 1 0 0 1 1 0 1 1 0 0 1 1 1 1 0 1 0 0 1 0 0 0 1 1 0 0 1 0 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n689_, new_n690_, new_n691_, new_n692_, new_n694_,
    new_n695_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n745_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n831_,
    new_n832_, new_n834_, new_n835_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n842_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n874_,
    new_n875_, new_n877_, new_n878_, new_n879_, new_n881_, new_n882_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_;
  NAND2_X1  g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202_));
  OR2_X1    g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G141gat), .A2(G148gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT3), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT2), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  OAI211_X1 g008(.A(new_n202_), .B(new_n203_), .C1(new_n206_), .C2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(new_n204_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n202_), .A2(KEYINPUT1), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(new_n203_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n202_), .A2(KEYINPUT1), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n211_), .B(new_n207_), .C1(new_n213_), .C2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n210_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT29), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT85), .ZN(new_n218_));
  XNOR2_X1  g017(.A(G197gat), .B(G204gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT21), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(G197gat), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n222_), .A2(G204gat), .ZN(new_n223_));
  INV_X1    g022(.A(G204gat), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n224_), .A2(G197gat), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT21), .B1(new_n223_), .B2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G211gat), .B(G218gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n221_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  XOR2_X1   g027(.A(G211gat), .B(G218gat), .Z(new_n229_));
  OAI211_X1 g028(.A(new_n229_), .B(KEYINPUT21), .C1(new_n223_), .C2(new_n225_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n217_), .A2(new_n218_), .A3(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G78gat), .B(G106gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT86), .ZN(new_n234_));
  XOR2_X1   g033(.A(new_n232_), .B(new_n234_), .Z(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G22gat), .B(G50gat), .ZN(new_n237_));
  OR3_X1    g036(.A1(new_n216_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n238_));
  OAI21_X1  g037(.A(KEYINPUT28), .B1(new_n216_), .B2(KEYINPUT29), .ZN(new_n239_));
  NAND2_X1  g038(.A1(KEYINPUT84), .A2(G233gat), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(KEYINPUT84), .A2(G233gat), .ZN(new_n242_));
  OAI21_X1  g041(.A(G228gat), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n238_), .A2(new_n239_), .A3(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n244_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n237_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NOR3_X1   g048(.A1(new_n246_), .A2(new_n247_), .A3(new_n237_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n236_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n250_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n252_), .A2(new_n235_), .A3(new_n248_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT101), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT27), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G169gat), .A2(G176gat), .ZN(new_n258_));
  INV_X1    g057(.A(G176gat), .ZN(new_n259_));
  AND2_X1   g058(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n260_));
  NOR2_X1   g059(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n259_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT78), .ZN(new_n263_));
  INV_X1    g062(.A(G183gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(KEYINPUT78), .A2(G183gat), .ZN(new_n266_));
  AOI21_X1  g065(.A(G190gat), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G183gat), .A2(G190gat), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT23), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  OAI211_X1 g071(.A(new_n258_), .B(new_n262_), .C1(new_n267_), .C2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(G190gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT26), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT26), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(G190gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n265_), .A2(KEYINPUT25), .A3(new_n266_), .ZN(new_n279_));
  OR2_X1    g078(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n278_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n271_), .ZN(new_n282_));
  AOI21_X1  g081(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  OR2_X1    g083(.A1(G169gat), .A2(G176gat), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n285_), .A2(KEYINPUT24), .A3(new_n258_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT24), .ZN(new_n287_));
  INV_X1    g086(.A(G169gat), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n287_), .A2(new_n288_), .A3(new_n259_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n284_), .A2(new_n286_), .A3(new_n289_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n273_), .B1(new_n281_), .B2(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT20), .B1(new_n291_), .B2(new_n231_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT88), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G226gat), .A2(G233gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n258_), .A2(KEYINPUT24), .ZN(new_n297_));
  OR2_X1    g096(.A1(new_n297_), .A2(KEYINPUT89), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(KEYINPUT89), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n298_), .A2(new_n299_), .A3(new_n285_), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n284_), .A2(new_n289_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n278_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT25), .B(G183gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n300_), .A2(new_n301_), .A3(new_n304_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n284_), .B1(G183gat), .B2(G190gat), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n306_), .A2(new_n258_), .A3(new_n262_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(new_n231_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT88), .ZN(new_n310_));
  OAI211_X1 g109(.A(new_n310_), .B(KEYINPUT20), .C1(new_n291_), .C2(new_n231_), .ZN(new_n311_));
  NAND4_X1  g110(.A1(new_n293_), .A2(new_n296_), .A3(new_n309_), .A4(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n291_), .A2(new_n231_), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n313_), .B(KEYINPUT20), .C1(new_n308_), .C2(new_n231_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n296_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n312_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G8gat), .B(G36gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT91), .ZN(new_n319_));
  XOR2_X1   g118(.A(KEYINPUT90), .B(KEYINPUT18), .Z(new_n320_));
  OR2_X1    g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n319_), .A2(new_n320_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G64gat), .B(G92gat), .ZN(new_n323_));
  AND3_X1   g122(.A1(new_n321_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n323_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n257_), .B1(new_n317_), .B2(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n293_), .A2(new_n309_), .A3(new_n311_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(new_n315_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n326_), .ZN(new_n330_));
  OR2_X1    g129(.A1(new_n314_), .A2(new_n315_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n329_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n332_));
  AND3_X1   g131(.A1(new_n327_), .A2(KEYINPUT99), .A3(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(KEYINPUT99), .B1(new_n327_), .B2(new_n332_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n332_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n330_), .B1(new_n329_), .B2(new_n331_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n257_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n256_), .B1(new_n335_), .B2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n327_), .A2(new_n332_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT99), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n327_), .A2(KEYINPUT99), .A3(new_n332_), .ZN(new_n343_));
  AND4_X1   g142(.A1(new_n256_), .A2(new_n342_), .A3(new_n338_), .A4(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n255_), .B1(new_n339_), .B2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT102), .ZN(new_n346_));
  AND2_X1   g145(.A1(G127gat), .A2(G134gat), .ZN(new_n347_));
  NOR2_X1   g146(.A1(G127gat), .A2(G134gat), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  AND2_X1   g149(.A1(G113gat), .A2(G120gat), .ZN(new_n351_));
  NOR2_X1   g150(.A1(G113gat), .A2(G120gat), .ZN(new_n352_));
  NOR3_X1   g151(.A1(new_n351_), .A2(new_n352_), .A3(KEYINPUT81), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT81), .ZN(new_n354_));
  OR2_X1    g153(.A1(G113gat), .A2(G120gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G113gat), .A2(G120gat), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n354_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n350_), .B1(new_n353_), .B2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT82), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n355_), .A2(new_n354_), .A3(new_n356_), .ZN(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT81), .B1(new_n351_), .B2(new_n352_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n360_), .A2(new_n361_), .A3(new_n349_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n358_), .A2(new_n359_), .A3(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n349_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(KEYINPUT82), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT4), .ZN(new_n367_));
  AND4_X1   g166(.A1(KEYINPUT92), .A2(new_n366_), .A3(new_n367_), .A4(new_n216_), .ZN(new_n368_));
  AOI22_X1  g167(.A1(new_n363_), .A2(new_n365_), .B1(new_n215_), .B2(new_n210_), .ZN(new_n369_));
  AOI21_X1  g168(.A(KEYINPUT92), .B1(new_n369_), .B2(new_n367_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G225gat), .A2(G233gat), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  AND3_X1   g172(.A1(new_n360_), .A2(new_n361_), .A3(new_n349_), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n210_), .B(new_n215_), .C1(new_n364_), .C2(new_n374_), .ZN(new_n375_));
  AOI211_X1 g174(.A(new_n359_), .B(new_n349_), .C1(new_n361_), .C2(new_n360_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n374_), .A2(new_n364_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n376_), .B1(new_n377_), .B2(new_n359_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n216_), .ZN(new_n379_));
  OAI211_X1 g178(.A(KEYINPUT4), .B(new_n375_), .C1(new_n378_), .C2(new_n379_), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n371_), .A2(KEYINPUT93), .A3(new_n373_), .A4(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G1gat), .B(G29gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT0), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G57gat), .B(G85gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(KEYINPUT94), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n383_), .B(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT95), .B(KEYINPUT96), .ZN(new_n387_));
  XOR2_X1   g186(.A(new_n386_), .B(new_n387_), .Z(new_n388_));
  NAND3_X1  g187(.A1(new_n366_), .A2(new_n367_), .A3(new_n216_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT92), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n369_), .A2(KEYINPUT92), .A3(new_n367_), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n391_), .A2(new_n380_), .A3(new_n373_), .A4(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n375_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n394_), .A2(new_n369_), .ZN(new_n395_));
  AOI21_X1  g194(.A(KEYINPUT93), .B1(new_n395_), .B2(new_n372_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n393_), .A2(new_n396_), .ZN(new_n397_));
  AND3_X1   g196(.A1(new_n381_), .A2(new_n388_), .A3(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n388_), .B1(new_n381_), .B2(new_n397_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n378_), .B(KEYINPUT31), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT80), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  OR2_X1    g202(.A1(new_n403_), .A2(KEYINPUT83), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n401_), .A2(KEYINPUT83), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G227gat), .A2(G233gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n291_), .B(new_n407_), .ZN(new_n408_));
  XOR2_X1   g207(.A(G15gat), .B(G43gat), .Z(new_n409_));
  XNOR2_X1  g208(.A(G71gat), .B(G99gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  XOR2_X1   g210(.A(KEYINPUT79), .B(KEYINPUT30), .Z(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  XOR2_X1   g212(.A(new_n408_), .B(new_n413_), .Z(new_n414_));
  NAND2_X1  g213(.A1(new_n406_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n414_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n404_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n415_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT102), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n419_), .B(new_n255_), .C1(new_n339_), .C2(new_n344_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n346_), .A2(new_n400_), .A3(new_n418_), .A4(new_n420_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n400_), .A2(new_n338_), .A3(new_n343_), .A4(new_n342_), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT100), .B1(new_n422_), .B2(new_n255_), .ZN(new_n423_));
  AND3_X1   g222(.A1(new_n342_), .A2(new_n338_), .A3(new_n343_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT100), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n424_), .A2(new_n254_), .A3(new_n425_), .A4(new_n400_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n423_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n381_), .A2(new_n397_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n388_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT33), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n391_), .A2(new_n380_), .A3(new_n372_), .A4(new_n392_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n395_), .A2(new_n373_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n388_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT97), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n336_), .A2(new_n337_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n399_), .A2(KEYINPUT33), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n432_), .A2(new_n437_), .A3(new_n438_), .A4(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT98), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(KEYINPUT33), .B1(new_n428_), .B2(new_n429_), .ZN(new_n443_));
  AOI211_X1 g242(.A(new_n431_), .B(new_n388_), .C1(new_n381_), .C2(new_n397_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n445_), .A2(KEYINPUT98), .A3(new_n438_), .A4(new_n437_), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n330_), .A2(KEYINPUT32), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(new_n317_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n329_), .A2(new_n331_), .ZN(new_n449_));
  OAI221_X1 g248(.A(new_n448_), .B1(new_n449_), .B2(new_n447_), .C1(new_n398_), .C2(new_n399_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n442_), .A2(new_n446_), .A3(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n427_), .B1(new_n255_), .B2(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n421_), .B1(new_n452_), .B2(new_n418_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  XOR2_X1   g253(.A(G71gat), .B(G78gat), .Z(new_n455_));
  XNOR2_X1  g254(.A(G57gat), .B(G64gat), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n456_), .A2(KEYINPUT11), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n456_), .A2(KEYINPUT11), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n455_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n459_), .B1(new_n457_), .B2(new_n455_), .ZN(new_n460_));
  OR2_X1    g259(.A1(new_n460_), .A2(KEYINPUT64), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(KEYINPUT64), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  XOR2_X1   g262(.A(G85gat), .B(G92gat), .Z(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT9), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G99gat), .A2(G106gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(KEYINPUT6), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n465_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(G85gat), .A2(G92gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT10), .B(G99gat), .ZN(new_n470_));
  OAI221_X1 g269(.A(new_n468_), .B1(KEYINPUT9), .B2(new_n469_), .C1(G106gat), .C2(new_n470_), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n472_));
  OR3_X1    g271(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n467_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(new_n464_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT8), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n463_), .A2(new_n471_), .A3(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n471_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n478_), .A2(new_n462_), .A3(new_n461_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G230gat), .A2(G233gat), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  OR2_X1    g282(.A1(new_n483_), .A2(KEYINPUT65), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(KEYINPUT65), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n478_), .A2(KEYINPUT66), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT66), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n476_), .A2(new_n487_), .A3(new_n471_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n460_), .B(KEYINPUT67), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n489_), .A2(KEYINPUT12), .A3(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT12), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n479_), .A2(new_n492_), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n491_), .A2(new_n481_), .A3(new_n477_), .A4(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n484_), .A2(new_n485_), .A3(new_n494_), .ZN(new_n495_));
  XOR2_X1   g294(.A(G176gat), .B(G204gat), .Z(new_n496_));
  XNOR2_X1  g295(.A(G120gat), .B(G148gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n495_), .A2(new_n501_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n484_), .A2(new_n494_), .A3(new_n485_), .A4(new_n500_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n502_), .A2(KEYINPUT69), .A3(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(KEYINPUT69), .B1(new_n502_), .B2(new_n503_), .ZN(new_n506_));
  OAI21_X1  g305(.A(KEYINPUT13), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n502_), .A2(new_n503_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT69), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT13), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n510_), .A2(new_n511_), .A3(new_n504_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n507_), .A2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G15gat), .B(G22gat), .ZN(new_n514_));
  INV_X1    g313(.A(G1gat), .ZN(new_n515_));
  INV_X1    g314(.A(G8gat), .ZN(new_n516_));
  OAI21_X1  g315(.A(KEYINPUT14), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n514_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G1gat), .B(G8gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G43gat), .B(G50gat), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G29gat), .B(G36gat), .ZN(new_n523_));
  OR2_X1    g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n523_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  XOR2_X1   g325(.A(new_n520_), .B(new_n526_), .Z(new_n527_));
  NAND2_X1  g326(.A1(G229gat), .A2(G233gat), .ZN(new_n528_));
  OR2_X1    g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  XOR2_X1   g328(.A(new_n526_), .B(KEYINPUT15), .Z(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(new_n520_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n531_), .B1(new_n526_), .B2(new_n520_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n528_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n529_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G113gat), .B(G141gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G169gat), .B(G197gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT76), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(new_n534_), .B(new_n539_), .Z(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT77), .ZN(new_n541_));
  NOR3_X1   g340(.A1(new_n454_), .A2(new_n513_), .A3(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G232gat), .A2(G233gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT34), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT35), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n489_), .A2(new_n530_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT70), .ZN(new_n549_));
  OAI22_X1  g348(.A1(new_n478_), .A2(new_n526_), .B1(KEYINPUT35), .B2(new_n544_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n548_), .B1(new_n549_), .B2(new_n551_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n550_), .A2(KEYINPUT70), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n547_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT71), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n547_), .B1(new_n489_), .B2(new_n530_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n555_), .B1(new_n556_), .B2(new_n551_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n556_), .A2(new_n555_), .A3(new_n551_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n554_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  XOR2_X1   g359(.A(G190gat), .B(G218gat), .Z(new_n561_));
  XNOR2_X1  g360(.A(G134gat), .B(G162gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT36), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n563_), .A2(new_n564_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n560_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n559_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n568_), .A2(new_n557_), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n569_), .A2(new_n564_), .A3(new_n563_), .A4(new_n554_), .ZN(new_n570_));
  AND3_X1   g369(.A1(new_n567_), .A2(new_n570_), .A3(KEYINPUT37), .ZN(new_n571_));
  AOI21_X1  g370(.A(KEYINPUT37), .B1(new_n567_), .B2(new_n570_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(G231gat), .A2(G233gat), .ZN(new_n574_));
  XOR2_X1   g373(.A(new_n574_), .B(KEYINPUT72), .Z(new_n575_));
  XOR2_X1   g374(.A(new_n520_), .B(new_n575_), .Z(new_n576_));
  XNOR2_X1  g375(.A(new_n490_), .B(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(G183gat), .B(G211gat), .Z(new_n578_));
  XNOR2_X1  g377(.A(G127gat), .B(G155gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(KEYINPUT17), .ZN(new_n583_));
  OR2_X1    g382(.A1(new_n583_), .A2(KEYINPUT74), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(KEYINPUT74), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n577_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n586_), .B(KEYINPUT75), .Z(new_n587_));
  XNOR2_X1  g386(.A(new_n463_), .B(new_n576_), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n582_), .A2(KEYINPUT17), .ZN(new_n589_));
  AND3_X1   g388(.A1(new_n588_), .A2(new_n583_), .A3(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n587_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n573_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n542_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n400_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n594_), .A2(new_n515_), .A3(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT38), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n567_), .A2(new_n570_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n453_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT103), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n453_), .A2(KEYINPUT103), .A3(new_n598_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n540_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n591_), .ZN(new_n605_));
  NOR3_X1   g404(.A1(new_n513_), .A2(new_n604_), .A3(new_n605_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n603_), .A2(new_n595_), .A3(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n597_), .B1(new_n515_), .B2(new_n607_), .ZN(G1324gat));
  NOR2_X1   g407(.A1(new_n339_), .A2(new_n344_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n602_), .ZN(new_n610_));
  AOI21_X1  g409(.A(KEYINPUT103), .B1(new_n453_), .B2(new_n598_), .ZN(new_n611_));
  OAI211_X1 g410(.A(new_n609_), .B(new_n606_), .C1(new_n610_), .C2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT104), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n603_), .A2(KEYINPUT104), .A3(new_n609_), .A4(new_n606_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n614_), .A2(new_n615_), .A3(G8gat), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(KEYINPUT39), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT39), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n614_), .A2(new_n615_), .A3(new_n618_), .A4(G8gat), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n594_), .A2(new_n516_), .A3(new_n609_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT40), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n620_), .A2(KEYINPUT40), .A3(new_n621_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(G1325gat));
  INV_X1    g425(.A(G15gat), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n594_), .A2(new_n627_), .A3(new_n418_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT105), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n603_), .A2(new_n418_), .A3(new_n606_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(G15gat), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n631_), .A2(KEYINPUT41), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(KEYINPUT41), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n629_), .A2(new_n632_), .A3(new_n633_), .ZN(G1326gat));
  INV_X1    g433(.A(G22gat), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n594_), .A2(new_n635_), .A3(new_n254_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n603_), .A2(new_n254_), .A3(new_n606_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT42), .ZN(new_n638_));
  AND3_X1   g437(.A1(new_n637_), .A2(new_n638_), .A3(G22gat), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n638_), .B1(new_n637_), .B2(G22gat), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n636_), .B1(new_n639_), .B2(new_n640_), .ZN(G1327gat));
  NOR3_X1   g440(.A1(new_n513_), .A2(new_n604_), .A3(new_n591_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n451_), .A2(new_n255_), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n423_), .A2(new_n426_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n418_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  AOI211_X1 g446(.A(KEYINPUT43), .B(new_n573_), .C1(new_n647_), .C2(new_n421_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT43), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n571_), .A2(new_n572_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n649_), .B1(new_n453_), .B2(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n642_), .B1(new_n648_), .B2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(KEYINPUT106), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT44), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT106), .ZN(new_n655_));
  OAI211_X1 g454(.A(new_n655_), .B(new_n642_), .C1(new_n648_), .C2(new_n651_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n653_), .A2(new_n654_), .A3(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n642_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n651_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n453_), .A2(new_n649_), .A3(new_n650_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n658_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(KEYINPUT44), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n657_), .A2(new_n595_), .A3(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(G29gat), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n598_), .A2(new_n591_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n542_), .A2(new_n665_), .ZN(new_n666_));
  OR3_X1    g465(.A1(new_n666_), .A2(G29gat), .A3(new_n400_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n664_), .A2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(KEYINPUT107), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT107), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n664_), .A2(new_n670_), .A3(new_n667_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(G1328gat));
  INV_X1    g471(.A(KEYINPUT108), .ZN(new_n673_));
  INV_X1    g472(.A(G36gat), .ZN(new_n674_));
  INV_X1    g473(.A(new_n609_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n675_), .B1(new_n661_), .B2(KEYINPUT44), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n674_), .B1(new_n657_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n666_), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n678_), .A2(KEYINPUT45), .A3(new_n674_), .A4(new_n609_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT45), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n542_), .A2(new_n674_), .A3(new_n665_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n680_), .B1(new_n681_), .B2(new_n675_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n679_), .A2(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n673_), .B1(new_n677_), .B2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT46), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n673_), .B(KEYINPUT46), .C1(new_n677_), .C2(new_n683_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n686_), .A2(new_n687_), .ZN(G1329gat));
  NOR3_X1   g487(.A1(new_n666_), .A2(G43gat), .A3(new_n646_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n657_), .A2(new_n418_), .A3(new_n662_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n689_), .B1(new_n690_), .B2(G43gat), .ZN(new_n691_));
  XOR2_X1   g490(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n692_));
  XNOR2_X1  g491(.A(new_n691_), .B(new_n692_), .ZN(G1330gat));
  AND4_X1   g492(.A1(G50gat), .A2(new_n657_), .A3(new_n254_), .A4(new_n662_), .ZN(new_n694_));
  AOI21_X1  g493(.A(G50gat), .B1(new_n678_), .B2(new_n254_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n694_), .A2(new_n695_), .ZN(G1331gat));
  INV_X1    g495(.A(new_n513_), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n454_), .A2(new_n540_), .A3(new_n697_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n698_), .A2(new_n593_), .ZN(new_n699_));
  AOI21_X1  g498(.A(G57gat), .B1(new_n699_), .B2(new_n595_), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n603_), .A2(new_n513_), .A3(new_n591_), .A4(new_n541_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT110), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n701_), .B(new_n702_), .ZN(new_n703_));
  XOR2_X1   g502(.A(KEYINPUT111), .B(G57gat), .Z(new_n704_));
  NAND3_X1  g503(.A1(new_n703_), .A2(new_n595_), .A3(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT112), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n703_), .A2(KEYINPUT112), .A3(new_n595_), .A4(new_n704_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n700_), .B1(new_n707_), .B2(new_n708_), .ZN(G1332gat));
  INV_X1    g508(.A(G64gat), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n699_), .A2(new_n710_), .A3(new_n609_), .ZN(new_n711_));
  OR2_X1    g510(.A1(new_n701_), .A2(KEYINPUT110), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n701_), .A2(KEYINPUT110), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n712_), .A2(new_n609_), .A3(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT48), .ZN(new_n715_));
  AND3_X1   g514(.A1(new_n714_), .A2(new_n715_), .A3(G64gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n715_), .B1(new_n714_), .B2(G64gat), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n711_), .B1(new_n716_), .B2(new_n717_), .ZN(G1333gat));
  INV_X1    g517(.A(G71gat), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n699_), .A2(new_n719_), .A3(new_n418_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n712_), .A2(new_n418_), .A3(new_n713_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT49), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n721_), .A2(new_n722_), .A3(G71gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n722_), .B1(new_n721_), .B2(G71gat), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n720_), .B1(new_n723_), .B2(new_n724_), .ZN(G1334gat));
  INV_X1    g524(.A(G78gat), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n699_), .A2(new_n726_), .A3(new_n254_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n712_), .A2(new_n254_), .A3(new_n713_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT50), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n728_), .A2(new_n729_), .A3(G78gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n728_), .B2(G78gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n727_), .B1(new_n730_), .B2(new_n731_), .ZN(G1335gat));
  NAND2_X1  g531(.A1(new_n698_), .A2(new_n665_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(KEYINPUT113), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT113), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n698_), .A2(new_n735_), .A3(new_n665_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(G85gat), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n737_), .A2(new_n738_), .A3(new_n595_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n513_), .A2(new_n604_), .A3(new_n605_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n741_), .A2(new_n595_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n739_), .B1(new_n742_), .B2(new_n738_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT114), .ZN(G1336gat));
  NAND3_X1  g543(.A1(new_n741_), .A2(G92gat), .A3(new_n609_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n675_), .B1(new_n734_), .B2(new_n736_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n745_), .B1(new_n746_), .B2(G92gat), .ZN(new_n747_));
  XOR2_X1   g546(.A(new_n747_), .B(KEYINPUT115), .Z(G1337gat));
  INV_X1    g547(.A(new_n470_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n737_), .A2(new_n418_), .A3(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n741_), .A2(new_n418_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(G99gat), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND2_X1  g553(.A1(new_n741_), .A2(new_n254_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(KEYINPUT116), .A2(KEYINPUT52), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n755_), .A2(G106gat), .A3(new_n756_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(KEYINPUT116), .A2(KEYINPUT52), .ZN(new_n758_));
  OR2_X1    g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(G106gat), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n737_), .A2(new_n760_), .A3(new_n254_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n757_), .A2(new_n758_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n759_), .A2(new_n761_), .A3(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT53), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT53), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n759_), .A2(new_n765_), .A3(new_n761_), .A4(new_n762_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(G1339gat));
  AND3_X1   g566(.A1(new_n346_), .A2(new_n418_), .A3(new_n420_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n598_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT55), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n491_), .A2(new_n477_), .A3(new_n493_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n771_), .B2(new_n482_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n494_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NOR3_X1   g573(.A1(new_n771_), .A2(new_n770_), .A3(new_n482_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n501_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(KEYINPUT56), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT56), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n778_), .B(new_n501_), .C1(new_n774_), .C2(new_n775_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n777_), .A2(new_n540_), .A3(new_n503_), .A4(new_n779_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n534_), .A2(new_n537_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n527_), .A2(new_n528_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n532_), .B(KEYINPUT117), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n782_), .B1(new_n783_), .B2(new_n528_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n781_), .B1(new_n784_), .B2(new_n537_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n510_), .A2(new_n504_), .A3(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n769_), .B1(new_n780_), .B2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT57), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n787_), .B(new_n788_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n777_), .A2(new_n503_), .A3(new_n785_), .A4(new_n779_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT118), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT58), .ZN(new_n792_));
  OR3_X1    g591(.A1(new_n790_), .A2(new_n791_), .A3(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n573_), .B1(new_n792_), .B2(new_n790_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n791_), .B1(new_n790_), .B2(new_n792_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n793_), .A2(new_n794_), .A3(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n591_), .B1(new_n789_), .B2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT54), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n507_), .A2(new_n512_), .A3(new_n541_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n798_), .B1(new_n593_), .B2(new_n800_), .ZN(new_n801_));
  NOR3_X1   g600(.A1(new_n592_), .A2(new_n799_), .A3(KEYINPUT54), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n595_), .B(new_n768_), .C1(new_n797_), .C2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(G113gat), .B1(new_n805_), .B2(new_n540_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(KEYINPUT59), .ZN(new_n807_));
  OR2_X1    g606(.A1(new_n787_), .A2(KEYINPUT57), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n787_), .A2(KEYINPUT57), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n796_), .A2(new_n808_), .A3(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n605_), .ZN(new_n811_));
  OR2_X1    g610(.A1(new_n801_), .A2(new_n802_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT59), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n813_), .A2(new_n814_), .A3(new_n595_), .A4(new_n768_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n807_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(KEYINPUT119), .B(G113gat), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n541_), .A2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n806_), .B1(new_n817_), .B2(new_n819_), .ZN(G1340gat));
  XNOR2_X1  g619(.A(KEYINPUT120), .B(G120gat), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(KEYINPUT60), .B1(new_n513_), .B2(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n513_), .B1(new_n804_), .B2(new_n823_), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n804_), .A2(KEYINPUT60), .A3(new_n823_), .ZN(new_n825_));
  OAI22_X1  g624(.A1(new_n816_), .A2(new_n824_), .B1(new_n825_), .B2(new_n821_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(KEYINPUT121), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT121), .ZN(new_n828_));
  OAI221_X1 g627(.A(new_n828_), .B1(new_n825_), .B2(new_n821_), .C1(new_n816_), .C2(new_n824_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n827_), .A2(new_n829_), .ZN(G1341gat));
  AOI21_X1  g629(.A(G127gat), .B1(new_n805_), .B2(new_n591_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n591_), .A2(G127gat), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n831_), .B1(new_n817_), .B2(new_n832_), .ZN(G1342gat));
  AOI21_X1  g632(.A(G134gat), .B1(new_n805_), .B2(new_n769_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n650_), .A2(G134gat), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n834_), .B1(new_n817_), .B2(new_n835_), .ZN(G1343gat));
  AOI21_X1  g635(.A(new_n400_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n418_), .A2(new_n255_), .ZN(new_n838_));
  AND3_X1   g637(.A1(new_n837_), .A2(new_n675_), .A3(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n540_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g640(.A1(new_n839_), .A2(new_n513_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(G148gat), .ZN(G1345gat));
  NAND4_X1  g642(.A1(new_n837_), .A2(new_n675_), .A3(new_n591_), .A4(new_n838_), .ZN(new_n844_));
  XOR2_X1   g643(.A(KEYINPUT122), .B(KEYINPUT123), .Z(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  AOI211_X1 g645(.A(new_n400_), .B(new_n609_), .C1(new_n811_), .C2(new_n812_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n845_), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n847_), .A2(new_n591_), .A3(new_n838_), .A4(new_n848_), .ZN(new_n849_));
  XOR2_X1   g648(.A(KEYINPUT61), .B(G155gat), .Z(new_n850_));
  AND3_X1   g649(.A1(new_n846_), .A2(new_n849_), .A3(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n850_), .B1(new_n846_), .B2(new_n849_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n851_), .A2(new_n852_), .ZN(G1346gat));
  INV_X1    g652(.A(G162gat), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n854_), .B1(new_n839_), .B2(new_n650_), .ZN(new_n855_));
  AND4_X1   g654(.A1(new_n854_), .A2(new_n847_), .A3(new_n769_), .A4(new_n838_), .ZN(new_n856_));
  OAI21_X1  g655(.A(KEYINPUT124), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n847_), .A2(new_n650_), .A3(new_n838_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(G162gat), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n839_), .A2(new_n854_), .A3(new_n769_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT124), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n859_), .A2(new_n860_), .A3(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n857_), .A2(new_n862_), .ZN(G1347gat));
  AOI21_X1  g662(.A(new_n595_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n675_), .A2(new_n646_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n864_), .A2(new_n255_), .A3(new_n540_), .A4(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(G169gat), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n867_), .A2(KEYINPUT62), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT62), .ZN(new_n869_));
  INV_X1    g668(.A(new_n866_), .ZN(new_n870_));
  OR2_X1    g669(.A1(new_n260_), .A2(new_n261_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n869_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n868_), .B1(new_n872_), .B2(new_n867_), .ZN(G1348gat));
  NAND3_X1  g672(.A1(new_n864_), .A2(new_n255_), .A3(new_n865_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n874_), .A2(new_n697_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(new_n259_), .ZN(G1349gat));
  INV_X1    g675(.A(new_n874_), .ZN(new_n877_));
  AOI22_X1  g676(.A1(new_n877_), .A2(new_n591_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n874_), .A2(new_n303_), .A3(new_n605_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1350gat));
  NAND3_X1  g679(.A1(new_n877_), .A2(new_n302_), .A3(new_n769_), .ZN(new_n881_));
  OAI21_X1  g680(.A(G190gat), .B1(new_n874_), .B2(new_n573_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(G1351gat));
  INV_X1    g682(.A(KEYINPUT125), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n400_), .B(new_n609_), .C1(new_n797_), .C2(new_n803_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n838_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n540_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n884_), .B1(new_n888_), .B2(new_n222_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n222_), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n887_), .A2(KEYINPUT125), .A3(G197gat), .A4(new_n540_), .ZN(new_n891_));
  AND3_X1   g690(.A1(new_n889_), .A2(new_n890_), .A3(new_n891_), .ZN(G1352gat));
  NAND4_X1  g691(.A1(new_n813_), .A2(new_n400_), .A3(new_n609_), .A4(new_n838_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n893_), .A2(new_n697_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(new_n224_), .ZN(G1353gat));
  INV_X1    g694(.A(KEYINPUT63), .ZN(new_n896_));
  INV_X1    g695(.A(G211gat), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT126), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n885_), .A2(new_n605_), .A3(new_n886_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n896_), .A2(new_n897_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n899_), .B1(new_n900_), .B2(new_n902_), .ZN(new_n903_));
  NOR4_X1   g702(.A1(new_n893_), .A2(KEYINPUT126), .A3(new_n605_), .A4(new_n901_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n898_), .B1(new_n903_), .B2(new_n904_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n900_), .A2(new_n899_), .A3(new_n902_), .ZN(new_n906_));
  NAND4_X1  g705(.A1(new_n864_), .A2(new_n609_), .A3(new_n591_), .A4(new_n838_), .ZN(new_n907_));
  OAI21_X1  g706(.A(KEYINPUT126), .B1(new_n907_), .B2(new_n901_), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n906_), .A2(new_n908_), .A3(new_n896_), .A4(new_n897_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n905_), .A2(new_n909_), .ZN(G1354gat));
  INV_X1    g709(.A(KEYINPUT127), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n887_), .A2(new_n911_), .A3(new_n769_), .ZN(new_n912_));
  OAI21_X1  g711(.A(KEYINPUT127), .B1(new_n893_), .B2(new_n598_), .ZN(new_n913_));
  INV_X1    g712(.A(G218gat), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n912_), .A2(new_n913_), .A3(new_n914_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n887_), .A2(G218gat), .A3(new_n650_), .ZN(new_n916_));
  AND2_X1   g715(.A1(new_n915_), .A2(new_n916_), .ZN(G1355gat));
endmodule


