//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 0 1 1 0 0 0 1 0 0 1 0 0 1 1 0 0 0 1 1 1 1 0 0 0 0 1 1 0 0 0 1 0 1 1 1 1 1 1 1 1 0 1 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n676_,
    new_n677_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n705_, new_n706_, new_n707_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n718_,
    new_n719_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n844_, new_n845_, new_n846_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n863_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_, new_n890_, new_n891_, new_n893_,
    new_n894_, new_n895_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n902_, new_n903_, new_n904_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_, new_n922_;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(new_n202_), .B(KEYINPUT11), .Z(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT66), .B(G71gat), .ZN(new_n204_));
  INV_X1    g003(.A(G78gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n203_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n207_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT12), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G99gat), .A2(G106gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT6), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT6), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n215_), .A2(G99gat), .A3(G106gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  OR2_X1    g016(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n218_));
  INV_X1    g017(.A(G106gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(G85gat), .ZN(new_n222_));
  INV_X1    g021(.A(G92gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G85gat), .A2(G92gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(KEYINPUT9), .A3(new_n225_), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n225_), .A2(KEYINPUT9), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n217_), .A2(new_n221_), .A3(new_n226_), .A4(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n228_), .B(KEYINPUT68), .ZN(new_n229_));
  NOR2_X1   g028(.A1(G99gat), .A2(G106gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT64), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT7), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT7), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT64), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n230_), .B1(new_n232_), .B2(new_n234_), .ZN(new_n235_));
  AOI211_X1 g034(.A(G99gat), .B(G106gat), .C1(new_n231_), .C2(KEYINPUT7), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(new_n217_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT8), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n224_), .A2(new_n225_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n238_), .A2(new_n239_), .A3(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(KEYINPUT65), .B1(new_n214_), .B2(new_n216_), .ZN(new_n243_));
  NOR3_X1   g042(.A1(new_n243_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n214_), .A2(new_n216_), .A3(KEYINPUT65), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n240_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n242_), .B1(new_n246_), .B2(new_n239_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT67), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n229_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  OAI211_X1 g048(.A(KEYINPUT67), .B(new_n242_), .C1(new_n246_), .C2(new_n239_), .ZN(new_n250_));
  AOI21_X1  g049(.A(KEYINPUT69), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT65), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n217_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n232_), .A2(new_n234_), .ZN(new_n254_));
  OR2_X1    g053(.A1(G99gat), .A2(G106gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n236_), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n253_), .A2(new_n256_), .A3(new_n257_), .A4(new_n245_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n239_), .B1(new_n258_), .B2(new_n241_), .ZN(new_n259_));
  AOI211_X1 g058(.A(KEYINPUT8), .B(new_n240_), .C1(new_n237_), .C2(new_n217_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n248_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n229_), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n261_), .A2(new_n250_), .A3(KEYINPUT69), .A4(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n212_), .B1(new_n251_), .B2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n247_), .A2(new_n228_), .ZN(new_n266_));
  AOI21_X1  g065(.A(KEYINPUT12), .B1(new_n266_), .B2(new_n210_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n259_), .A2(new_n260_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n228_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n210_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G230gat), .A2(G233gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n265_), .A2(new_n268_), .A3(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT70), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n266_), .A2(new_n210_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n273_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n274_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n261_), .A2(new_n250_), .A3(new_n262_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT69), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(new_n263_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n267_), .B1(new_n286_), .B2(new_n212_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT70), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n287_), .A2(new_n288_), .A3(new_n276_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n278_), .A2(new_n282_), .A3(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G120gat), .B(G148gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT5), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G176gat), .B(G204gat), .ZN(new_n293_));
  XOR2_X1   g092(.A(new_n292_), .B(new_n293_), .Z(new_n294_));
  NAND2_X1  g093(.A1(new_n290_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n294_), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n278_), .A2(new_n282_), .A3(new_n289_), .A4(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT71), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT72), .ZN(new_n299_));
  AND3_X1   g098(.A1(new_n297_), .A2(new_n298_), .A3(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n299_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n295_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n297_), .A2(new_n298_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT72), .ZN(new_n304_));
  INV_X1    g103(.A(new_n295_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n297_), .A2(new_n298_), .A3(new_n299_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n304_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n302_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT13), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n302_), .A2(new_n307_), .A3(KEYINPUT13), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT73), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n310_), .A2(KEYINPUT73), .A3(new_n311_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT23), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n318_), .A2(G183gat), .A3(G190gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT81), .ZN(new_n320_));
  INV_X1    g119(.A(G183gat), .ZN(new_n321_));
  INV_X1    g120(.A(G190gat), .ZN(new_n322_));
  OAI21_X1  g121(.A(KEYINPUT23), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n320_), .A2(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(G169gat), .A2(G176gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT80), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT24), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT26), .B(G190gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT25), .B(G183gat), .ZN(new_n329_));
  AOI22_X1  g128(.A1(new_n326_), .A2(new_n327_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n326_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G169gat), .A2(G176gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n324_), .B(new_n330_), .C1(new_n333_), .C2(new_n327_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(KEYINPUT22), .B(G169gat), .ZN(new_n335_));
  INV_X1    g134(.A(G176gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  OR2_X1    g136(.A1(new_n337_), .A2(KEYINPUT82), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n323_), .A2(new_n319_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n339_), .B1(G183gat), .B2(G190gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n337_), .A2(KEYINPUT82), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n338_), .A2(new_n332_), .A3(new_n340_), .A4(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n334_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT83), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G15gat), .B(G43gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT84), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(G71gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(G99gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n345_), .B(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  XOR2_X1   g150(.A(G127gat), .B(G134gat), .Z(new_n352_));
  XOR2_X1   g151(.A(G113gat), .B(G120gat), .Z(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  XOR2_X1   g153(.A(new_n354_), .B(KEYINPUT87), .Z(new_n355_));
  INV_X1    g154(.A(KEYINPUT31), .ZN(new_n356_));
  AOI21_X1  g155(.A(KEYINPUT86), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n357_), .B1(new_n356_), .B2(new_n355_), .ZN(new_n358_));
  OR2_X1    g157(.A1(new_n358_), .A2(KEYINPUT88), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(KEYINPUT88), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G227gat), .A2(G233gat), .ZN(new_n361_));
  XOR2_X1   g160(.A(new_n361_), .B(KEYINPUT85), .Z(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT30), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n359_), .A2(new_n360_), .A3(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n364_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n351_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n367_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n369_), .A2(new_n350_), .A3(new_n365_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G226gat), .A2(G233gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT19), .ZN(new_n374_));
  XOR2_X1   g173(.A(KEYINPUT97), .B(KEYINPUT24), .Z(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(new_n325_), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n339_), .B(new_n376_), .C1(new_n333_), .C2(new_n375_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n329_), .B(KEYINPUT96), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n377_), .B1(new_n328_), .B2(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n324_), .B1(G183gat), .B2(G190gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n335_), .B(KEYINPUT98), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(new_n336_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n380_), .A2(new_n332_), .A3(new_n382_), .ZN(new_n383_));
  OR2_X1    g182(.A1(new_n383_), .A2(KEYINPUT99), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(KEYINPUT99), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n379_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  XOR2_X1   g185(.A(KEYINPUT92), .B(G204gat), .Z(new_n387_));
  XOR2_X1   g186(.A(KEYINPUT91), .B(G197gat), .Z(new_n388_));
  AOI22_X1  g187(.A1(G197gat), .A2(new_n387_), .B1(new_n388_), .B2(G204gat), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT21), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G211gat), .B(G218gat), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n388_), .A2(G204gat), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n387_), .A2(G197gat), .ZN(new_n394_));
  OAI21_X1  g193(.A(KEYINPUT21), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT93), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n395_), .A2(new_n396_), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n391_), .B(new_n392_), .C1(new_n397_), .C2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT94), .ZN(new_n400_));
  AOI211_X1 g199(.A(new_n390_), .B(new_n392_), .C1(new_n389_), .C2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n401_), .B1(new_n400_), .B2(new_n389_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n399_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(KEYINPUT20), .B1(new_n386_), .B2(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n345_), .A2(new_n403_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n374_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G8gat), .B(G36gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT18), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G64gat), .B(G92gat), .ZN(new_n410_));
  XOR2_X1   g209(.A(new_n409_), .B(new_n410_), .Z(new_n411_));
  NAND2_X1  g210(.A1(new_n386_), .A2(new_n404_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n345_), .A2(new_n403_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n374_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n412_), .A2(KEYINPUT20), .A3(new_n413_), .A4(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n407_), .A2(new_n411_), .A3(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT100), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT100), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n407_), .A2(new_n418_), .A3(new_n411_), .A4(new_n415_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n407_), .A2(new_n415_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n411_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n417_), .A2(new_n419_), .A3(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G1gat), .B(G29gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(new_n222_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(KEYINPUT0), .B(G57gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n425_), .B(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G225gat), .A2(G233gat), .ZN(new_n428_));
  NOR2_X1   g227(.A1(G155gat), .A2(G162gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(KEYINPUT89), .ZN(new_n430_));
  NAND2_X1  g229(.A1(G155gat), .A2(G162gat), .ZN(new_n431_));
  INV_X1    g230(.A(G141gat), .ZN(new_n432_));
  INV_X1    g231(.A(G148gat), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT3), .ZN(new_n435_));
  NOR2_X1   g234(.A1(G141gat), .A2(G148gat), .ZN(new_n436_));
  AOI22_X1  g235(.A1(new_n434_), .A2(KEYINPUT2), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n437_), .B1(KEYINPUT2), .B2(new_n434_), .ZN(new_n438_));
  OAI21_X1  g237(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(KEYINPUT90), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n430_), .B(new_n431_), .C1(new_n438_), .C2(new_n440_), .ZN(new_n441_));
  XOR2_X1   g240(.A(new_n431_), .B(KEYINPUT1), .Z(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(new_n430_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n434_), .A2(new_n436_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n441_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n354_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n448_), .A2(KEYINPUT4), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n441_), .A2(new_n354_), .A3(new_n445_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n448_), .A2(KEYINPUT4), .A3(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n449_), .B1(KEYINPUT101), .B2(new_n451_), .ZN(new_n452_));
  AND2_X1   g251(.A1(new_n448_), .A2(new_n450_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT101), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n453_), .A2(new_n454_), .A3(KEYINPUT4), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n428_), .B1(new_n452_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n428_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n453_), .A2(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n427_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n452_), .A2(new_n455_), .A3(new_n428_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n427_), .B1(new_n453_), .B2(new_n457_), .ZN(new_n461_));
  AND2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT33), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n459_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n464_), .B1(new_n463_), .B2(new_n459_), .ZN(new_n465_));
  OR3_X1    g264(.A1(new_n456_), .A2(new_n427_), .A3(new_n458_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT102), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n466_), .A2(new_n459_), .A3(new_n467_), .ZN(new_n468_));
  OAI211_X1 g267(.A(KEYINPUT102), .B(new_n427_), .C1(new_n456_), .C2(new_n458_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n411_), .A2(KEYINPUT32), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n407_), .A2(new_n471_), .A3(new_n415_), .ZN(new_n472_));
  NOR3_X1   g271(.A1(new_n405_), .A2(new_n374_), .A3(new_n406_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT20), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n382_), .A2(new_n332_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n379_), .B1(new_n380_), .B2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n474_), .B1(new_n404_), .B2(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n414_), .B1(new_n477_), .B2(new_n413_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n473_), .A2(new_n478_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n472_), .B1(new_n479_), .B2(new_n471_), .ZN(new_n480_));
  OAI22_X1  g279(.A1(new_n423_), .A2(new_n465_), .B1(new_n470_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G228gat), .A2(G233gat), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT29), .ZN(new_n483_));
  INV_X1    g282(.A(new_n446_), .ZN(new_n484_));
  OAI211_X1 g283(.A(new_n403_), .B(new_n482_), .C1(new_n483_), .C2(new_n484_), .ZN(new_n485_));
  XOR2_X1   g284(.A(KEYINPUT95), .B(KEYINPUT29), .Z(new_n486_));
  AOI22_X1  g285(.A1(new_n399_), .A2(new_n402_), .B1(new_n446_), .B2(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n485_), .B1(new_n487_), .B2(new_n482_), .ZN(new_n488_));
  XOR2_X1   g287(.A(G78gat), .B(G106gat), .Z(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n489_), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n485_), .B(new_n491_), .C1(new_n487_), .C2(new_n482_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n484_), .A2(new_n483_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT28), .ZN(new_n495_));
  XOR2_X1   g294(.A(G22gat), .B(G50gat), .Z(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n493_), .A2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n497_), .A2(new_n490_), .A3(new_n492_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n481_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT27), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n423_), .A2(new_n504_), .ZN(new_n505_));
  AND2_X1   g304(.A1(new_n416_), .A2(KEYINPUT27), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n421_), .B1(new_n473_), .B2(new_n478_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  AOI22_X1  g307(.A1(new_n469_), .A2(new_n468_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n505_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n372_), .B1(new_n503_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n470_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n512_), .A2(new_n371_), .ZN(new_n513_));
  AOI22_X1  g312(.A1(new_n423_), .A2(new_n504_), .B1(new_n507_), .B2(new_n506_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n513_), .A2(new_n514_), .A3(new_n502_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n511_), .A2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G29gat), .B(G36gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G43gat), .B(G50gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT15), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n286_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G232gat), .A2(G233gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT34), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT35), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n271_), .A2(new_n520_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT75), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n530_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n529_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n522_), .A2(new_n528_), .A3(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n521_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n535_), .B1(new_n285_), .B2(new_n263_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n527_), .B1(new_n536_), .B2(new_n532_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n534_), .A2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G190gat), .B(G218gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT74), .ZN(new_n540_));
  XOR2_X1   g339(.A(G134gat), .B(G162gat), .Z(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n543_), .A2(KEYINPUT36), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n538_), .A2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n534_), .A2(new_n544_), .A3(new_n537_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n543_), .A2(KEYINPUT36), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n547_), .A2(KEYINPUT76), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(KEYINPUT37), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n548_), .A2(KEYINPUT37), .A3(new_n549_), .A4(new_n551_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G127gat), .B(G155gat), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT16), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G183gat), .B(G211gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT17), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT77), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G15gat), .B(G22gat), .ZN(new_n565_));
  INV_X1    g364(.A(G1gat), .ZN(new_n566_));
  INV_X1    g365(.A(G8gat), .ZN(new_n567_));
  OAI21_X1  g366(.A(KEYINPUT14), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n565_), .A2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G1gat), .B(G8gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G231gat), .A2(G233gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n272_), .B(new_n573_), .ZN(new_n574_));
  AND2_X1   g373(.A1(new_n564_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(KEYINPUT78), .ZN(new_n576_));
  INV_X1    g375(.A(new_n561_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(KEYINPUT17), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n576_), .B1(new_n574_), .B2(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n575_), .A2(KEYINPUT78), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n556_), .A2(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n571_), .B(new_n520_), .Z(new_n583_));
  NAND2_X1  g382(.A1(G229gat), .A2(G233gat), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n521_), .A2(new_n571_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n571_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n588_), .A2(new_n520_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n587_), .A2(new_n589_), .A3(new_n584_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n586_), .A2(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G113gat), .B(G141gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G169gat), .B(G197gat), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n592_), .B(new_n593_), .Z(new_n594_));
  OR2_X1    g393(.A1(new_n594_), .A2(KEYINPUT79), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n591_), .B(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n582_), .A2(new_n597_), .ZN(new_n598_));
  NOR3_X1   g397(.A1(new_n317_), .A2(new_n517_), .A3(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n599_), .A2(new_n566_), .A3(new_n512_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT38), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  AOI22_X1  g401(.A1(new_n481_), .A2(new_n502_), .B1(new_n514_), .B2(new_n509_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n515_), .B1(new_n603_), .B2(new_n372_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n581_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n550_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n604_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n312_), .A2(new_n596_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(G1gat), .B1(new_n610_), .B2(new_n470_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n600_), .A2(new_n601_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n602_), .A2(new_n611_), .A3(new_n612_), .ZN(G1324gat));
  NOR2_X1   g412(.A1(new_n610_), .A2(new_n514_), .ZN(new_n614_));
  OR3_X1    g413(.A1(new_n614_), .A2(KEYINPUT39), .A3(new_n567_), .ZN(new_n615_));
  OAI21_X1  g414(.A(KEYINPUT39), .B1(new_n614_), .B2(new_n567_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n514_), .A2(G8gat), .ZN(new_n617_));
  AOI22_X1  g416(.A1(new_n615_), .A2(new_n616_), .B1(new_n599_), .B2(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n618_), .B(new_n620_), .ZN(G1325gat));
  INV_X1    g420(.A(G15gat), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n599_), .A2(new_n622_), .A3(new_n372_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n608_), .A2(new_n372_), .A3(new_n609_), .ZN(new_n624_));
  AND3_X1   g423(.A1(new_n624_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n625_));
  AOI21_X1  g424(.A(KEYINPUT41), .B1(new_n624_), .B2(G15gat), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n623_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT104), .ZN(G1326gat));
  XNOR2_X1  g427(.A(new_n501_), .B(KEYINPUT105), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(G22gat), .B1(new_n610_), .B2(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT42), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n630_), .A2(G22gat), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n633_), .B(KEYINPUT106), .Z(new_n634_));
  NAND2_X1  g433(.A1(new_n599_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n632_), .A2(new_n635_), .ZN(G1327gat));
  NAND2_X1  g435(.A1(new_n609_), .A2(new_n581_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n604_), .A2(new_n550_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  AOI21_X1  g438(.A(G29gat), .B1(new_n639_), .B2(new_n512_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(KEYINPUT108), .B(KEYINPUT44), .ZN(new_n641_));
  XNOR2_X1  g440(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n642_), .B1(new_n604_), .B2(new_n556_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n517_), .A2(new_n555_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT107), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(KEYINPUT43), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n643_), .B1(new_n644_), .B2(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n641_), .B1(new_n647_), .B2(new_n637_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n604_), .A2(new_n556_), .A3(new_n646_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n649_), .B1(new_n644_), .B2(new_n642_), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n650_), .A2(KEYINPUT44), .A3(new_n581_), .A4(new_n609_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n648_), .A2(new_n651_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n512_), .A2(G29gat), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n640_), .B1(new_n652_), .B2(new_n653_), .ZN(G1328gat));
  INV_X1    g453(.A(new_n514_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n648_), .A2(new_n655_), .A3(new_n651_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(G36gat), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n514_), .A2(G36gat), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n639_), .A2(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT45), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n657_), .A2(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(KEYINPUT46), .B1(new_n661_), .B2(KEYINPUT109), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT109), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT46), .ZN(new_n664_));
  AOI211_X1 g463(.A(new_n663_), .B(new_n664_), .C1(new_n657_), .C2(new_n660_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n662_), .A2(new_n665_), .ZN(G1329gat));
  NAND3_X1  g465(.A1(new_n652_), .A2(G43gat), .A3(new_n372_), .ZN(new_n667_));
  INV_X1    g466(.A(G43gat), .ZN(new_n668_));
  INV_X1    g467(.A(new_n639_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n668_), .B1(new_n669_), .B2(new_n371_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n667_), .A2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(KEYINPUT47), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT47), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n667_), .A2(new_n673_), .A3(new_n670_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n672_), .A2(new_n674_), .ZN(G1330gat));
  AOI21_X1  g474(.A(G50gat), .B1(new_n639_), .B2(new_n629_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n501_), .A2(G50gat), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n676_), .B1(new_n652_), .B2(new_n677_), .ZN(G1331gat));
  NAND3_X1  g477(.A1(new_n317_), .A2(new_n596_), .A3(new_n608_), .ZN(new_n679_));
  OAI21_X1  g478(.A(G57gat), .B1(new_n679_), .B2(new_n470_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n312_), .A2(new_n582_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT110), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n683_), .A2(new_n604_), .A3(new_n596_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n681_), .A2(new_n682_), .ZN(new_n685_));
  OR3_X1    g484(.A1(new_n684_), .A2(KEYINPUT111), .A3(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(KEYINPUT111), .B1(new_n684_), .B2(new_n685_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  OR2_X1    g487(.A1(new_n470_), .A2(G57gat), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n680_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT112), .ZN(G1332gat));
  OR2_X1    g490(.A1(new_n679_), .A2(new_n514_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT48), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n692_), .A2(new_n693_), .A3(G64gat), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n693_), .B1(new_n692_), .B2(G64gat), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n514_), .A2(G64gat), .ZN(new_n697_));
  OAI22_X1  g496(.A1(new_n695_), .A2(new_n696_), .B1(new_n688_), .B2(new_n697_), .ZN(G1333gat));
  OAI21_X1  g497(.A(G71gat), .B1(new_n679_), .B2(new_n371_), .ZN(new_n699_));
  OR2_X1    g498(.A1(new_n699_), .A2(KEYINPUT49), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n699_), .A2(KEYINPUT49), .ZN(new_n702_));
  OR2_X1    g501(.A1(new_n371_), .A2(G71gat), .ZN(new_n703_));
  OAI22_X1  g502(.A1(new_n701_), .A2(new_n702_), .B1(new_n688_), .B2(new_n703_), .ZN(G1334gat));
  OAI21_X1  g503(.A(G78gat), .B1(new_n679_), .B2(new_n630_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT50), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n629_), .A2(new_n205_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n706_), .B1(new_n688_), .B2(new_n707_), .ZN(G1335gat));
  NOR2_X1   g507(.A1(new_n605_), .A2(new_n597_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n650_), .A2(new_n312_), .A3(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(G85gat), .B1(new_n710_), .B2(new_n470_), .ZN(new_n711_));
  OAI211_X1 g510(.A(new_n581_), .B(new_n550_), .C1(new_n511_), .C2(new_n516_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n713_), .A2(new_n315_), .A3(new_n314_), .A4(new_n596_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT113), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n512_), .A2(new_n222_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n711_), .B1(new_n715_), .B2(new_n716_), .ZN(G1336gat));
  OAI21_X1  g516(.A(G92gat), .B1(new_n710_), .B2(new_n514_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n655_), .A2(new_n223_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n718_), .B1(new_n715_), .B2(new_n719_), .ZN(G1337gat));
  NAND3_X1  g519(.A1(new_n372_), .A2(new_n218_), .A3(new_n220_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT113), .ZN(new_n722_));
  OR2_X1    g521(.A1(new_n714_), .A2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n714_), .A2(new_n722_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n721_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n650_), .A2(new_n312_), .A3(new_n372_), .A4(new_n709_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n726_), .A2(G99gat), .ZN(new_n727_));
  OAI21_X1  g526(.A(KEYINPUT115), .B1(new_n725_), .B2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT115), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n726_), .A2(G99gat), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n729_), .B(new_n730_), .C1(new_n715_), .C2(new_n721_), .ZN(new_n731_));
  AND2_X1   g530(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n732_));
  AND3_X1   g531(.A1(new_n728_), .A2(new_n731_), .A3(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n728_), .B2(new_n731_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n733_), .A2(new_n734_), .ZN(G1338gat));
  NAND4_X1  g534(.A1(new_n650_), .A2(new_n312_), .A3(new_n501_), .A4(new_n709_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT52), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n736_), .A2(new_n737_), .A3(G106gat), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n737_), .B1(new_n736_), .B2(G106gat), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n501_), .A2(new_n219_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n715_), .A2(new_n741_), .ZN(new_n742_));
  OR3_X1    g541(.A1(new_n740_), .A2(KEYINPUT53), .A3(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(KEYINPUT53), .B1(new_n740_), .B2(new_n742_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(G1339gat));
  INV_X1    g544(.A(G113gat), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n596_), .A2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT117), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n583_), .A2(new_n584_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n587_), .A2(new_n589_), .A3(new_n585_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n594_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(new_n594_), .B2(new_n591_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n288_), .B1(new_n287_), .B2(new_n276_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n211_), .B1(new_n285_), .B2(new_n263_), .ZN(new_n755_));
  NOR4_X1   g554(.A1(new_n755_), .A2(KEYINPUT70), .A3(new_n275_), .A4(new_n267_), .ZN(new_n756_));
  NOR3_X1   g555(.A1(new_n754_), .A2(new_n756_), .A3(KEYINPUT55), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n287_), .A2(new_n273_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(new_n281_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n755_), .A2(new_n267_), .A3(new_n275_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT55), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n294_), .B1(new_n757_), .B2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT56), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  OAI211_X1 g564(.A(KEYINPUT56), .B(new_n294_), .C1(new_n757_), .C2(new_n762_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n765_), .A2(KEYINPUT116), .A3(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n297_), .A2(new_n597_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n278_), .A2(new_n769_), .A3(new_n289_), .ZN(new_n770_));
  AOI22_X1  g569(.A1(new_n758_), .A2(new_n281_), .B1(new_n760_), .B2(KEYINPUT55), .ZN(new_n771_));
  AOI211_X1 g570(.A(new_n764_), .B(new_n296_), .C1(new_n770_), .C2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT116), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n768_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  AOI22_X1  g573(.A1(new_n308_), .A2(new_n753_), .B1(new_n767_), .B2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT57), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n550_), .A2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n748_), .B1(new_n775_), .B2(new_n778_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n767_), .A2(new_n774_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n752_), .B1(new_n302_), .B2(new_n307_), .ZN(new_n781_));
  OAI211_X1 g580(.A(KEYINPUT117), .B(new_n777_), .C1(new_n780_), .C2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n779_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n765_), .A2(new_n766_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n297_), .A2(new_n753_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT58), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n784_), .A2(KEYINPUT58), .A3(new_n785_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n788_), .A2(new_n556_), .A3(new_n789_), .ZN(new_n790_));
  NOR3_X1   g589(.A1(new_n300_), .A2(new_n301_), .A3(new_n295_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n305_), .B1(new_n304_), .B2(new_n306_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n753_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n767_), .A2(new_n774_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n550_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n790_), .B1(new_n795_), .B2(KEYINPUT57), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n581_), .B1(new_n783_), .B2(new_n796_), .ZN(new_n797_));
  AOI211_X1 g596(.A(new_n597_), .B(new_n581_), .C1(new_n553_), .C2(new_n554_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n310_), .A2(new_n311_), .A3(new_n798_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n799_), .B(KEYINPUT54), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n797_), .A2(new_n800_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n655_), .A2(new_n501_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n802_), .A2(new_n512_), .A3(new_n372_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(KEYINPUT59), .B1(new_n801_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT59), .ZN(new_n806_));
  AOI211_X1 g605(.A(new_n806_), .B(new_n803_), .C1(new_n797_), .C2(new_n800_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n747_), .B1(new_n805_), .B2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n803_), .B1(new_n797_), .B2(new_n800_), .ZN(new_n809_));
  AOI211_X1 g608(.A(KEYINPUT118), .B(G113gat), .C1(new_n809_), .C2(new_n597_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT118), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n793_), .A2(new_n794_), .ZN(new_n812_));
  AOI21_X1  g611(.A(KEYINPUT117), .B1(new_n812_), .B2(new_n777_), .ZN(new_n813_));
  AOI211_X1 g612(.A(new_n748_), .B(new_n778_), .C1(new_n793_), .C2(new_n794_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n606_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n555_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n817_));
  AOI22_X1  g616(.A1(new_n816_), .A2(new_n776_), .B1(new_n789_), .B2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n605_), .B1(new_n815_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n799_), .B(new_n820_), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n597_), .B(new_n804_), .C1(new_n819_), .C2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n811_), .B1(new_n822_), .B2(new_n746_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n808_), .B1(new_n810_), .B2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(KEYINPUT119), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT119), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n808_), .B(new_n826_), .C1(new_n810_), .C2(new_n823_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n825_), .A2(new_n827_), .ZN(G1340gat));
  OAI21_X1  g627(.A(new_n776_), .B1(new_n775_), .B2(new_n550_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n829_), .A2(new_n779_), .A3(new_n790_), .A4(new_n782_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n821_), .B1(new_n581_), .B2(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n806_), .B1(new_n831_), .B2(new_n803_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n801_), .A2(KEYINPUT59), .A3(new_n804_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(G120gat), .B1(new_n835_), .B2(new_n316_), .ZN(new_n836_));
  INV_X1    g635(.A(G120gat), .ZN(new_n837_));
  INV_X1    g636(.A(new_n312_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n837_), .B1(new_n838_), .B2(KEYINPUT60), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n809_), .B(new_n839_), .C1(KEYINPUT60), .C2(new_n837_), .ZN(new_n840_));
  AND2_X1   g639(.A1(new_n840_), .A2(KEYINPUT120), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n840_), .A2(KEYINPUT120), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n836_), .B1(new_n841_), .B2(new_n842_), .ZN(G1341gat));
  OAI21_X1  g642(.A(G127gat), .B1(new_n835_), .B2(new_n581_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n809_), .ZN(new_n845_));
  OR3_X1    g644(.A1(new_n845_), .A2(G127gat), .A3(new_n581_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n846_), .ZN(G1342gat));
  INV_X1    g646(.A(KEYINPUT121), .ZN(new_n848_));
  INV_X1    g647(.A(G134gat), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n849_), .B1(new_n834_), .B2(new_n556_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n550_), .A2(new_n849_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n845_), .A2(new_n851_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n848_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n555_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n854_));
  OAI221_X1 g653(.A(KEYINPUT121), .B1(new_n845_), .B2(new_n851_), .C1(new_n854_), .C2(new_n849_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n853_), .A2(new_n855_), .ZN(G1343gat));
  NOR2_X1   g655(.A1(new_n372_), .A2(new_n502_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n801_), .A2(new_n857_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n655_), .A2(new_n470_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n860_), .A2(new_n596_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(new_n432_), .ZN(G1344gat));
  NOR2_X1   g661(.A1(new_n860_), .A2(new_n316_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(new_n433_), .ZN(G1345gat));
  NAND4_X1  g663(.A1(new_n801_), .A2(new_n605_), .A3(new_n857_), .A4(new_n859_), .ZN(new_n865_));
  OR2_X1    g664(.A1(new_n865_), .A2(KEYINPUT122), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(KEYINPUT122), .ZN(new_n867_));
  XNOR2_X1  g666(.A(KEYINPUT61), .B(G155gat), .ZN(new_n868_));
  AND3_X1   g667(.A1(new_n866_), .A2(new_n867_), .A3(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n868_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1346gat));
  OAI21_X1  g670(.A(G162gat), .B1(new_n860_), .B2(new_n555_), .ZN(new_n872_));
  OR2_X1    g671(.A1(new_n606_), .A2(G162gat), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n860_), .B2(new_n873_), .ZN(G1347gat));
  NOR3_X1   g673(.A1(new_n514_), .A2(new_n512_), .A3(new_n371_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n801_), .A2(new_n630_), .A3(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(G169gat), .B1(new_n876_), .B2(new_n596_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(KEYINPUT123), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT123), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n879_), .B(G169gat), .C1(new_n876_), .C2(new_n596_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n878_), .A2(KEYINPUT62), .A3(new_n880_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n876_), .B(KEYINPUT124), .ZN(new_n882_));
  AND2_X1   g681(.A1(new_n597_), .A2(new_n381_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT62), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n877_), .A2(KEYINPUT123), .A3(new_n885_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n881_), .A2(new_n884_), .A3(new_n886_), .ZN(G1348gat));
  NOR2_X1   g686(.A1(new_n316_), .A2(new_n336_), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n801_), .A2(new_n502_), .A3(new_n875_), .A4(new_n888_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(KEYINPUT125), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n882_), .A2(new_n312_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n890_), .B1(new_n891_), .B2(new_n336_), .ZN(G1349gat));
  AND3_X1   g691(.A1(new_n801_), .A2(new_n502_), .A3(new_n875_), .ZN(new_n893_));
  AOI21_X1  g692(.A(G183gat), .B1(new_n893_), .B2(new_n605_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n581_), .A2(new_n378_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n894_), .B1(new_n882_), .B2(new_n895_), .ZN(G1350gat));
  NAND3_X1  g695(.A1(new_n882_), .A2(new_n328_), .A3(new_n550_), .ZN(new_n897_));
  OR2_X1    g696(.A1(new_n876_), .A2(KEYINPUT124), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n876_), .A2(KEYINPUT124), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n555_), .B1(new_n898_), .B2(new_n899_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n897_), .B1(new_n322_), .B2(new_n900_), .ZN(G1351gat));
  NOR2_X1   g700(.A1(new_n514_), .A2(new_n512_), .ZN(new_n902_));
  AND3_X1   g701(.A1(new_n858_), .A2(new_n597_), .A3(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(G197gat), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n903_), .B(new_n904_), .ZN(G1352gat));
  NAND3_X1  g704(.A1(new_n858_), .A2(new_n317_), .A3(new_n902_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n387_), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n906_), .A2(KEYINPUT126), .A3(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT126), .ZN(new_n909_));
  AND3_X1   g708(.A1(new_n858_), .A2(new_n317_), .A3(new_n902_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n909_), .B1(new_n910_), .B2(new_n387_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n906_), .A2(G204gat), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n908_), .B1(new_n911_), .B2(new_n912_), .ZN(G1353gat));
  NAND3_X1  g712(.A1(new_n858_), .A2(new_n605_), .A3(new_n902_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n915_));
  AND2_X1   g714(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n914_), .A2(new_n915_), .A3(new_n916_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n917_), .B1(new_n914_), .B2(new_n915_), .ZN(G1354gat));
  AND2_X1   g717(.A1(new_n858_), .A2(new_n902_), .ZN(new_n919_));
  AOI21_X1  g718(.A(G218gat), .B1(new_n919_), .B2(new_n550_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n556_), .A2(G218gat), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(KEYINPUT127), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n920_), .B1(new_n919_), .B2(new_n922_), .ZN(G1355gat));
endmodule


