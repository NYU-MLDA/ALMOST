//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 1 1 1 0 1 1 0 0 0 1 1 1 1 1 0 1 0 0 1 1 0 1 1 1 0 0 1 1 1 0 1 1 1 0 0 1 1 1 0 0 0 0 0 1 1 1 0 1 1 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n720_, new_n721_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n816_, new_n817_, new_n818_, new_n820_,
    new_n821_, new_n823_, new_n824_, new_n825_, new_n826_, new_n828_,
    new_n830_, new_n831_, new_n833_, new_n834_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n861_, new_n862_, new_n863_, new_n864_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_;
  NOR2_X1   g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203_));
  AOI21_X1  g002(.A(new_n202_), .B1(KEYINPUT1), .B2(new_n203_), .ZN(new_n204_));
  OAI21_X1  g003(.A(new_n204_), .B1(KEYINPUT1), .B2(new_n203_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206_));
  INV_X1    g005(.A(G141gat), .ZN(new_n207_));
  INV_X1    g006(.A(G148gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n205_), .A2(new_n206_), .A3(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT3), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n211_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n206_), .A2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n212_), .A2(new_n214_), .A3(new_n215_), .A4(new_n216_), .ZN(new_n217_));
  XOR2_X1   g016(.A(G155gat), .B(G162gat), .Z(new_n218_));
  AND3_X1   g017(.A1(new_n217_), .A2(KEYINPUT85), .A3(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(KEYINPUT85), .B1(new_n217_), .B2(new_n218_), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n210_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  OR3_X1    g020(.A1(new_n221_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT28), .B1(new_n221_), .B2(KEYINPUT29), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G22gat), .B(G50gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n224_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT90), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n227_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT90), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n229_), .A2(new_n230_), .A3(new_n225_), .ZN(new_n231_));
  INV_X1    g030(.A(G218gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(G211gat), .ZN(new_n233_));
  INV_X1    g032(.A(G211gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(G218gat), .ZN(new_n235_));
  AND2_X1   g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  OR2_X1    g035(.A1(G197gat), .A2(G204gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G197gat), .A2(G204gat), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n237_), .A2(KEYINPUT21), .A3(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT21), .ZN(new_n240_));
  AND2_X1   g039(.A1(G197gat), .A2(G204gat), .ZN(new_n241_));
  NOR2_X1   g040(.A1(G197gat), .A2(G204gat), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n240_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n236_), .A2(new_n239_), .A3(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n240_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT88), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n247_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n237_), .A2(KEYINPUT88), .A3(new_n238_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n246_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT89), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT89), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n246_), .A2(new_n249_), .A3(new_n248_), .A4(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n245_), .B1(new_n251_), .B2(new_n253_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n254_), .A2(KEYINPUT87), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n221_), .A2(KEYINPUT29), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(G106gat), .ZN(new_n258_));
  AND2_X1   g057(.A1(KEYINPUT86), .A2(G233gat), .ZN(new_n259_));
  NOR2_X1   g058(.A1(KEYINPUT86), .A2(G233gat), .ZN(new_n260_));
  OAI21_X1  g059(.A(G228gat), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(G78gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n261_), .B(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(G106gat), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n255_), .A2(new_n265_), .A3(new_n256_), .ZN(new_n266_));
  AND3_X1   g065(.A1(new_n258_), .A2(new_n264_), .A3(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n264_), .B1(new_n258_), .B2(new_n266_), .ZN(new_n268_));
  OAI211_X1 g067(.A(new_n228_), .B(new_n231_), .C1(new_n267_), .C2(new_n268_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n267_), .A2(new_n268_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n230_), .B1(new_n229_), .B2(new_n225_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  XOR2_X1   g071(.A(G127gat), .B(G134gat), .Z(new_n273_));
  XOR2_X1   g072(.A(G113gat), .B(G120gat), .Z(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n221_), .A2(new_n276_), .ZN(new_n277_));
  OAI211_X1 g076(.A(new_n275_), .B(new_n210_), .C1(new_n219_), .C2(new_n220_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G225gat), .A2(G233gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT95), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n280_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT4), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n221_), .A2(new_n285_), .A3(new_n276_), .ZN(new_n286_));
  OAI211_X1 g085(.A(new_n282_), .B(new_n286_), .C1(new_n279_), .C2(new_n285_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G1gat), .B(G29gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT96), .B(G85gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT0), .B(G57gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n284_), .A2(new_n287_), .A3(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n284_), .A2(new_n287_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n292_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n269_), .A2(new_n272_), .A3(new_n293_), .A4(new_n296_), .ZN(new_n297_));
  XOR2_X1   g096(.A(G8gat), .B(G36gat), .Z(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G64gat), .B(G92gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G226gat), .A2(G233gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT19), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT20), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n251_), .A2(new_n253_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(new_n244_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G183gat), .A2(G190gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT23), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT23), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n312_), .A2(G183gat), .A3(G190gat), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT24), .ZN(new_n314_));
  NOR2_X1   g113(.A1(G169gat), .A2(G176gat), .ZN(new_n315_));
  AOI22_X1  g114(.A1(new_n311_), .A2(new_n313_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(G183gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT25), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT25), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(G183gat), .ZN(new_n320_));
  INV_X1    g119(.A(G190gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT26), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT26), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(G190gat), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n318_), .A2(new_n320_), .A3(new_n322_), .A4(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n314_), .B1(G169gat), .B2(G176gat), .ZN(new_n326_));
  INV_X1    g125(.A(new_n315_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n316_), .A2(new_n325_), .A3(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT91), .ZN(new_n330_));
  XNOR2_X1  g129(.A(KEYINPUT25), .B(G183gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT26), .B(G190gat), .ZN(new_n332_));
  AOI22_X1  g131(.A1(new_n331_), .A2(new_n332_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT91), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n333_), .A2(new_n334_), .A3(new_n316_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n310_), .A2(new_n312_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n337_));
  OAI211_X1 g136(.A(new_n336_), .B(new_n337_), .C1(G183gat), .C2(G190gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G169gat), .A2(G176gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT92), .ZN(new_n340_));
  XOR2_X1   g139(.A(KEYINPUT22), .B(G169gat), .Z(new_n341_));
  OAI211_X1 g140(.A(new_n338_), .B(new_n340_), .C1(G176gat), .C2(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n330_), .A2(new_n335_), .A3(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n307_), .B1(new_n309_), .B2(new_n343_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(G169gat), .ZN(new_n346_));
  AOI22_X1  g145(.A1(new_n333_), .A2(new_n316_), .B1(new_n346_), .B2(new_n338_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n308_), .A2(new_n347_), .A3(new_n244_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n306_), .B1(new_n344_), .B2(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n306_), .B1(new_n309_), .B2(new_n343_), .ZN(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT20), .B1(new_n254_), .B2(new_n347_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n303_), .B1(new_n349_), .B2(new_n352_), .ZN(new_n353_));
  AND3_X1   g152(.A1(new_n330_), .A2(new_n335_), .A3(new_n342_), .ZN(new_n354_));
  OAI211_X1 g153(.A(KEYINPUT20), .B(new_n348_), .C1(new_n354_), .C2(new_n254_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(new_n305_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n305_), .B1(new_n354_), .B2(new_n254_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n347_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n307_), .B1(new_n309_), .B2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n357_), .A2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n356_), .A2(new_n302_), .A3(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n353_), .A2(KEYINPUT94), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT27), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n356_), .A2(new_n360_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT94), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n364_), .A2(new_n365_), .A3(new_n303_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n362_), .A2(new_n363_), .A3(new_n366_), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n254_), .A2(new_n329_), .A3(new_n342_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n305_), .B1(new_n368_), .B2(new_n351_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n344_), .A2(new_n306_), .A3(new_n348_), .ZN(new_n370_));
  AND2_X1   g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  OAI211_X1 g170(.A(KEYINPUT27), .B(new_n361_), .C1(new_n371_), .C2(new_n302_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n367_), .A2(new_n372_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n297_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT98), .ZN(new_n375_));
  AND2_X1   g174(.A1(new_n362_), .A2(new_n366_), .ZN(new_n376_));
  XOR2_X1   g175(.A(KEYINPUT97), .B(KEYINPUT33), .Z(new_n377_));
  NAND2_X1  g176(.A1(new_n293_), .A2(new_n377_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n284_), .A2(new_n287_), .A3(KEYINPUT33), .A4(new_n292_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n292_), .B1(new_n280_), .B2(new_n282_), .ZN(new_n380_));
  OAI211_X1 g179(.A(new_n283_), .B(new_n286_), .C1(new_n279_), .C2(new_n285_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n378_), .A2(new_n379_), .A3(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n375_), .B1(new_n376_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n362_), .A2(new_n366_), .ZN(new_n385_));
  AOI22_X1  g184(.A1(new_n293_), .A2(new_n377_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n385_), .A2(KEYINPUT98), .A3(new_n386_), .A4(new_n379_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n302_), .A2(KEYINPUT32), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n371_), .B(new_n389_), .C1(KEYINPUT99), .C2(new_n364_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT99), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n388_), .B1(new_n364_), .B2(new_n391_), .ZN(new_n392_));
  AOI22_X1  g191(.A1(new_n390_), .A2(new_n392_), .B1(new_n296_), .B2(new_n293_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n384_), .A2(new_n387_), .A3(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n269_), .A2(new_n272_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n374_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n347_), .B(KEYINPUT30), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT82), .B(G15gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  XOR2_X1   g199(.A(G71gat), .B(G99gat), .Z(new_n401_));
  XNOR2_X1  g200(.A(KEYINPUT81), .B(G43gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n401_), .B(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G227gat), .A2(G233gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n400_), .B(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n275_), .B(KEYINPUT31), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT83), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT84), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  OR2_X1    g209(.A1(new_n406_), .A2(new_n410_), .ZN(new_n411_));
  OAI211_X1 g210(.A(new_n406_), .B(new_n410_), .C1(KEYINPUT84), .C2(new_n408_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(KEYINPUT100), .B1(new_n397_), .B2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n296_), .A2(new_n293_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n413_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n396_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n418_), .A2(new_n373_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT100), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n385_), .A2(new_n379_), .A3(new_n386_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n393_), .B1(new_n422_), .B2(new_n375_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n418_), .B1(new_n423_), .B2(new_n387_), .ZN(new_n424_));
  OAI211_X1 g223(.A(new_n421_), .B(new_n413_), .C1(new_n424_), .C2(new_n374_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n415_), .A2(new_n420_), .A3(new_n425_), .ZN(new_n426_));
  XOR2_X1   g225(.A(KEYINPUT75), .B(G1gat), .Z(new_n427_));
  INV_X1    g226(.A(G8gat), .ZN(new_n428_));
  OAI21_X1  g227(.A(KEYINPUT14), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G15gat), .B(G22gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G1gat), .B(G8gat), .ZN(new_n432_));
  XOR2_X1   g231(.A(new_n431_), .B(new_n432_), .Z(new_n433_));
  XOR2_X1   g232(.A(G29gat), .B(G36gat), .Z(new_n434_));
  XOR2_X1   g233(.A(G43gat), .B(G50gat), .Z(new_n435_));
  XOR2_X1   g234(.A(new_n434_), .B(new_n435_), .Z(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n433_), .B(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n438_), .A2(G229gat), .A3(G233gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n436_), .B(KEYINPUT15), .ZN(new_n440_));
  OR2_X1    g239(.A1(new_n440_), .A2(new_n433_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n433_), .A2(new_n437_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G229gat), .A2(G233gat), .ZN(new_n443_));
  XOR2_X1   g242(.A(new_n443_), .B(KEYINPUT79), .Z(new_n444_));
  NAND3_X1  g243(.A1(new_n441_), .A2(new_n442_), .A3(new_n444_), .ZN(new_n445_));
  AND2_X1   g244(.A1(new_n439_), .A2(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G113gat), .B(G141gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(KEYINPUT80), .ZN(new_n448_));
  XOR2_X1   g247(.A(G169gat), .B(G197gat), .Z(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n446_), .B(new_n450_), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n426_), .A2(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G57gat), .B(G64gat), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT68), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(KEYINPUT11), .ZN(new_n456_));
  XOR2_X1   g255(.A(G71gat), .B(G78gat), .Z(new_n457_));
  OR2_X1    g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n453_), .B(KEYINPUT68), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT11), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n456_), .A2(new_n461_), .A3(new_n457_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n458_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  XOR2_X1   g263(.A(KEYINPUT10), .B(G99gat), .Z(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(new_n265_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT64), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n466_), .B(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(G99gat), .A2(G106gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n469_), .B(KEYINPUT6), .ZN(new_n470_));
  XOR2_X1   g269(.A(G85gat), .B(G92gat), .Z(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(KEYINPUT9), .ZN(new_n472_));
  INV_X1    g271(.A(G85gat), .ZN(new_n473_));
  INV_X1    g272(.A(G92gat), .ZN(new_n474_));
  OR3_X1    g273(.A1(new_n473_), .A2(new_n474_), .A3(KEYINPUT9), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n468_), .A2(new_n470_), .A3(new_n472_), .A4(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(KEYINPUT66), .B1(G99gat), .B2(G106gat), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NOR3_X1   g277(.A1(KEYINPUT66), .A2(G99gat), .A3(G106gat), .ZN(new_n479_));
  OR3_X1    g278(.A1(new_n478_), .A2(new_n479_), .A3(KEYINPUT7), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT65), .ZN(new_n482_));
  OR2_X1    g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n481_), .A2(new_n482_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n480_), .A2(new_n470_), .A3(new_n483_), .A4(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT8), .ZN(new_n486_));
  OR2_X1    g285(.A1(new_n486_), .A2(KEYINPUT67), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n485_), .A2(new_n471_), .A3(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n486_), .A2(KEYINPUT67), .ZN(new_n490_));
  AOI22_X1  g289(.A1(new_n485_), .A2(new_n471_), .B1(new_n490_), .B2(new_n487_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n476_), .B1(new_n489_), .B2(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n464_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n476_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n491_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT71), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n495_), .A2(new_n496_), .A3(new_n488_), .ZN(new_n497_));
  OAI21_X1  g296(.A(KEYINPUT71), .B1(new_n489_), .B2(new_n491_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n494_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT12), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n463_), .A2(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n493_), .B1(new_n500_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n495_), .A2(new_n488_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n463_), .B1(new_n504_), .B2(new_n476_), .ZN(new_n505_));
  OAI21_X1  g304(.A(KEYINPUT72), .B1(new_n505_), .B2(KEYINPUT12), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n464_), .A2(new_n492_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT72), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n507_), .A2(new_n508_), .A3(new_n501_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n506_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G230gat), .A2(G233gat), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n503_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n493_), .A2(KEYINPUT69), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT70), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n505_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n507_), .A2(KEYINPUT70), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT69), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n517_), .B1(new_n464_), .B2(new_n492_), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n513_), .A2(new_n515_), .A3(new_n516_), .A4(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n511_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n512_), .A2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G120gat), .B(G148gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT5), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G176gat), .B(G204gat), .ZN(new_n525_));
  XOR2_X1   g324(.A(new_n524_), .B(new_n525_), .Z(new_n526_));
  NAND2_X1  g325(.A1(new_n522_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n526_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n512_), .A2(new_n521_), .A3(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT13), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n527_), .A2(KEYINPUT13), .A3(new_n529_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G231gat), .A2(G233gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT76), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n433_), .B(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(new_n464_), .ZN(new_n539_));
  XOR2_X1   g338(.A(G183gat), .B(G211gat), .Z(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT78), .ZN(new_n541_));
  XOR2_X1   g340(.A(G127gat), .B(G155gat), .Z(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  XOR2_X1   g342(.A(KEYINPUT77), .B(KEYINPUT16), .Z(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT17), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n539_), .A2(new_n547_), .ZN(new_n548_));
  AND2_X1   g347(.A1(new_n545_), .A2(new_n546_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n539_), .B1(new_n547_), .B2(new_n549_), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT37), .ZN(new_n553_));
  XOR2_X1   g352(.A(G134gat), .B(G162gat), .Z(new_n554_));
  XNOR2_X1  g353(.A(G190gat), .B(G218gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT36), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n556_), .A2(new_n557_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(G232gat), .A2(G233gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT34), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT35), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n440_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n500_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT73), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n568_), .B1(new_n499_), .B2(new_n440_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n563_), .A2(new_n564_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n504_), .A2(new_n437_), .A3(new_n476_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n570_), .A2(new_n571_), .A3(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n565_), .B1(new_n569_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT74), .ZN(new_n575_));
  INV_X1    g374(.A(new_n565_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n572_), .A2(new_n576_), .A3(new_n571_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n575_), .B1(new_n567_), .B2(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n499_), .A2(new_n440_), .ZN(new_n580_));
  NOR3_X1   g379(.A1(new_n580_), .A2(new_n577_), .A3(KEYINPUT74), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  AOI211_X1 g381(.A(new_n559_), .B(new_n560_), .C1(new_n574_), .C2(new_n582_), .ZN(new_n583_));
  AND4_X1   g382(.A1(new_n557_), .A2(new_n574_), .A3(new_n582_), .A4(new_n556_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n553_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n560_), .B1(new_n574_), .B2(new_n582_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(new_n558_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n574_), .A2(new_n582_), .A3(new_n557_), .A4(new_n556_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n587_), .A2(KEYINPUT37), .A3(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n585_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n452_), .A2(new_n535_), .A3(new_n552_), .A4(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT101), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n594_), .A2(new_n416_), .A3(new_n427_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT38), .ZN(new_n596_));
  OR2_X1    g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT102), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n598_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n587_), .A2(KEYINPUT102), .A3(new_n588_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  AND2_X1   g400(.A1(new_n426_), .A2(new_n601_), .ZN(new_n602_));
  AND4_X1   g401(.A1(new_n451_), .A2(new_n602_), .A3(new_n535_), .A4(new_n552_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(new_n416_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(G1gat), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n595_), .A2(new_n596_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n597_), .A2(new_n605_), .A3(new_n606_), .ZN(G1324gat));
  NAND3_X1  g406(.A1(new_n594_), .A2(new_n428_), .A3(new_n373_), .ZN(new_n608_));
  AOI211_X1 g407(.A(KEYINPUT39), .B(new_n428_), .C1(new_n603_), .C2(new_n373_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT39), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n603_), .A2(new_n373_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n610_), .B1(new_n611_), .B2(G8gat), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n608_), .B1(new_n609_), .B2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT40), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  OAI211_X1 g414(.A(new_n608_), .B(KEYINPUT40), .C1(new_n612_), .C2(new_n609_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(G1325gat));
  INV_X1    g416(.A(G15gat), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n618_), .B1(new_n603_), .B2(new_n414_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT41), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n594_), .A2(new_n618_), .A3(new_n414_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(G1326gat));
  INV_X1    g421(.A(KEYINPUT42), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n603_), .A2(new_n418_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(G22gat), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT103), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n625_), .A2(KEYINPUT103), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n623_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n628_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n630_), .A2(KEYINPUT42), .A3(new_n626_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n396_), .A2(G22gat), .ZN(new_n632_));
  XOR2_X1   g431(.A(new_n632_), .B(KEYINPUT104), .Z(new_n633_));
  NAND2_X1  g432(.A1(new_n594_), .A2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n629_), .A2(new_n631_), .A3(new_n634_), .ZN(G1327gat));
  NOR3_X1   g434(.A1(new_n601_), .A2(new_n534_), .A3(new_n552_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n452_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(G29gat), .B1(new_n638_), .B2(new_n416_), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n532_), .A2(new_n451_), .A3(new_n533_), .A4(new_n551_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT105), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT43), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n426_), .A2(new_n642_), .A3(new_n590_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(KEYINPUT106), .B(KEYINPUT43), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n645_), .B1(new_n426_), .B2(new_n590_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n641_), .B1(new_n643_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT44), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  OAI211_X1 g448(.A(KEYINPUT44), .B(new_n641_), .C1(new_n643_), .C2(new_n646_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n416_), .A2(G29gat), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n639_), .B1(new_n651_), .B2(new_n652_), .ZN(G1328gat));
  INV_X1    g452(.A(new_n373_), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n637_), .A2(G36gat), .A3(new_n654_), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n655_), .B(KEYINPUT45), .Z(new_n656_));
  NAND3_X1  g455(.A1(new_n649_), .A2(new_n373_), .A3(new_n650_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(G36gat), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT46), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n656_), .A2(KEYINPUT46), .A3(new_n658_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1329gat));
  XNOR2_X1  g462(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(G43gat), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n413_), .A2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n649_), .A2(new_n650_), .A3(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT108), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n666_), .B1(new_n637_), .B2(new_n413_), .ZN(new_n670_));
  AND3_X1   g469(.A1(new_n668_), .A2(new_n669_), .A3(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n669_), .B1(new_n668_), .B2(new_n670_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n665_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n668_), .A2(new_n670_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(KEYINPUT108), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n668_), .A2(new_n669_), .A3(new_n670_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n675_), .A2(new_n676_), .A3(new_n664_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n673_), .A2(new_n677_), .ZN(G1330gat));
  OR3_X1    g477(.A1(new_n637_), .A2(G50gat), .A3(new_n396_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n651_), .A2(new_n418_), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n680_), .A2(KEYINPUT109), .A3(G50gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(KEYINPUT109), .B1(new_n680_), .B2(G50gat), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n679_), .B1(new_n681_), .B2(new_n682_), .ZN(G1331gat));
  INV_X1    g482(.A(new_n451_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n426_), .A2(new_n684_), .ZN(new_n685_));
  AND4_X1   g484(.A1(new_n534_), .A2(new_n685_), .A3(new_n552_), .A4(new_n591_), .ZN(new_n686_));
  INV_X1    g485(.A(G57gat), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n686_), .A2(new_n687_), .A3(new_n416_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n551_), .A2(new_n451_), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n602_), .A2(new_n534_), .A3(new_n689_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n690_), .A2(new_n416_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n688_), .B1(new_n691_), .B2(new_n687_), .ZN(G1332gat));
  INV_X1    g491(.A(G64gat), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n693_), .B1(new_n690_), .B2(new_n373_), .ZN(new_n694_));
  XOR2_X1   g493(.A(new_n694_), .B(KEYINPUT48), .Z(new_n695_));
  NAND3_X1  g494(.A1(new_n686_), .A2(new_n693_), .A3(new_n373_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(G1333gat));
  INV_X1    g496(.A(G71gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n698_), .B1(new_n690_), .B2(new_n414_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT49), .Z(new_n700_));
  NAND3_X1  g499(.A1(new_n686_), .A2(new_n698_), .A3(new_n414_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(G1334gat));
  NAND3_X1  g501(.A1(new_n686_), .A2(new_n262_), .A3(new_n418_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n690_), .A2(new_n418_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n704_), .A2(G78gat), .A3(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n705_), .B1(new_n704_), .B2(G78gat), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n703_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT111), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n708_), .B(new_n709_), .ZN(G1335gat));
  NOR2_X1   g509(.A1(new_n601_), .A2(new_n552_), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n685_), .A2(new_n534_), .A3(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(G85gat), .B1(new_n712_), .B2(new_n416_), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n713_), .B(KEYINPUT112), .Z(new_n714_));
  OR2_X1    g513(.A1(new_n643_), .A2(new_n646_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n535_), .A2(new_n451_), .A3(new_n552_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n473_), .B1(new_n296_), .B2(new_n293_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n714_), .B1(new_n717_), .B2(new_n718_), .ZN(G1336gat));
  NAND3_X1  g518(.A1(new_n712_), .A2(new_n474_), .A3(new_n373_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n717_), .A2(new_n373_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n720_), .B1(new_n721_), .B2(new_n474_), .ZN(G1337gat));
  NAND3_X1  g521(.A1(new_n715_), .A2(new_n414_), .A3(new_n716_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n414_), .A2(new_n465_), .ZN(new_n724_));
  AOI22_X1  g523(.A1(new_n723_), .A2(G99gat), .B1(new_n712_), .B2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT114), .ZN(new_n726_));
  XNOR2_X1  g525(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n725_), .A2(new_n726_), .A3(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT51), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n725_), .A2(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n726_), .B1(new_n725_), .B2(new_n727_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n728_), .B1(new_n730_), .B2(new_n731_), .ZN(G1338gat));
  NAND3_X1  g531(.A1(new_n712_), .A2(new_n265_), .A3(new_n418_), .ZN(new_n733_));
  OAI211_X1 g532(.A(new_n418_), .B(new_n716_), .C1(new_n643_), .C2(new_n646_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT52), .ZN(new_n735_));
  AND3_X1   g534(.A1(new_n734_), .A2(new_n735_), .A3(G106gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n734_), .B2(G106gat), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n733_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g538(.A(new_n444_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n441_), .A2(new_n442_), .A3(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n450_), .B1(new_n438_), .B2(new_n444_), .ZN(new_n742_));
  AOI22_X1  g541(.A1(new_n446_), .A2(new_n450_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n529_), .A2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT55), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n746_), .B1(new_n520_), .B2(KEYINPUT116), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n747_), .B1(new_n746_), .B2(new_n520_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n503_), .A2(new_n510_), .A3(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n502_), .ZN(new_n750_));
  OAI22_X1  g549(.A1(new_n499_), .A2(new_n750_), .B1(new_n464_), .B2(new_n492_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(new_n506_), .B2(new_n509_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n747_), .ZN(new_n753_));
  OAI211_X1 g552(.A(new_n749_), .B(new_n526_), .C1(new_n752_), .C2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT56), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n503_), .A2(new_n510_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n528_), .B1(new_n757_), .B2(new_n747_), .ZN(new_n758_));
  AOI21_X1  g557(.A(KEYINPUT56), .B1(new_n758_), .B2(new_n749_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n745_), .B1(new_n756_), .B2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT117), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT58), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n760_), .A2(new_n761_), .A3(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n754_), .A2(new_n755_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n758_), .A2(KEYINPUT56), .A3(new_n749_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n744_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  OAI21_X1  g565(.A(KEYINPUT58), .B1(new_n766_), .B2(KEYINPUT117), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n590_), .A2(new_n763_), .A3(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT118), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n590_), .A2(new_n763_), .A3(new_n767_), .A4(KEYINPUT118), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT57), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n599_), .A2(new_n600_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n764_), .A2(new_n765_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n451_), .A2(new_n529_), .ZN(new_n775_));
  AOI22_X1  g574(.A1(new_n774_), .A2(new_n775_), .B1(new_n530_), .B2(new_n743_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n772_), .B1(new_n773_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n776_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n601_), .A2(KEYINPUT57), .A3(new_n778_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n770_), .A2(new_n771_), .A3(new_n777_), .A4(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n532_), .A2(new_n533_), .A3(new_n689_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT115), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n532_), .A2(KEYINPUT115), .A3(new_n689_), .A4(new_n533_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n591_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT54), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT54), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n785_), .A2(new_n788_), .A3(new_n591_), .ZN(new_n789_));
  AOI22_X1  g588(.A1(new_n780_), .A2(new_n551_), .B1(new_n787_), .B2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n419_), .A2(new_n414_), .A3(new_n416_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(G113gat), .B1(new_n792_), .B2(new_n451_), .ZN(new_n793_));
  OAI21_X1  g592(.A(KEYINPUT59), .B1(new_n790_), .B2(new_n791_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT119), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n787_), .A2(new_n789_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n779_), .A2(new_n777_), .A3(new_n768_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n551_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n798_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n791_), .A2(KEYINPUT59), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n794_), .A2(new_n795_), .A3(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n795_), .B1(new_n794_), .B2(new_n801_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT120), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n451_), .A2(new_n805_), .A3(G113gat), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n806_), .B1(new_n805_), .B2(G113gat), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n793_), .B1(new_n804_), .B2(new_n807_), .ZN(G1340gat));
  NOR2_X1   g607(.A1(new_n535_), .A2(KEYINPUT60), .ZN(new_n809_));
  MUX2_X1   g608(.A(new_n809_), .B(KEYINPUT60), .S(G120gat), .Z(new_n810_));
  NAND2_X1  g609(.A1(new_n792_), .A2(new_n810_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n811_), .B(KEYINPUT121), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n794_), .A2(new_n534_), .A3(new_n801_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(G120gat), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(new_n814_), .ZN(G1341gat));
  AOI21_X1  g614(.A(G127gat), .B1(new_n792_), .B2(new_n552_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n552_), .A2(G127gat), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(KEYINPUT122), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n816_), .B1(new_n804_), .B2(new_n818_), .ZN(G1342gat));
  AOI21_X1  g618(.A(G134gat), .B1(new_n792_), .B2(new_n773_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n590_), .A2(G134gat), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n820_), .B1(new_n804_), .B2(new_n821_), .ZN(G1343gat));
  NAND4_X1  g621(.A1(new_n413_), .A2(new_n654_), .A3(new_n416_), .A4(new_n418_), .ZN(new_n823_));
  OR2_X1    g622(.A1(new_n790_), .A2(new_n823_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n824_), .A2(new_n684_), .ZN(new_n825_));
  XOR2_X1   g624(.A(KEYINPUT123), .B(G141gat), .Z(new_n826_));
  XNOR2_X1  g625(.A(new_n825_), .B(new_n826_), .ZN(G1344gat));
  NOR2_X1   g626(.A1(new_n824_), .A2(new_n535_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n828_), .B(new_n208_), .ZN(G1345gat));
  NOR2_X1   g628(.A1(new_n824_), .A2(new_n551_), .ZN(new_n830_));
  XOR2_X1   g629(.A(KEYINPUT61), .B(G155gat), .Z(new_n831_));
  XNOR2_X1  g630(.A(new_n830_), .B(new_n831_), .ZN(G1346gat));
  OAI21_X1  g631(.A(G162gat), .B1(new_n824_), .B2(new_n591_), .ZN(new_n833_));
  OR2_X1    g632(.A1(new_n601_), .A2(G162gat), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n833_), .B1(new_n824_), .B2(new_n834_), .ZN(G1347gat));
  NAND2_X1  g634(.A1(new_n417_), .A2(new_n373_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n836_), .A2(new_n418_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n799_), .A2(new_n451_), .A3(new_n837_), .ZN(new_n838_));
  XOR2_X1   g637(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n838_), .A2(G169gat), .A3(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n837_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n842_), .B1(new_n796_), .B2(new_n798_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n341_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n843_), .A2(new_n844_), .A3(new_n451_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n841_), .A2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n840_), .B1(new_n838_), .B2(G169gat), .ZN(new_n847_));
  OAI21_X1  g646(.A(KEYINPUT125), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n847_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT125), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n849_), .A2(new_n850_), .A3(new_n845_), .A4(new_n841_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n848_), .A2(new_n851_), .ZN(G1348gat));
  AOI21_X1  g651(.A(G176gat), .B1(new_n843_), .B2(new_n534_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n790_), .A2(new_n418_), .ZN(new_n854_));
  INV_X1    g653(.A(G176gat), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n535_), .A2(new_n855_), .A3(new_n836_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n853_), .B1(new_n854_), .B2(new_n856_), .ZN(G1349gat));
  NAND4_X1  g656(.A1(new_n854_), .A2(new_n373_), .A3(new_n417_), .A4(new_n552_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n551_), .A2(new_n331_), .ZN(new_n859_));
  AOI22_X1  g658(.A1(new_n858_), .A2(new_n317_), .B1(new_n843_), .B2(new_n859_), .ZN(G1350gat));
  NAND3_X1  g659(.A1(new_n843_), .A2(new_n332_), .A3(new_n773_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n843_), .A2(new_n590_), .ZN(new_n862_));
  AND3_X1   g661(.A1(new_n862_), .A2(KEYINPUT126), .A3(G190gat), .ZN(new_n863_));
  AOI21_X1  g662(.A(KEYINPUT126), .B1(new_n862_), .B2(G190gat), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n861_), .B1(new_n863_), .B2(new_n864_), .ZN(G1351gat));
  NOR4_X1   g664(.A1(new_n790_), .A2(new_n414_), .A3(new_n654_), .A4(new_n297_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n451_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n534_), .ZN(new_n869_));
  XOR2_X1   g668(.A(KEYINPUT127), .B(G204gat), .Z(new_n870_));
  XNOR2_X1  g669(.A(new_n869_), .B(new_n870_), .ZN(G1353gat));
  NAND2_X1  g670(.A1(new_n866_), .A2(new_n552_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(KEYINPUT63), .B(G211gat), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n874_), .B1(new_n872_), .B2(new_n875_), .ZN(G1354gat));
  NAND3_X1  g675(.A1(new_n866_), .A2(new_n232_), .A3(new_n773_), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n866_), .A2(new_n590_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n878_), .B2(new_n232_), .ZN(G1355gat));
endmodule


