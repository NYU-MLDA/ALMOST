//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 1 1 0 0 0 1 0 1 0 0 0 1 1 1 1 0 0 1 0 1 0 1 1 1 1 1 1 0 0 0 1 1 1 1 0 0 1 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n698_, new_n699_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n871_, new_n872_, new_n874_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n914_, new_n915_, new_n916_, new_n918_, new_n920_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n927_, new_n928_,
    new_n929_, new_n930_;
  INV_X1    g000(.A(KEYINPUT3), .ZN(new_n202_));
  INV_X1    g001(.A(G141gat), .ZN(new_n203_));
  INV_X1    g002(.A(G148gat), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n202_), .A2(new_n203_), .A3(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT2), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n205_), .A2(new_n208_), .A3(new_n209_), .A4(new_n210_), .ZN(new_n211_));
  OR2_X1    g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213_));
  AND2_X1   g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n211_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT81), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(G127gat), .ZN(new_n218_));
  INV_X1    g017(.A(G134gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G127gat), .A2(G134gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(G113gat), .ZN(new_n223_));
  INV_X1    g022(.A(G120gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G113gat), .A2(G120gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n222_), .A2(new_n227_), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n220_), .A2(new_n225_), .A3(new_n221_), .A4(new_n226_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  AND2_X1   g029(.A1(G155gat), .A2(G162gat), .ZN(new_n231_));
  AOI22_X1  g030(.A1(new_n231_), .A2(KEYINPUT1), .B1(new_n203_), .B2(new_n204_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT1), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n212_), .A2(new_n233_), .A3(new_n213_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n232_), .A2(new_n234_), .A3(new_n206_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n211_), .A2(KEYINPUT81), .A3(new_n214_), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n217_), .A2(new_n230_), .A3(new_n235_), .A4(new_n236_), .ZN(new_n237_));
  AND3_X1   g036(.A1(new_n211_), .A2(KEYINPUT81), .A3(new_n214_), .ZN(new_n238_));
  AOI21_X1  g037(.A(KEYINPUT81), .B1(new_n211_), .B2(new_n214_), .ZN(new_n239_));
  AND3_X1   g038(.A1(new_n232_), .A2(new_n234_), .A3(new_n206_), .ZN(new_n240_));
  NOR3_X1   g039(.A1(new_n238_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT79), .ZN(new_n242_));
  OR3_X1    g041(.A1(new_n222_), .A2(new_n227_), .A3(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n228_), .A2(new_n242_), .A3(new_n229_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  OAI211_X1 g045(.A(KEYINPUT4), .B(new_n237_), .C1(new_n241_), .C2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G225gat), .A2(G233gat), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n217_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT90), .B(KEYINPUT4), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n250_), .A2(new_n245_), .A3(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n247_), .A2(new_n249_), .A3(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT91), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n250_), .A2(new_n245_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n256_), .A2(new_n237_), .A3(new_n248_), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n247_), .A2(KEYINPUT91), .A3(new_n249_), .A4(new_n252_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n255_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G57gat), .B(G85gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT92), .B(KEYINPUT0), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G1gat), .B(G29gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(KEYINPUT96), .B1(new_n259_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n264_), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n255_), .A2(new_n257_), .A3(new_n258_), .A4(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n259_), .A2(KEYINPUT96), .A3(new_n264_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n266_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT80), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT31), .ZN(new_n272_));
  OR2_X1    g071(.A1(KEYINPUT76), .A2(G176gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(KEYINPUT76), .A2(G176gat), .ZN(new_n274_));
  OR2_X1    g073(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n276_));
  AOI22_X1  g075(.A1(new_n273_), .A2(new_n274_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G169gat), .A2(G176gat), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT77), .B1(new_n277_), .B2(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n283_));
  INV_X1    g082(.A(G183gat), .ZN(new_n284_));
  INV_X1    g083(.A(G190gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n282_), .A2(new_n283_), .A3(new_n286_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(KEYINPUT76), .A2(G176gat), .ZN(new_n288_));
  AND2_X1   g087(.A1(KEYINPUT76), .A2(G176gat), .ZN(new_n289_));
  AND2_X1   g088(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n290_));
  NOR2_X1   g089(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n291_));
  OAI22_X1  g090(.A1(new_n288_), .A2(new_n289_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT77), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n292_), .A2(new_n293_), .A3(new_n278_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n280_), .A2(new_n287_), .A3(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT30), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT75), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n297_), .B1(new_n285_), .B2(KEYINPUT26), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT25), .B(G183gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT26), .B(G190gat), .ZN(new_n300_));
  OAI211_X1 g099(.A(new_n298_), .B(new_n299_), .C1(new_n300_), .C2(new_n297_), .ZN(new_n301_));
  OR2_X1    g100(.A1(G169gat), .A2(G176gat), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n302_), .A2(KEYINPUT24), .A3(new_n278_), .ZN(new_n303_));
  NOR3_X1   g102(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n304_));
  AND3_X1   g103(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n305_));
  NOR3_X1   g104(.A1(new_n304_), .A2(new_n305_), .A3(new_n281_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n301_), .A2(new_n303_), .A3(new_n306_), .ZN(new_n307_));
  AND3_X1   g106(.A1(new_n295_), .A2(new_n296_), .A3(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n296_), .B1(new_n295_), .B2(new_n307_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n272_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n273_), .A2(new_n274_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT22), .B(G169gat), .ZN(new_n312_));
  AOI211_X1 g111(.A(KEYINPUT77), .B(new_n279_), .C1(new_n311_), .C2(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n293_), .B1(new_n292_), .B2(new_n278_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n287_), .ZN(new_n315_));
  NOR3_X1   g114(.A1(new_n313_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n307_), .ZN(new_n317_));
  OAI21_X1  g116(.A(KEYINPUT30), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n295_), .A2(new_n296_), .A3(new_n307_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n318_), .A2(KEYINPUT31), .A3(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G15gat), .B(G43gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n245_), .B(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  AND3_X1   g122(.A1(new_n310_), .A2(new_n320_), .A3(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n323_), .B1(new_n310_), .B2(new_n320_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G227gat), .A2(G233gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT78), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G71gat), .B(G99gat), .ZN(new_n328_));
  XOR2_X1   g127(.A(new_n327_), .B(new_n328_), .Z(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NOR3_X1   g129(.A1(new_n324_), .A2(new_n325_), .A3(new_n330_), .ZN(new_n331_));
  NOR3_X1   g130(.A1(new_n308_), .A2(new_n309_), .A3(new_n272_), .ZN(new_n332_));
  AOI21_X1  g131(.A(KEYINPUT31), .B1(new_n318_), .B2(new_n319_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n322_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n310_), .A2(new_n320_), .A3(new_n323_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n329_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n271_), .B1(new_n331_), .B2(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n330_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n334_), .A2(new_n329_), .A3(new_n335_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n338_), .A2(KEYINPUT80), .A3(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n250_), .A2(KEYINPUT29), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT21), .ZN(new_n342_));
  INV_X1    g141(.A(G204gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(G197gat), .ZN(new_n344_));
  INV_X1    g143(.A(G197gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(G204gat), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n342_), .B1(new_n344_), .B2(new_n346_), .ZN(new_n347_));
  AND2_X1   g146(.A1(G211gat), .A2(G218gat), .ZN(new_n348_));
  NOR2_X1   g147(.A1(G211gat), .A2(G218gat), .ZN(new_n349_));
  OAI21_X1  g148(.A(KEYINPUT83), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  OR2_X1    g149(.A1(G211gat), .A2(G218gat), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT83), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G211gat), .A2(G218gat), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n351_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n347_), .A2(new_n350_), .A3(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT84), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT84), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n347_), .A2(new_n354_), .A3(new_n350_), .A4(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  AND3_X1   g158(.A1(new_n344_), .A2(new_n346_), .A3(new_n342_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n348_), .A2(new_n349_), .ZN(new_n361_));
  NOR3_X1   g160(.A1(new_n360_), .A2(new_n347_), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n359_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(G228gat), .ZN(new_n365_));
  INV_X1    g164(.A(G233gat), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  AND3_X1   g167(.A1(new_n341_), .A2(new_n364_), .A3(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n368_), .B1(new_n341_), .B2(new_n364_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G78gat), .B(G106gat), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NOR3_X1   g171(.A1(new_n369_), .A2(new_n370_), .A3(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT29), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n238_), .A2(new_n239_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n374_), .B1(new_n375_), .B2(new_n235_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n362_), .B1(new_n356_), .B2(new_n358_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n367_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n341_), .A2(new_n364_), .A3(new_n368_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n371_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT85), .B1(new_n373_), .B2(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n372_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT85), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n378_), .A2(new_n379_), .A3(new_n371_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n382_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n241_), .A2(new_n374_), .ZN(new_n386_));
  XOR2_X1   g185(.A(G22gat), .B(G50gat), .Z(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT82), .B(KEYINPUT28), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n386_), .B(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n381_), .A2(new_n385_), .A3(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n390_), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n392_), .A2(new_n382_), .A3(new_n383_), .A4(new_n384_), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n337_), .A2(new_n340_), .A3(new_n391_), .A4(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n391_), .A2(new_n393_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n338_), .A2(new_n339_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n270_), .B1(new_n394_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT27), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G226gat), .A2(G233gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT19), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT20), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT87), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n278_), .A2(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n278_), .A2(new_n404_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n287_), .A2(new_n292_), .A3(new_n405_), .A4(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT88), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  AOI22_X1  g209(.A1(new_n311_), .A2(new_n312_), .B1(new_n404_), .B2(new_n278_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n411_), .A2(KEYINPUT88), .A3(new_n287_), .A4(new_n407_), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n282_), .B(new_n283_), .C1(new_n302_), .C2(KEYINPUT24), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n278_), .A2(KEYINPUT86), .A3(KEYINPUT24), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(KEYINPUT86), .B1(new_n278_), .B2(KEYINPUT24), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n413_), .B1(new_n417_), .B2(new_n302_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n299_), .A2(new_n300_), .ZN(new_n419_));
  AOI22_X1  g218(.A1(new_n410_), .A2(new_n412_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n403_), .B1(new_n420_), .B2(new_n377_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n295_), .A2(new_n307_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT89), .ZN(new_n423_));
  AND3_X1   g222(.A1(new_n422_), .A2(new_n364_), .A3(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n423_), .B1(new_n422_), .B2(new_n364_), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n402_), .B(new_n421_), .C1(new_n424_), .C2(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G8gat), .B(G36gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(G92gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(KEYINPUT18), .B(G64gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n428_), .B(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT20), .B1(new_n420_), .B2(new_n377_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n422_), .A2(new_n364_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n401_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  AND3_X1   g233(.A1(new_n426_), .A2(new_n431_), .A3(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n431_), .B1(new_n426_), .B2(new_n434_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n399_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT97), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  OAI211_X1 g238(.A(KEYINPUT97), .B(new_n399_), .C1(new_n435_), .C2(new_n436_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT95), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n305_), .A2(new_n281_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n406_), .B1(new_n442_), .B2(new_n286_), .ZN(new_n443_));
  AOI22_X1  g242(.A1(new_n418_), .A2(new_n419_), .B1(new_n411_), .B2(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n403_), .B1(new_n444_), .B2(new_n377_), .ZN(new_n445_));
  OAI22_X1  g244(.A1(new_n424_), .A2(new_n425_), .B1(new_n441_), .B2(new_n445_), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n445_), .A2(new_n441_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n401_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  OR3_X1    g247(.A1(new_n432_), .A2(new_n433_), .A3(new_n401_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n435_), .B1(new_n450_), .B2(new_n430_), .ZN(new_n451_));
  AOI22_X1  g250(.A1(new_n439_), .A2(new_n440_), .B1(new_n451_), .B2(KEYINPUT27), .ZN(new_n452_));
  INV_X1    g251(.A(new_n268_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT33), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n435_), .A2(new_n436_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n247_), .A2(new_n248_), .A3(new_n252_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n256_), .A2(new_n237_), .A3(new_n249_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n456_), .A2(new_n264_), .A3(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(KEYINPUT93), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT33), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n268_), .A2(new_n460_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n454_), .A2(new_n455_), .A3(new_n459_), .A4(new_n461_), .ZN(new_n462_));
  AND3_X1   g261(.A1(new_n259_), .A2(KEYINPUT96), .A3(new_n264_), .ZN(new_n463_));
  NOR3_X1   g262(.A1(new_n463_), .A2(new_n265_), .A3(new_n453_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT94), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n426_), .A2(new_n465_), .A3(new_n434_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n448_), .A2(new_n466_), .A3(new_n449_), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n431_), .A2(KEYINPUT32), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n468_), .A2(new_n465_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n470_), .A2(new_n426_), .A3(new_n434_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n462_), .B1(new_n464_), .B2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n395_), .A2(new_n340_), .A3(new_n337_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  AOI22_X1  g274(.A1(new_n398_), .A2(new_n452_), .B1(new_n473_), .B2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G15gat), .B(G22gat), .ZN(new_n477_));
  INV_X1    g276(.A(G1gat), .ZN(new_n478_));
  INV_X1    g277(.A(G8gat), .ZN(new_n479_));
  OAI21_X1  g278(.A(KEYINPUT14), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G1gat), .B(G8gat), .ZN(new_n482_));
  OR2_X1    g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n481_), .A2(new_n482_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G231gat), .A2(G233gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT69), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n485_), .B(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G57gat), .B(G64gat), .ZN(new_n489_));
  OR2_X1    g288(.A1(new_n489_), .A2(KEYINPUT11), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(KEYINPUT11), .ZN(new_n491_));
  XOR2_X1   g290(.A(G71gat), .B(G78gat), .Z(new_n492_));
  NAND3_X1  g291(.A1(new_n490_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n493_));
  OR2_X1    g292(.A1(new_n491_), .A2(new_n492_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n488_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n488_), .A2(new_n496_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  XOR2_X1   g299(.A(KEYINPUT71), .B(KEYINPUT16), .Z(new_n501_));
  XNOR2_X1  g300(.A(G183gat), .B(G211gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  XOR2_X1   g302(.A(G127gat), .B(G155gat), .Z(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT17), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n500_), .A2(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(KEYINPUT70), .B1(new_n498_), .B2(new_n499_), .ZN(new_n508_));
  AND2_X1   g307(.A1(new_n505_), .A2(KEYINPUT17), .ZN(new_n509_));
  OR2_X1    g308(.A1(new_n488_), .A2(new_n496_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT70), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n510_), .A2(new_n511_), .A3(new_n497_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n508_), .A2(new_n509_), .A3(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT72), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n508_), .A2(new_n512_), .A3(KEYINPUT72), .A4(new_n509_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n507_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT73), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  AOI211_X1 g318(.A(KEYINPUT73), .B(new_n507_), .C1(new_n515_), .C2(new_n516_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n476_), .A2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT68), .B(KEYINPUT37), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  XOR2_X1   g323(.A(G85gat), .B(G92gat), .Z(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(KEYINPUT9), .ZN(new_n526_));
  XOR2_X1   g325(.A(KEYINPUT10), .B(G99gat), .Z(new_n527_));
  INV_X1    g326(.A(G106gat), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G99gat), .A2(G106gat), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT6), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n533_));
  AND2_X1   g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT9), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n535_), .A2(G85gat), .A3(G92gat), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n526_), .A2(new_n529_), .A3(new_n534_), .A4(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT7), .ZN(new_n538_));
  INV_X1    g337(.A(G99gat), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n538_), .A2(new_n539_), .A3(new_n528_), .A4(KEYINPUT64), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT64), .ZN(new_n541_));
  OAI22_X1  g340(.A1(new_n541_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n541_), .A2(KEYINPUT7), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n532_), .A2(new_n533_), .A3(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n525_), .B1(new_n543_), .B2(new_n545_), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n546_), .A2(KEYINPUT8), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT8), .ZN(new_n548_));
  OAI211_X1 g347(.A(new_n548_), .B(new_n525_), .C1(new_n543_), .C2(new_n545_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n537_), .B1(new_n547_), .B2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G29gat), .B(G36gat), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G43gat), .B(G50gat), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n554_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(new_n552_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT15), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n555_), .A2(new_n557_), .A3(KEYINPUT15), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n551_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G232gat), .A2(G233gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT34), .ZN(new_n565_));
  XNOR2_X1  g364(.A(KEYINPUT66), .B(KEYINPUT67), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  OAI221_X1 g366(.A(new_n563_), .B1(KEYINPUT35), .B2(new_n567_), .C1(new_n558_), .C2(new_n551_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(KEYINPUT35), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G190gat), .B(G218gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G134gat), .B(G162gat), .ZN(new_n572_));
  XOR2_X1   g371(.A(new_n571_), .B(new_n572_), .Z(new_n573_));
  INV_X1    g372(.A(KEYINPUT36), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n570_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n573_), .B(KEYINPUT36), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n570_), .A2(new_n578_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n524_), .B1(new_n577_), .B2(new_n579_), .ZN(new_n580_));
  OAI211_X1 g379(.A(new_n576_), .B(new_n523_), .C1(new_n578_), .C2(new_n570_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n522_), .A2(new_n582_), .ZN(new_n583_));
  AOI22_X1  g382(.A1(new_n560_), .A2(new_n561_), .B1(new_n484_), .B2(new_n483_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n485_), .A2(new_n558_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G229gat), .A2(G233gat), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NOR3_X1   g386(.A1(new_n584_), .A2(new_n585_), .A3(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n485_), .B(new_n558_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n588_), .B1(new_n587_), .B2(new_n589_), .ZN(new_n590_));
  XOR2_X1   g389(.A(G169gat), .B(G197gat), .Z(new_n591_));
  XNOR2_X1  g390(.A(G113gat), .B(G141gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n593_), .A2(KEYINPUT74), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n590_), .B(new_n594_), .Z(new_n595_));
  NAND2_X1  g394(.A1(G230gat), .A2(G233gat), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n551_), .A2(new_n496_), .ZN(new_n598_));
  OAI211_X1 g397(.A(new_n495_), .B(new_n537_), .C1(new_n547_), .C2(new_n550_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n598_), .A2(KEYINPUT12), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT12), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n551_), .A2(new_n601_), .A3(new_n496_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n597_), .B1(new_n600_), .B2(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n596_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(KEYINPUT65), .B(KEYINPUT5), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G176gat), .B(G204gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G120gat), .B(G148gat), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n608_), .B(new_n609_), .Z(new_n610_));
  XNOR2_X1  g409(.A(new_n605_), .B(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT13), .ZN(new_n612_));
  NOR3_X1   g411(.A1(new_n583_), .A2(new_n595_), .A3(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n613_), .A2(new_n478_), .A3(new_n270_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT38), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n394_), .A2(new_n397_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n616_), .A2(new_n464_), .A3(new_n452_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n473_), .A2(new_n475_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n577_), .A2(new_n579_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT98), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n612_), .A2(new_n595_), .ZN(new_n623_));
  AND3_X1   g422(.A1(new_n622_), .A2(new_n517_), .A3(new_n623_), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n624_), .A2(new_n270_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n615_), .B1(new_n478_), .B2(new_n625_), .ZN(G1324gat));
  INV_X1    g425(.A(new_n452_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n613_), .A2(new_n479_), .A3(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT39), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n624_), .A2(new_n627_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n629_), .B1(new_n630_), .B2(G8gat), .ZN(new_n631_));
  AOI211_X1 g430(.A(KEYINPUT39), .B(new_n479_), .C1(new_n624_), .C2(new_n627_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n628_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT40), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  OAI211_X1 g434(.A(KEYINPUT40), .B(new_n628_), .C1(new_n631_), .C2(new_n632_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(G1325gat));
  INV_X1    g436(.A(G15gat), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n337_), .A2(new_n340_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n638_), .B1(new_n624_), .B2(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT41), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n613_), .A2(new_n638_), .A3(new_n639_), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n642_), .B(KEYINPUT99), .Z(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n643_), .ZN(G1326gat));
  INV_X1    g443(.A(G22gat), .ZN(new_n645_));
  INV_X1    g444(.A(new_n395_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n645_), .B1(new_n624_), .B2(new_n646_), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n647_), .B(KEYINPUT42), .Z(new_n648_));
  NOR2_X1   g447(.A1(new_n395_), .A2(G22gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT100), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n613_), .A2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n648_), .A2(new_n651_), .ZN(G1327gat));
  INV_X1    g451(.A(new_n620_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n619_), .A2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n623_), .A2(new_n521_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(G29gat), .B1(new_n656_), .B2(new_n270_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT43), .ZN(new_n658_));
  INV_X1    g457(.A(new_n582_), .ZN(new_n659_));
  AND3_X1   g458(.A1(new_n616_), .A2(new_n464_), .A3(new_n452_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n270_), .A2(new_n469_), .A3(new_n471_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n474_), .B1(new_n661_), .B2(new_n462_), .ZN(new_n662_));
  OAI211_X1 g461(.A(new_n658_), .B(new_n659_), .C1(new_n660_), .C2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(KEYINPUT102), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n582_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT102), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n665_), .A2(new_n666_), .A3(new_n658_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n664_), .A2(new_n667_), .ZN(new_n668_));
  OAI21_X1  g467(.A(KEYINPUT101), .B1(new_n665_), .B2(new_n658_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT101), .ZN(new_n670_));
  OAI211_X1 g469(.A(new_n670_), .B(KEYINPUT43), .C1(new_n476_), .C2(new_n582_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n655_), .B1(new_n668_), .B2(new_n672_), .ZN(new_n673_));
  OR2_X1    g472(.A1(new_n673_), .A2(KEYINPUT44), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n674_), .A2(G29gat), .A3(new_n270_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n655_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n668_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n672_), .ZN(new_n678_));
  OAI211_X1 g477(.A(KEYINPUT44), .B(new_n676_), .C1(new_n677_), .C2(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n657_), .B1(new_n675_), .B2(new_n679_), .ZN(G1328gat));
  NAND3_X1  g479(.A1(new_n674_), .A2(new_n627_), .A3(new_n679_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(G36gat), .ZN(new_n682_));
  OR2_X1    g481(.A1(new_n452_), .A2(KEYINPUT103), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n452_), .A2(KEYINPUT103), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NOR4_X1   g484(.A1(new_n654_), .A2(new_n655_), .A3(G36gat), .A4(new_n685_), .ZN(new_n686_));
  XOR2_X1   g485(.A(new_n686_), .B(KEYINPUT45), .Z(new_n687_));
  NAND2_X1  g486(.A1(new_n682_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT46), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n682_), .A2(KEYINPUT46), .A3(new_n687_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1329gat));
  NAND4_X1  g491(.A1(new_n674_), .A2(G43gat), .A3(new_n396_), .A4(new_n679_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n639_), .ZN(new_n694_));
  NOR3_X1   g493(.A1(new_n654_), .A2(new_n655_), .A3(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n693_), .B1(G43gat), .B2(new_n695_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g496(.A(G50gat), .B1(new_n656_), .B2(new_n646_), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n674_), .A2(G50gat), .A3(new_n679_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n698_), .B1(new_n699_), .B2(new_n646_), .ZN(G1331gat));
  INV_X1    g499(.A(new_n595_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n515_), .A2(new_n516_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n507_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(KEYINPUT73), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n517_), .A2(new_n518_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n701_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n622_), .A2(new_n612_), .A3(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n709_), .A2(G57gat), .A3(new_n270_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT105), .ZN(new_n711_));
  INV_X1    g510(.A(new_n612_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n712_), .A2(new_n701_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n522_), .A2(new_n582_), .A3(new_n713_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT104), .ZN(new_n715_));
  AOI21_X1  g514(.A(G57gat), .B1(new_n715_), .B2(new_n270_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n711_), .A2(new_n716_), .ZN(G1332gat));
  OAI21_X1  g516(.A(G64gat), .B1(new_n708_), .B2(new_n685_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT48), .ZN(new_n719_));
  OR3_X1    g518(.A1(new_n714_), .A2(G64gat), .A3(new_n685_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(KEYINPUT106), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT106), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n719_), .A2(new_n723_), .A3(new_n720_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n722_), .A2(new_n724_), .ZN(G1333gat));
  OR3_X1    g524(.A1(new_n714_), .A2(G71gat), .A3(new_n694_), .ZN(new_n726_));
  OAI21_X1  g525(.A(G71gat), .B1(new_n708_), .B2(new_n694_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n727_), .A2(KEYINPUT49), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n727_), .A2(KEYINPUT49), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n726_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT107), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  OAI211_X1 g531(.A(KEYINPUT107), .B(new_n726_), .C1(new_n728_), .C2(new_n729_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1334gat));
  OAI21_X1  g533(.A(G78gat), .B1(new_n708_), .B2(new_n395_), .ZN(new_n735_));
  XOR2_X1   g534(.A(KEYINPUT108), .B(KEYINPUT50), .Z(new_n736_));
  XNOR2_X1  g535(.A(new_n735_), .B(new_n736_), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n395_), .A2(G78gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n737_), .B1(new_n714_), .B2(new_n738_), .ZN(G1335gat));
  NAND2_X1  g538(.A1(new_n713_), .A2(new_n521_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n740_), .A2(new_n654_), .ZN(new_n741_));
  AOI21_X1  g540(.A(G85gat), .B1(new_n741_), .B2(new_n270_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n740_), .B1(new_n668_), .B2(new_n672_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n270_), .A2(G85gat), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n742_), .B1(new_n743_), .B2(new_n744_), .ZN(G1336gat));
  AOI21_X1  g544(.A(G92gat), .B1(new_n741_), .B2(new_n627_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n685_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(G92gat), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT109), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n746_), .B1(new_n743_), .B2(new_n749_), .ZN(G1337gat));
  INV_X1    g549(.A(KEYINPUT110), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n539_), .B1(new_n743_), .B2(new_n639_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n741_), .A2(new_n527_), .A3(new_n396_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n751_), .B1(new_n752_), .B2(new_n754_), .ZN(new_n755_));
  AOI211_X1 g554(.A(new_n694_), .B(new_n740_), .C1(new_n668_), .C2(new_n672_), .ZN(new_n756_));
  OAI211_X1 g555(.A(KEYINPUT110), .B(new_n753_), .C1(new_n756_), .C2(new_n539_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n755_), .A2(KEYINPUT51), .A3(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT111), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n755_), .A2(KEYINPUT111), .A3(new_n757_), .A4(KEYINPUT51), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  NOR3_X1   g561(.A1(new_n752_), .A2(KEYINPUT51), .A3(new_n754_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT112), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n763_), .B(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n762_), .A2(new_n765_), .ZN(G1338gat));
  NAND3_X1  g565(.A1(new_n741_), .A2(new_n528_), .A3(new_n646_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n743_), .A2(new_n646_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n768_), .B1(new_n769_), .B2(G106gat), .ZN(new_n770_));
  AOI211_X1 g569(.A(KEYINPUT52), .B(new_n528_), .C1(new_n743_), .C2(new_n646_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n767_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g572(.A1(new_n627_), .A2(new_n464_), .A3(new_n397_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT57), .ZN(new_n776_));
  NOR3_X1   g575(.A1(new_n603_), .A2(new_n604_), .A3(new_n610_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n595_), .A2(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n600_), .A2(new_n597_), .A3(new_n602_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT55), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n603_), .A2(new_n780_), .ZN(new_n781_));
  AOI211_X1 g580(.A(KEYINPUT55), .B(new_n597_), .C1(new_n600_), .C2(new_n602_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n779_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n783_), .A2(KEYINPUT56), .A3(new_n610_), .ZN(new_n784_));
  AOI21_X1  g583(.A(KEYINPUT56), .B1(new_n783_), .B2(new_n610_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n778_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n562_), .A2(new_n485_), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n787_), .B(KEYINPUT116), .C1(new_n485_), .C2(new_n558_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT116), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n789_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n788_), .A2(new_n790_), .A3(new_n587_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n593_), .B1(new_n589_), .B2(new_n586_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT117), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n590_), .A2(new_n593_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT117), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n791_), .A2(new_n796_), .A3(new_n792_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n794_), .A2(new_n795_), .A3(new_n797_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n611_), .A2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n786_), .A2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(new_n620_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n776_), .B1(new_n802_), .B2(KEYINPUT118), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n653_), .B1(new_n786_), .B2(new_n800_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT118), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n804_), .A2(new_n805_), .A3(KEYINPUT57), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n803_), .A2(new_n806_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n798_), .A2(new_n777_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT119), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n808_), .B(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n783_), .A2(KEYINPUT56), .A3(new_n610_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n811_), .B1(new_n785_), .B2(KEYINPUT120), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT120), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n783_), .A2(new_n813_), .A3(KEYINPUT56), .A4(new_n610_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n810_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT58), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n582_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n810_), .A2(new_n815_), .A3(KEYINPUT58), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT121), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT121), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n810_), .A2(new_n815_), .A3(new_n821_), .A4(KEYINPUT58), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n818_), .A2(new_n820_), .A3(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n807_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT122), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n807_), .A2(new_n823_), .A3(KEYINPUT122), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(new_n704_), .A3(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n707_), .A2(new_n712_), .A3(KEYINPUT113), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT113), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n595_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n830_), .B1(new_n831_), .B2(new_n612_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n829_), .A2(new_n832_), .A3(new_n582_), .ZN(new_n833_));
  XOR2_X1   g632(.A(KEYINPUT114), .B(KEYINPUT54), .Z(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT115), .ZN(new_n836_));
  OR2_X1    g635(.A1(new_n833_), .A2(new_n834_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT115), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n833_), .A2(new_n838_), .A3(new_n834_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n836_), .A2(new_n837_), .A3(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n775_), .B1(new_n828_), .B2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(G113gat), .B1(new_n841_), .B2(new_n701_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n841_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n521_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n824_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n840_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n775_), .A2(KEYINPUT59), .ZN(new_n847_));
  AOI22_X1  g646(.A1(new_n843_), .A2(KEYINPUT59), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n595_), .A2(new_n223_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n842_), .B1(new_n848_), .B2(new_n849_), .ZN(G1340gat));
  NAND2_X1  g649(.A1(new_n846_), .A2(new_n847_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT59), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n612_), .B(new_n851_), .C1(new_n841_), .C2(new_n852_), .ZN(new_n853_));
  AND3_X1   g652(.A1(new_n836_), .A2(new_n837_), .A3(new_n839_), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n807_), .A2(new_n823_), .A3(KEYINPUT122), .ZN(new_n855_));
  AOI21_X1  g654(.A(KEYINPUT122), .B1(new_n807_), .B2(new_n823_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n854_), .B1(new_n857_), .B2(new_n704_), .ZN(new_n858_));
  AOI21_X1  g657(.A(KEYINPUT60), .B1(new_n612_), .B2(new_n224_), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n858_), .A2(new_n775_), .A3(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(G120gat), .B1(new_n853_), .B2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT60), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n863_), .ZN(G1341gat));
  AOI21_X1  g663(.A(G127gat), .B1(new_n841_), .B2(new_n844_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n704_), .A2(new_n218_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n865_), .B1(new_n848_), .B2(new_n866_), .ZN(G1342gat));
  AOI21_X1  g666(.A(G134gat), .B1(new_n841_), .B2(new_n653_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n582_), .A2(new_n219_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n868_), .B1(new_n848_), .B2(new_n869_), .ZN(G1343gat));
  AOI21_X1  g669(.A(new_n394_), .B1(new_n828_), .B2(new_n840_), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n871_), .A2(new_n270_), .A3(new_n701_), .A4(new_n685_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(G141gat), .ZN(G1344gat));
  NAND4_X1  g672(.A1(new_n871_), .A2(new_n270_), .A3(new_n612_), .A4(new_n685_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(G148gat), .ZN(G1345gat));
  NAND4_X1  g674(.A1(new_n871_), .A2(new_n270_), .A3(new_n844_), .A4(new_n685_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(KEYINPUT61), .B(G155gat), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n876_), .B(new_n877_), .ZN(G1346gat));
  INV_X1    g677(.A(new_n871_), .ZN(new_n879_));
  NOR3_X1   g678(.A1(new_n879_), .A2(new_n464_), .A3(new_n747_), .ZN(new_n880_));
  INV_X1    g679(.A(G162gat), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n582_), .A2(new_n881_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(KEYINPUT123), .ZN(new_n883_));
  NAND4_X1  g682(.A1(new_n871_), .A2(new_n270_), .A3(new_n653_), .A4(new_n685_), .ZN(new_n884_));
  AOI22_X1  g683(.A1(new_n880_), .A2(new_n883_), .B1(new_n881_), .B2(new_n884_), .ZN(G1347gat));
  NOR2_X1   g684(.A1(new_n685_), .A2(new_n270_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n887_), .A2(new_n694_), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n846_), .A2(new_n395_), .A3(new_n701_), .A4(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(G169gat), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT62), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n890_), .A2(KEYINPUT124), .A3(new_n891_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n846_), .A2(new_n395_), .A3(new_n888_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n894_), .A2(new_n312_), .A3(new_n701_), .ZN(new_n895_));
  OR2_X1    g694(.A1(new_n891_), .A2(KEYINPUT124), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n891_), .A2(KEYINPUT124), .ZN(new_n897_));
  NAND4_X1  g696(.A1(new_n889_), .A2(G169gat), .A3(new_n896_), .A4(new_n897_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n892_), .A2(new_n895_), .A3(new_n898_), .ZN(G1348gat));
  AOI22_X1  g698(.A1(new_n894_), .A2(new_n612_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n828_), .A2(new_n840_), .ZN(new_n901_));
  AOI21_X1  g700(.A(KEYINPUT125), .B1(new_n901_), .B2(new_n395_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT125), .ZN(new_n903_));
  AOI211_X1 g702(.A(new_n903_), .B(new_n646_), .C1(new_n828_), .C2(new_n840_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n888_), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n902_), .A2(new_n904_), .A3(new_n905_), .ZN(new_n906_));
  AND2_X1   g705(.A1(new_n612_), .A2(G176gat), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n900_), .B1(new_n906_), .B2(new_n907_), .ZN(G1349gat));
  NOR3_X1   g707(.A1(new_n893_), .A2(new_n704_), .A3(new_n299_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n903_), .B1(new_n858_), .B2(new_n646_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n901_), .A2(KEYINPUT125), .A3(new_n395_), .ZN(new_n911_));
  NAND4_X1  g710(.A1(new_n910_), .A2(new_n844_), .A3(new_n888_), .A4(new_n911_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n909_), .B1(new_n912_), .B2(new_n284_), .ZN(G1350gat));
  OAI21_X1  g712(.A(G190gat), .B1(new_n893_), .B2(new_n582_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n653_), .A2(new_n300_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(KEYINPUT126), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n914_), .B1(new_n893_), .B2(new_n916_), .ZN(G1351gat));
  NAND3_X1  g716(.A1(new_n871_), .A2(new_n701_), .A3(new_n886_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g718(.A1(new_n871_), .A2(new_n612_), .A3(new_n886_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g720(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n922_));
  NAND4_X1  g721(.A1(new_n871_), .A2(new_n517_), .A3(new_n886_), .A4(new_n922_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n924_));
  XOR2_X1   g723(.A(new_n924_), .B(KEYINPUT127), .Z(new_n925_));
  XNOR2_X1  g724(.A(new_n923_), .B(new_n925_), .ZN(G1354gat));
  NOR2_X1   g725(.A1(new_n879_), .A2(new_n887_), .ZN(new_n927_));
  INV_X1    g726(.A(G218gat), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n582_), .A2(new_n928_), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n871_), .A2(new_n653_), .A3(new_n886_), .ZN(new_n930_));
  AOI22_X1  g729(.A1(new_n927_), .A2(new_n929_), .B1(new_n930_), .B2(new_n928_), .ZN(G1355gat));
endmodule


