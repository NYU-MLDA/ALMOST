//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 1 1 0 0 1 0 0 1 0 0 0 0 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 0 1 1 0 1 1 0 0 1 0 0 1 0 0 0 1 0 0 1 1 1 1 1 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n808_,
    new_n809_, new_n810_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n823_, new_n824_, new_n825_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n863_, new_n864_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n935_, new_n936_, new_n937_, new_n939_,
    new_n940_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n956_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n974_,
    new_n975_, new_n976_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n989_, new_n990_, new_n992_, new_n993_, new_n994_, new_n995_,
    new_n997_, new_n998_, new_n999_, new_n1001_, new_n1002_, new_n1003_,
    new_n1005_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1012_, new_n1013_, new_n1015_, new_n1016_, new_n1017_;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT32), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G226gat), .A2(G233gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT19), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  OR2_X1    g010(.A1(KEYINPUT83), .A2(G169gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(KEYINPUT83), .A2(G169gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NOR2_X1   g013(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n212_), .A2(new_n215_), .A3(new_n213_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G183gat), .A2(G190gat), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G183gat), .A2(G190gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT81), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT81), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n225_), .A2(G183gat), .A3(G190gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n222_), .B1(new_n227_), .B2(KEYINPUT23), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n219_), .B1(new_n221_), .B2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT79), .ZN(new_n230_));
  INV_X1    g029(.A(G169gat), .ZN(new_n231_));
  INV_X1    g030(.A(G176gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n230_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT79), .B1(G169gat), .B2(G176gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G169gat), .A2(G176gat), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n233_), .A2(KEYINPUT24), .A3(new_n234_), .A4(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(KEYINPUT26), .B(G190gat), .ZN(new_n237_));
  INV_X1    g036(.A(G183gat), .ZN(new_n238_));
  OAI21_X1  g037(.A(KEYINPUT78), .B1(new_n238_), .B2(KEYINPUT25), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT25), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(G183gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n238_), .A2(KEYINPUT25), .ZN(new_n243_));
  AOI21_X1  g042(.A(KEYINPUT78), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n236_), .B1(new_n240_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT24), .ZN(new_n246_));
  INV_X1    g045(.A(new_n234_), .ZN(new_n247_));
  NOR3_X1   g046(.A1(KEYINPUT79), .A2(G169gat), .A3(G176gat), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n246_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n223_), .A2(KEYINPUT23), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT80), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT80), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n223_), .A2(new_n252_), .A3(KEYINPUT23), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(KEYINPUT23), .B1(new_n224_), .B2(new_n226_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n249_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT82), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n245_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  OAI211_X1 g057(.A(KEYINPUT82), .B(new_n249_), .C1(new_n254_), .C2(new_n255_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n229_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(G197gat), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n261_), .A2(KEYINPUT91), .A3(G204gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G197gat), .B(G204gat), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  OAI211_X1 g063(.A(KEYINPUT21), .B(new_n262_), .C1(new_n264_), .C2(KEYINPUT91), .ZN(new_n265_));
  XOR2_X1   g064(.A(G211gat), .B(G218gat), .Z(new_n266_));
  INV_X1    g065(.A(KEYINPUT21), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n266_), .B1(new_n267_), .B2(new_n263_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n263_), .A2(new_n267_), .ZN(new_n269_));
  AOI22_X1  g068(.A1(new_n265_), .A2(new_n268_), .B1(new_n266_), .B2(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT93), .B1(new_n260_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n229_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n244_), .ZN(new_n273_));
  INV_X1    g072(.A(G190gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT26), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT26), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(G190gat), .ZN(new_n277_));
  AND3_X1   g076(.A1(new_n239_), .A2(new_n275_), .A3(new_n277_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n247_), .A2(new_n248_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n235_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n280_), .A2(new_n246_), .ZN(new_n281_));
  AOI22_X1  g080(.A1(new_n273_), .A2(new_n278_), .B1(new_n279_), .B2(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(KEYINPUT24), .B1(new_n233_), .B2(new_n234_), .ZN(new_n283_));
  AND3_X1   g082(.A1(new_n223_), .A2(new_n252_), .A3(KEYINPUT23), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n252_), .B1(new_n223_), .B2(KEYINPUT23), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT23), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n227_), .A2(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n283_), .B1(new_n286_), .B2(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n282_), .B1(new_n289_), .B2(KEYINPUT82), .ZN(new_n290_));
  INV_X1    g089(.A(new_n259_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n272_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT93), .ZN(new_n293_));
  INV_X1    g092(.A(new_n270_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n292_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n271_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n242_), .A2(new_n243_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT92), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT92), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n242_), .A2(new_n243_), .A3(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n298_), .A2(new_n300_), .A3(new_n237_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n246_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n301_), .A2(new_n228_), .A3(new_n236_), .A4(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n221_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT22), .B(G169gat), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n280_), .B1(new_n305_), .B2(new_n232_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n303_), .A2(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n308_), .A2(new_n294_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT20), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n211_), .B1(new_n296_), .B2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n260_), .A2(new_n270_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n310_), .B1(new_n308_), .B2(new_n294_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n315_), .A2(new_n210_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n208_), .B1(new_n312_), .B2(new_n316_), .ZN(new_n317_));
  OAI211_X1 g116(.A(KEYINPUT20), .B(new_n211_), .C1(new_n308_), .C2(new_n294_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n296_), .A2(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n211_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n320_), .A2(new_n322_), .A3(new_n207_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT87), .ZN(new_n324_));
  INV_X1    g123(.A(G134gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(G127gat), .ZN(new_n326_));
  INV_X1    g125(.A(G127gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(G134gat), .ZN(new_n328_));
  AND3_X1   g127(.A1(new_n326_), .A2(new_n328_), .A3(KEYINPUT86), .ZN(new_n329_));
  AOI21_X1  g128(.A(KEYINPUT86), .B1(new_n326_), .B2(new_n328_), .ZN(new_n330_));
  INV_X1    g129(.A(G120gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(G113gat), .ZN(new_n332_));
  INV_X1    g131(.A(G113gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(G120gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  NOR3_X1   g134(.A1(new_n329_), .A2(new_n330_), .A3(new_n335_), .ZN(new_n336_));
  AND2_X1   g135(.A1(new_n332_), .A2(new_n334_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT86), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n327_), .A2(G134gat), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n325_), .A2(G127gat), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n338_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n326_), .A2(new_n328_), .A3(KEYINPUT86), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n337_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n324_), .B1(new_n336_), .B2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT88), .ZN(new_n345_));
  OR2_X1    g144(.A1(G155gat), .A2(G162gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G155gat), .A2(G162gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NOR3_X1   g149(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n348_), .B1(new_n352_), .B2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(G141gat), .ZN(new_n358_));
  INV_X1    g157(.A(G148gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G141gat), .A2(G148gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(G155gat), .A2(G162gat), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n363_), .B1(KEYINPUT1), .B2(new_n347_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT1), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n365_), .A2(G155gat), .A3(G162gat), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n362_), .B1(new_n364_), .B2(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n345_), .B1(new_n357_), .B2(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n335_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n341_), .A2(new_n342_), .A3(new_n337_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n369_), .A2(new_n370_), .A3(KEYINPUT87), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT3), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n372_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT2), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n361_), .A2(new_n374_), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n373_), .A2(new_n375_), .A3(new_n353_), .A4(new_n349_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n348_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n347_), .A2(KEYINPUT1), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n379_), .A2(new_n366_), .A3(new_n346_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n380_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n378_), .A2(new_n381_), .A3(KEYINPUT88), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n344_), .A2(new_n368_), .A3(new_n371_), .A4(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G225gat), .A2(G233gat), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n357_), .A2(new_n367_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n385_), .B1(new_n336_), .B2(new_n343_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n383_), .A2(new_n384_), .A3(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT96), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT94), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n390_), .B1(new_n383_), .B2(KEYINPUT4), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n369_), .A2(KEYINPUT87), .A3(new_n370_), .ZN(new_n392_));
  AOI21_X1  g191(.A(KEYINPUT87), .B1(new_n369_), .B2(new_n370_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT4), .ZN(new_n395_));
  AND3_X1   g194(.A1(new_n378_), .A2(new_n381_), .A3(KEYINPUT88), .ZN(new_n396_));
  AOI21_X1  g195(.A(KEYINPUT88), .B1(new_n378_), .B2(new_n381_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n394_), .A2(KEYINPUT94), .A3(new_n395_), .A4(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n391_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n384_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n383_), .A2(KEYINPUT4), .A3(new_n386_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n400_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  XOR2_X1   g202(.A(G1gat), .B(G29gat), .Z(new_n404_));
  XNOR2_X1  g203(.A(KEYINPUT95), .B(G85gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT0), .B(G57gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  AND3_X1   g207(.A1(new_n389_), .A2(new_n403_), .A3(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n408_), .B1(new_n389_), .B2(new_n403_), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n317_), .B(new_n323_), .C1(new_n409_), .C2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n389_), .A2(new_n403_), .A3(new_n408_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT33), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n389_), .A2(new_n403_), .A3(KEYINPUT33), .A4(new_n408_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n400_), .A2(new_n384_), .A3(new_n402_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n408_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n383_), .A2(new_n401_), .A3(new_n386_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n417_), .A2(new_n418_), .A3(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n320_), .A2(new_n206_), .A3(new_n322_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n318_), .B1(new_n271_), .B2(new_n295_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n205_), .B1(new_n422_), .B2(new_n321_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n420_), .A2(new_n421_), .A3(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n411_), .B1(new_n416_), .B2(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(KEYINPUT84), .B(KEYINPUT30), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  XOR2_X1   g226(.A(KEYINPUT85), .B(G43gat), .Z(new_n428_));
  AOI211_X1 g227(.A(new_n428_), .B(new_n229_), .C1(new_n258_), .C2(new_n259_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n428_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n256_), .A2(new_n257_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n431_), .A2(new_n259_), .A3(new_n282_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n430_), .B1(new_n432_), .B2(new_n272_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n427_), .B1(new_n429_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n292_), .A2(new_n428_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n432_), .A2(new_n272_), .A3(new_n430_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n435_), .A2(new_n426_), .A3(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G227gat), .A2(G233gat), .ZN(new_n438_));
  INV_X1    g237(.A(G15gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n438_), .B(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(G71gat), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  AND3_X1   g241(.A1(new_n434_), .A2(new_n437_), .A3(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n442_), .B1(new_n434_), .B2(new_n437_), .ZN(new_n444_));
  OAI21_X1  g243(.A(KEYINPUT31), .B1(new_n392_), .B2(new_n393_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  NOR3_X1   g245(.A1(new_n392_), .A2(new_n393_), .A3(KEYINPUT31), .ZN(new_n447_));
  OAI21_X1  g246(.A(G99gat), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n447_), .ZN(new_n449_));
  INV_X1    g248(.A(G99gat), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n449_), .A2(new_n450_), .A3(new_n445_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n448_), .A2(new_n451_), .ZN(new_n452_));
  NOR3_X1   g251(.A1(new_n443_), .A2(new_n444_), .A3(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n452_), .ZN(new_n454_));
  NOR3_X1   g253(.A1(new_n429_), .A2(new_n433_), .A3(new_n427_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n426_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n441_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n434_), .A2(new_n437_), .A3(new_n442_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n454_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G22gat), .B(G50gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(KEYINPUT90), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n461_), .B1(new_n398_), .B2(KEYINPUT29), .ZN(new_n462_));
  XOR2_X1   g261(.A(KEYINPUT89), .B(KEYINPUT28), .Z(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n368_), .A2(new_n382_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT29), .ZN(new_n466_));
  INV_X1    g265(.A(new_n461_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n465_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n462_), .A2(new_n464_), .A3(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n464_), .B1(new_n462_), .B2(new_n468_), .ZN(new_n471_));
  INV_X1    g270(.A(G228gat), .ZN(new_n472_));
  INV_X1    g271(.A(G233gat), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  OAI211_X1 g274(.A(new_n294_), .B(new_n475_), .C1(new_n465_), .C2(new_n466_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n385_), .A2(new_n466_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n474_), .B1(new_n477_), .B2(new_n270_), .ZN(new_n478_));
  XOR2_X1   g277(.A(G78gat), .B(G106gat), .Z(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  AND3_X1   g279(.A1(new_n476_), .A2(new_n478_), .A3(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n480_), .B1(new_n476_), .B2(new_n478_), .ZN(new_n482_));
  OAI22_X1  g281(.A1(new_n470_), .A2(new_n471_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n482_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n462_), .A2(new_n468_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(new_n463_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n476_), .A2(new_n480_), .A3(new_n478_), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n484_), .A2(new_n486_), .A3(new_n469_), .A4(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n483_), .A2(new_n488_), .ZN(new_n489_));
  NOR3_X1   g288(.A1(new_n453_), .A2(new_n459_), .A3(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n425_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT97), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n421_), .A2(new_n492_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n205_), .B1(new_n312_), .B2(new_n316_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n492_), .B(new_n205_), .C1(new_n312_), .C2(new_n316_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n495_), .A2(KEYINPUT27), .A3(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT98), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n421_), .A2(new_n423_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT27), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n498_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  AOI211_X1 g300(.A(KEYINPUT98), .B(KEYINPUT27), .C1(new_n421_), .C2(new_n423_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n497_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n409_), .A2(new_n410_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n452_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n457_), .A2(new_n454_), .A3(new_n458_), .ZN(new_n506_));
  AND3_X1   g305(.A1(new_n505_), .A2(new_n489_), .A3(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n489_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n504_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n491_), .B1(new_n503_), .B2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G99gat), .A2(G106gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT6), .ZN(new_n512_));
  INV_X1    g311(.A(G85gat), .ZN(new_n513_));
  INV_X1    g312(.A(G92gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G85gat), .A2(G92gat), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n515_), .A2(KEYINPUT9), .A3(new_n516_), .ZN(new_n517_));
  OR2_X1    g316(.A1(new_n516_), .A2(KEYINPUT9), .ZN(new_n518_));
  AND3_X1   g317(.A1(new_n512_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(KEYINPUT10), .B(G99gat), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT64), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  OR2_X1    g321(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n523_), .A2(KEYINPUT64), .A3(new_n524_), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n522_), .A2(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n519_), .B1(new_n526_), .B2(G106gat), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT8), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT66), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NOR3_X1   g330(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n529_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT7), .ZN(new_n534_));
  INV_X1    g333(.A(G106gat), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(new_n450_), .A3(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n536_), .A2(KEYINPUT66), .A3(new_n530_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n533_), .A2(new_n512_), .A3(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n516_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(G85gat), .A2(G92gat), .ZN(new_n540_));
  OAI21_X1  g339(.A(KEYINPUT65), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT65), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n515_), .A2(new_n542_), .A3(new_n516_), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n541_), .A2(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n528_), .B1(new_n538_), .B2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n541_), .A2(new_n543_), .A3(new_n528_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n531_), .A2(new_n532_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n546_), .B1(new_n512_), .B2(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n527_), .B1(new_n545_), .B2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G57gat), .B(G64gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G71gat), .B(G78gat), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n550_), .A2(new_n551_), .A3(KEYINPUT11), .ZN(new_n552_));
  XOR2_X1   g351(.A(G71gat), .B(G78gat), .Z(new_n553_));
  INV_X1    g352(.A(G64gat), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(G57gat), .ZN(new_n555_));
  INV_X1    g354(.A(G57gat), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(G64gat), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n555_), .A2(new_n557_), .A3(KEYINPUT11), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n553_), .A2(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n550_), .A2(KEYINPUT11), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n552_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n549_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT12), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G230gat), .A2(G233gat), .ZN(new_n566_));
  OAI211_X1 g365(.A(new_n527_), .B(new_n561_), .C1(new_n545_), .C2(new_n548_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT67), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n519_), .B(new_n568_), .C1(new_n526_), .C2(G106gat), .ZN(new_n569_));
  AOI21_X1  g368(.A(G106gat), .B1(new_n522_), .B2(new_n525_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n512_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n571_));
  OAI21_X1  g370(.A(KEYINPUT67), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  OAI211_X1 g371(.A(new_n569_), .B(new_n572_), .C1(new_n545_), .C2(new_n548_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n561_), .A2(KEYINPUT68), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT68), .ZN(new_n575_));
  OAI211_X1 g374(.A(new_n575_), .B(new_n552_), .C1(new_n559_), .C2(new_n560_), .ZN(new_n576_));
  AND3_X1   g375(.A1(new_n574_), .A2(KEYINPUT12), .A3(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n573_), .A2(new_n577_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n565_), .A2(new_n566_), .A3(new_n567_), .A4(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n563_), .A2(new_n567_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n566_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G120gat), .B(G148gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT5), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G176gat), .B(G204gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n579_), .A2(new_n582_), .A3(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT69), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n579_), .A2(KEYINPUT69), .A3(new_n582_), .A4(new_n586_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n579_), .A2(new_n582_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n586_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n591_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT13), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n591_), .A2(KEYINPUT13), .A3(new_n594_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT70), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(G229gat), .A2(G233gat), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G1gat), .B(G8gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(KEYINPUT72), .B(G1gat), .ZN(new_n605_));
  INV_X1    g404(.A(G8gat), .ZN(new_n606_));
  OAI21_X1  g405(.A(KEYINPUT14), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G15gat), .B(G22gat), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(KEYINPUT73), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT73), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n607_), .A2(new_n611_), .A3(new_n608_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n604_), .B1(new_n610_), .B2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n610_), .A2(new_n612_), .A3(new_n604_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G29gat), .B(G36gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G43gat), .B(G50gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n616_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n616_), .A2(new_n620_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n603_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n615_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n625_), .A2(new_n613_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(new_n619_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n619_), .B(KEYINPUT15), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n616_), .A2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n627_), .A2(new_n629_), .A3(new_n602_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(G113gat), .B(G141gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(G169gat), .B(G197gat), .ZN(new_n632_));
  XOR2_X1   g431(.A(new_n631_), .B(new_n632_), .Z(new_n633_));
  NAND3_X1  g432(.A1(new_n624_), .A2(new_n630_), .A3(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n633_), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n627_), .A2(new_n629_), .A3(new_n602_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n602_), .B1(new_n627_), .B2(new_n621_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n635_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n634_), .A2(new_n638_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n574_), .A2(new_n576_), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT75), .Z(new_n641_));
  NAND2_X1  g440(.A1(G231gat), .A2(G233gat), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n642_), .B(KEYINPUT74), .Z(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n616_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n626_), .A2(new_n643_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n641_), .A2(new_n645_), .A3(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n645_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n640_), .B(KEYINPUT75), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(G127gat), .B(G155gat), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT16), .ZN(new_n652_));
  XNOR2_X1  g451(.A(G183gat), .B(G211gat), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n652_), .B(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(KEYINPUT17), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT76), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n647_), .A2(new_n650_), .A3(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n648_), .A2(new_n562_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n646_), .A2(new_n645_), .A3(new_n561_), .ZN(new_n659_));
  XOR2_X1   g458(.A(new_n654_), .B(KEYINPUT17), .Z(new_n660_));
  NAND3_X1  g459(.A1(new_n658_), .A2(new_n659_), .A3(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT77), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n657_), .A2(new_n661_), .A3(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n662_), .B1(new_n657_), .B2(new_n661_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  OR2_X1    g465(.A1(new_n549_), .A2(new_n620_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n573_), .A2(new_n628_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n669_));
  NAND2_X1  g468(.A1(G232gat), .A2(G233gat), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n669_), .B(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT35), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n667_), .A2(new_n668_), .A3(new_n674_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n672_), .A2(new_n673_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(G190gat), .B(G218gat), .ZN(new_n678_));
  XNOR2_X1  g477(.A(G134gat), .B(G162gat), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n678_), .B(new_n679_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n680_), .A2(KEYINPUT36), .ZN(new_n681_));
  INV_X1    g480(.A(new_n676_), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n667_), .A2(new_n668_), .A3(new_n682_), .A4(new_n674_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n677_), .A2(new_n681_), .A3(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  XOR2_X1   g484(.A(new_n680_), .B(KEYINPUT36), .Z(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n687_), .B1(new_n677_), .B2(new_n683_), .ZN(new_n688_));
  OAI21_X1  g487(.A(KEYINPUT37), .B1(new_n685_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n688_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT37), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n690_), .A2(new_n691_), .A3(new_n684_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n689_), .A2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n666_), .A2(new_n694_), .ZN(new_n695_));
  AND4_X1   g494(.A1(new_n510_), .A2(new_n601_), .A3(new_n639_), .A4(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n504_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n696_), .A2(new_n697_), .A3(new_n605_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT38), .ZN(new_n699_));
  OR2_X1    g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n639_), .ZN(new_n701_));
  OR3_X1    g500(.A1(new_n599_), .A2(KEYINPUT99), .A3(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(KEYINPUT99), .B1(new_n599_), .B2(new_n701_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n685_), .A2(new_n688_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n666_), .A2(new_n704_), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n702_), .A2(new_n510_), .A3(new_n703_), .A4(new_n705_), .ZN(new_n706_));
  OAI21_X1  g505(.A(G1gat), .B1(new_n706_), .B2(new_n504_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n698_), .A2(new_n699_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n700_), .A2(new_n707_), .A3(new_n708_), .ZN(G1324gat));
  INV_X1    g508(.A(KEYINPUT39), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n206_), .B1(new_n320_), .B2(new_n322_), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n422_), .A2(new_n205_), .A3(new_n321_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n500_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(KEYINPUT98), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n499_), .A2(new_n498_), .A3(new_n500_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n500_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n716_));
  AOI22_X1  g515(.A1(new_n714_), .A2(new_n715_), .B1(new_n716_), .B2(new_n496_), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n710_), .B(G8gat), .C1(new_n706_), .C2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT101), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n718_), .B(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT100), .ZN(new_n721_));
  OR2_X1    g520(.A1(new_n706_), .A2(new_n717_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(G8gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n721_), .B1(new_n723_), .B2(KEYINPUT39), .ZN(new_n724_));
  AOI211_X1 g523(.A(KEYINPUT100), .B(new_n710_), .C1(new_n722_), .C2(G8gat), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n720_), .A2(new_n724_), .A3(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT40), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n717_), .A2(G8gat), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n696_), .A2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  OR3_X1    g529(.A1(new_n726_), .A2(new_n727_), .A3(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n727_), .B1(new_n726_), .B2(new_n730_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(G1325gat));
  NOR2_X1   g532(.A1(new_n453_), .A2(new_n459_), .ZN(new_n734_));
  OAI21_X1  g533(.A(G15gat), .B1(new_n706_), .B2(new_n734_), .ZN(new_n735_));
  XOR2_X1   g534(.A(new_n735_), .B(KEYINPUT41), .Z(new_n736_));
  INV_X1    g535(.A(new_n734_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n696_), .A2(new_n439_), .A3(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(G1326gat));
  INV_X1    g538(.A(new_n489_), .ZN(new_n740_));
  OAI21_X1  g539(.A(G22gat), .B1(new_n706_), .B2(new_n740_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n741_), .B(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(G22gat), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n696_), .A2(new_n744_), .A3(new_n489_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1327gat));
  INV_X1    g545(.A(new_n599_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n704_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n665_), .A2(new_n748_), .ZN(new_n749_));
  AND4_X1   g548(.A1(new_n510_), .A2(new_n639_), .A3(new_n747_), .A4(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(G29gat), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n750_), .A2(new_n751_), .A3(new_n697_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n702_), .A2(new_n703_), .A3(new_n666_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n510_), .A2(new_n694_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT103), .ZN(new_n756_));
  AOI21_X1  g555(.A(KEYINPUT43), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT43), .ZN(new_n758_));
  AOI211_X1 g557(.A(KEYINPUT103), .B(new_n758_), .C1(new_n510_), .C2(new_n694_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n754_), .B1(new_n757_), .B2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT104), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT44), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n740_), .B1(new_n453_), .B2(new_n459_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n505_), .A2(new_n489_), .A3(new_n506_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n714_), .A2(new_n715_), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n765_), .A2(new_n766_), .A3(new_n497_), .A4(new_n504_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n693_), .B1(new_n767_), .B2(new_n491_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n758_), .B1(new_n768_), .B2(KEYINPUT103), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n697_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n770_));
  AOI22_X1  g569(.A1(new_n717_), .A2(new_n770_), .B1(new_n425_), .B2(new_n490_), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n756_), .B(KEYINPUT43), .C1(new_n771_), .C2(new_n693_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n753_), .B1(new_n769_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT104), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n761_), .A2(new_n762_), .A3(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n773_), .A2(KEYINPUT44), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n776_), .A2(new_n697_), .A3(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT105), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n778_), .A2(new_n779_), .A3(G29gat), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n779_), .B1(new_n778_), .B2(G29gat), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n752_), .B1(new_n780_), .B2(new_n781_), .ZN(G1328gat));
  INV_X1    g581(.A(G36gat), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n750_), .A2(new_n783_), .A3(new_n503_), .ZN(new_n784_));
  XOR2_X1   g583(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n785_));
  XNOR2_X1  g584(.A(new_n784_), .B(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT106), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n717_), .B1(new_n773_), .B2(KEYINPUT44), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n762_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n789_));
  AOI211_X1 g588(.A(KEYINPUT104), .B(new_n753_), .C1(new_n769_), .C2(new_n772_), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n787_), .B(new_n788_), .C1(new_n789_), .C2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(G36gat), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n787_), .B1(new_n776_), .B2(new_n788_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n786_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT46), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  OAI211_X1 g595(.A(KEYINPUT46), .B(new_n786_), .C1(new_n792_), .C2(new_n793_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(G1329gat));
  OAI211_X1 g597(.A(new_n737_), .B(new_n777_), .C1(new_n789_), .C2(new_n790_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(G43gat), .ZN(new_n800_));
  INV_X1    g599(.A(G43gat), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n750_), .A2(new_n801_), .A3(new_n737_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT47), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n800_), .A2(KEYINPUT47), .A3(new_n802_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(G1330gat));
  AOI21_X1  g606(.A(G50gat), .B1(new_n750_), .B2(new_n489_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n776_), .A2(new_n777_), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n489_), .A2(G50gat), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n808_), .B1(new_n809_), .B2(new_n810_), .ZN(G1331gat));
  NOR2_X1   g610(.A1(new_n771_), .A2(new_n639_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n812_), .A2(new_n600_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n813_), .A2(new_n705_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(G57gat), .B1(new_n815_), .B2(new_n504_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n695_), .A2(new_n599_), .ZN(new_n817_));
  OR2_X1    g616(.A1(new_n817_), .A2(KEYINPUT108), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(KEYINPUT108), .ZN(new_n819_));
  AND3_X1   g618(.A1(new_n818_), .A2(new_n812_), .A3(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n820_), .A2(new_n556_), .A3(new_n697_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n816_), .A2(new_n821_), .ZN(G1332gat));
  AOI21_X1  g621(.A(new_n554_), .B1(new_n814_), .B2(new_n503_), .ZN(new_n823_));
  XOR2_X1   g622(.A(new_n823_), .B(KEYINPUT48), .Z(new_n824_));
  NAND3_X1  g623(.A1(new_n820_), .A2(new_n554_), .A3(new_n503_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(G1333gat));
  INV_X1    g625(.A(G71gat), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n827_), .B1(new_n814_), .B2(new_n737_), .ZN(new_n828_));
  XOR2_X1   g627(.A(new_n828_), .B(KEYINPUT49), .Z(new_n829_));
  NAND3_X1  g628(.A1(new_n820_), .A2(new_n827_), .A3(new_n737_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(G1334gat));
  INV_X1    g630(.A(G78gat), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n820_), .A2(new_n832_), .A3(new_n489_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT50), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n814_), .A2(new_n489_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n834_), .B1(new_n835_), .B2(G78gat), .ZN(new_n836_));
  AOI211_X1 g635(.A(KEYINPUT50), .B(new_n832_), .C1(new_n814_), .C2(new_n489_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n833_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT109), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n838_), .B(new_n839_), .ZN(G1335gat));
  NOR2_X1   g639(.A1(new_n757_), .A2(new_n759_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n599_), .A2(new_n666_), .A3(new_n701_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n513_), .B1(new_n843_), .B2(new_n697_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n813_), .A2(new_n749_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n504_), .A2(G85gat), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n844_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n847_), .B(KEYINPUT110), .ZN(G1336gat));
  NAND3_X1  g647(.A1(new_n843_), .A2(G92gat), .A3(new_n503_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n845_), .A2(new_n503_), .ZN(new_n850_));
  AND3_X1   g649(.A1(new_n850_), .A2(KEYINPUT111), .A3(new_n514_), .ZN(new_n851_));
  AOI21_X1  g650(.A(KEYINPUT111), .B1(new_n850_), .B2(new_n514_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n849_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT112), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n853_), .B(new_n854_), .ZN(G1337gat));
  INV_X1    g654(.A(new_n845_), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n856_), .A2(new_n734_), .A3(new_n526_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n450_), .B1(new_n843_), .B2(new_n737_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT113), .ZN(new_n859_));
  OAI22_X1  g658(.A1(new_n857_), .A2(new_n858_), .B1(new_n859_), .B2(KEYINPUT51), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(KEYINPUT51), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n860_), .B(new_n861_), .ZN(G1338gat));
  XNOR2_X1  g661(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n863_));
  NOR3_X1   g662(.A1(new_n841_), .A2(new_n740_), .A3(new_n842_), .ZN(new_n864_));
  OR2_X1    g663(.A1(KEYINPUT114), .A2(KEYINPUT52), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n535_), .B1(KEYINPUT114), .B2(KEYINPUT52), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  OR3_X1    g666(.A1(new_n864_), .A2(new_n865_), .A3(new_n867_), .ZN(new_n868_));
  OAI22_X1  g667(.A1(new_n864_), .A2(new_n867_), .B1(KEYINPUT114), .B2(KEYINPUT52), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n856_), .A2(G106gat), .A3(new_n740_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n863_), .B1(new_n870_), .B2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n863_), .ZN(new_n874_));
  AOI211_X1 g673(.A(new_n871_), .B(new_n874_), .C1(new_n868_), .C2(new_n869_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n873_), .A2(new_n875_), .ZN(G1339gat));
  NAND2_X1  g675(.A1(new_n717_), .A2(new_n697_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n565_), .A2(new_n567_), .A3(new_n578_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT55), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n880_), .B1(new_n581_), .B2(KEYINPUT116), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n881_), .B1(new_n880_), .B2(new_n581_), .ZN(new_n883_));
  NAND4_X1  g682(.A1(new_n565_), .A2(new_n567_), .A3(new_n578_), .A4(new_n883_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n882_), .A2(new_n593_), .A3(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(KEYINPUT56), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT56), .ZN(new_n887_));
  NAND4_X1  g686(.A1(new_n882_), .A2(new_n887_), .A3(new_n593_), .A4(new_n884_), .ZN(new_n888_));
  AND4_X1   g687(.A1(new_n639_), .A2(new_n591_), .A3(new_n886_), .A4(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n602_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n627_), .A2(new_n629_), .A3(new_n603_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n890_), .A2(new_n635_), .A3(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n634_), .A2(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n893_), .B1(new_n591_), .B2(new_n594_), .ZN(new_n894_));
  OAI211_X1 g693(.A(KEYINPUT57), .B(new_n748_), .C1(new_n889_), .C2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT118), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(new_n897_));
  AND2_X1   g696(.A1(new_n634_), .A2(new_n892_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n595_), .A2(new_n898_), .ZN(new_n899_));
  NAND4_X1  g698(.A1(new_n639_), .A2(new_n591_), .A3(new_n886_), .A4(new_n888_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n704_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n901_), .A2(KEYINPUT118), .A3(KEYINPUT57), .ZN(new_n902_));
  NAND4_X1  g701(.A1(new_n898_), .A2(new_n591_), .A3(new_n886_), .A4(new_n888_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT58), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n693_), .B1(new_n903_), .B2(new_n904_), .ZN(new_n905_));
  AND2_X1   g704(.A1(new_n886_), .A2(new_n888_), .ZN(new_n906_));
  NAND4_X1  g705(.A1(new_n906_), .A2(KEYINPUT58), .A3(new_n591_), .A4(new_n898_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n905_), .A2(new_n907_), .ZN(new_n908_));
  AND3_X1   g707(.A1(new_n897_), .A2(new_n902_), .A3(new_n908_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n748_), .B1(new_n889_), .B2(new_n894_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT117), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT57), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n901_), .A2(KEYINPUT117), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n912_), .A2(new_n913_), .A3(new_n914_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n665_), .B1(new_n909_), .B2(new_n915_), .ZN(new_n916_));
  AND3_X1   g715(.A1(new_n665_), .A2(new_n701_), .A3(new_n693_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT54), .ZN(new_n918_));
  AND3_X1   g717(.A1(new_n917_), .A2(new_n747_), .A3(new_n918_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n918_), .B1(new_n917_), .B2(new_n747_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  OAI211_X1 g720(.A(new_n508_), .B(new_n878_), .C1(new_n916_), .C2(new_n921_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n922_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n923_), .A2(new_n333_), .A3(new_n639_), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT59), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n922_), .A2(new_n925_), .ZN(new_n926_));
  AND3_X1   g725(.A1(new_n912_), .A2(new_n913_), .A3(new_n914_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n897_), .A2(new_n902_), .A3(new_n908_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n666_), .B1(new_n927_), .B2(new_n928_), .ZN(new_n929_));
  INV_X1    g728(.A(new_n921_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n877_), .B1(new_n929_), .B2(new_n930_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n931_), .A2(KEYINPUT59), .A3(new_n508_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n701_), .B1(new_n926_), .B2(new_n932_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n924_), .B1(new_n933_), .B2(new_n333_), .ZN(G1340gat));
  AOI21_X1  g733(.A(new_n601_), .B1(new_n926_), .B2(new_n932_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n331_), .B1(new_n747_), .B2(KEYINPUT60), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n936_), .B1(KEYINPUT60), .B2(new_n331_), .ZN(new_n937_));
  OAI22_X1  g736(.A1(new_n935_), .A2(new_n331_), .B1(new_n922_), .B2(new_n937_), .ZN(G1341gat));
  NAND3_X1  g737(.A1(new_n923_), .A2(new_n327_), .A3(new_n665_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n666_), .B1(new_n926_), .B2(new_n932_), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n939_), .B1(new_n940_), .B2(new_n327_), .ZN(G1342gat));
  NAND3_X1  g740(.A1(new_n923_), .A2(new_n325_), .A3(new_n704_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n693_), .B1(new_n926_), .B2(new_n932_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n942_), .B1(new_n943_), .B2(new_n325_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n944_), .A2(KEYINPUT119), .ZN(new_n945_));
  INV_X1    g744(.A(KEYINPUT119), .ZN(new_n946_));
  OAI211_X1 g745(.A(new_n942_), .B(new_n946_), .C1(new_n943_), .C2(new_n325_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n945_), .A2(new_n947_), .ZN(G1343gat));
  OAI211_X1 g747(.A(new_n507_), .B(new_n878_), .C1(new_n916_), .C2(new_n921_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n949_), .A2(KEYINPUT120), .ZN(new_n950_));
  INV_X1    g749(.A(KEYINPUT120), .ZN(new_n951_));
  NAND3_X1  g750(.A1(new_n931_), .A2(new_n951_), .A3(new_n507_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n950_), .A2(new_n952_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n953_), .A2(new_n639_), .ZN(new_n954_));
  XNOR2_X1  g753(.A(new_n954_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g754(.A1(new_n953_), .A2(new_n600_), .ZN(new_n956_));
  XNOR2_X1  g755(.A(new_n956_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g756(.A(KEYINPUT61), .B(G155gat), .ZN(new_n958_));
  INV_X1    g757(.A(new_n958_), .ZN(new_n959_));
  INV_X1    g758(.A(KEYINPUT121), .ZN(new_n960_));
  AOI21_X1  g759(.A(new_n960_), .B1(new_n953_), .B2(new_n665_), .ZN(new_n961_));
  AOI211_X1 g760(.A(KEYINPUT121), .B(new_n666_), .C1(new_n950_), .C2(new_n952_), .ZN(new_n962_));
  OAI21_X1  g761(.A(new_n959_), .B1(new_n961_), .B2(new_n962_), .ZN(new_n963_));
  AOI21_X1  g762(.A(new_n951_), .B1(new_n931_), .B2(new_n507_), .ZN(new_n964_));
  AOI22_X1  g763(.A1(new_n895_), .A2(new_n896_), .B1(new_n905_), .B2(new_n907_), .ZN(new_n965_));
  NAND3_X1  g764(.A1(new_n915_), .A2(new_n902_), .A3(new_n965_), .ZN(new_n966_));
  AOI21_X1  g765(.A(new_n921_), .B1(new_n966_), .B2(new_n666_), .ZN(new_n967_));
  NOR4_X1   g766(.A1(new_n967_), .A2(KEYINPUT120), .A3(new_n764_), .A4(new_n877_), .ZN(new_n968_));
  OAI21_X1  g767(.A(new_n665_), .B1(new_n964_), .B2(new_n968_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n969_), .A2(KEYINPUT121), .ZN(new_n970_));
  NAND3_X1  g769(.A1(new_n953_), .A2(new_n960_), .A3(new_n665_), .ZN(new_n971_));
  NAND3_X1  g770(.A1(new_n970_), .A2(new_n958_), .A3(new_n971_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n963_), .A2(new_n972_), .ZN(G1346gat));
  INV_X1    g772(.A(new_n953_), .ZN(new_n974_));
  OR3_X1    g773(.A1(new_n974_), .A2(G162gat), .A3(new_n748_), .ZN(new_n975_));
  OAI21_X1  g774(.A(G162gat), .B1(new_n974_), .B2(new_n693_), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n975_), .A2(new_n976_), .ZN(G1347gat));
  INV_X1    g776(.A(KEYINPUT122), .ZN(new_n978_));
  NAND2_X1  g777(.A1(new_n929_), .A2(new_n930_), .ZN(new_n979_));
  NAND2_X1  g778(.A1(new_n503_), .A2(new_n504_), .ZN(new_n980_));
  NOR2_X1   g779(.A1(new_n980_), .A2(new_n763_), .ZN(new_n981_));
  NAND2_X1  g780(.A1(new_n979_), .A2(new_n981_), .ZN(new_n982_));
  NOR2_X1   g781(.A1(new_n982_), .A2(new_n701_), .ZN(new_n983_));
  OAI21_X1  g782(.A(new_n978_), .B1(new_n983_), .B2(new_n231_), .ZN(new_n984_));
  OAI211_X1 g783(.A(KEYINPUT122), .B(G169gat), .C1(new_n982_), .C2(new_n701_), .ZN(new_n985_));
  NAND3_X1  g784(.A1(new_n984_), .A2(KEYINPUT62), .A3(new_n985_), .ZN(new_n986_));
  NAND2_X1  g785(.A1(new_n983_), .A2(new_n305_), .ZN(new_n987_));
  OAI211_X1 g786(.A(new_n986_), .B(new_n987_), .C1(KEYINPUT62), .C2(new_n984_), .ZN(G1348gat));
  OAI21_X1  g787(.A(G176gat), .B1(new_n982_), .B2(new_n601_), .ZN(new_n989_));
  NAND2_X1  g788(.A1(new_n599_), .A2(new_n232_), .ZN(new_n990_));
  OAI21_X1  g789(.A(new_n989_), .B1(new_n982_), .B2(new_n990_), .ZN(G1349gat));
  OAI21_X1  g790(.A(new_n238_), .B1(new_n982_), .B2(new_n666_), .ZN(new_n992_));
  NAND2_X1  g791(.A1(new_n298_), .A2(new_n300_), .ZN(new_n993_));
  NAND4_X1  g792(.A1(new_n979_), .A2(new_n993_), .A3(new_n665_), .A4(new_n981_), .ZN(new_n994_));
  NAND2_X1  g793(.A1(new_n992_), .A2(new_n994_), .ZN(new_n995_));
  XOR2_X1   g794(.A(new_n995_), .B(KEYINPUT123), .Z(G1350gat));
  OAI21_X1  g795(.A(G190gat), .B1(new_n982_), .B2(new_n693_), .ZN(new_n997_));
  NAND2_X1  g796(.A1(new_n704_), .A2(new_n237_), .ZN(new_n998_));
  XOR2_X1   g797(.A(new_n998_), .B(KEYINPUT124), .Z(new_n999_));
  OAI21_X1  g798(.A(new_n997_), .B1(new_n982_), .B2(new_n999_), .ZN(G1351gat));
  NOR3_X1   g799(.A1(new_n967_), .A2(new_n764_), .A3(new_n980_), .ZN(new_n1001_));
  NAND2_X1  g800(.A1(new_n1001_), .A2(new_n639_), .ZN(new_n1002_));
  XNOR2_X1  g801(.A(KEYINPUT125), .B(G197gat), .ZN(new_n1003_));
  XNOR2_X1  g802(.A(new_n1002_), .B(new_n1003_), .ZN(G1352gat));
  NAND2_X1  g803(.A1(new_n1001_), .A2(new_n600_), .ZN(new_n1005_));
  XNOR2_X1  g804(.A(new_n1005_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g805(.A(new_n666_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n1007_));
  NAND2_X1  g806(.A1(new_n1001_), .A2(new_n1007_), .ZN(new_n1008_));
  INV_X1    g807(.A(KEYINPUT127), .ZN(new_n1009_));
  NOR2_X1   g808(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1010_));
  XOR2_X1   g809(.A(new_n1010_), .B(KEYINPUT126), .Z(new_n1011_));
  AOI21_X1  g810(.A(new_n1008_), .B1(new_n1009_), .B2(new_n1011_), .ZN(new_n1012_));
  XOR2_X1   g811(.A(new_n1011_), .B(KEYINPUT127), .Z(new_n1013_));
  AOI21_X1  g812(.A(new_n1012_), .B1(new_n1008_), .B2(new_n1013_), .ZN(G1354gat));
  INV_X1    g813(.A(G218gat), .ZN(new_n1015_));
  NAND3_X1  g814(.A1(new_n1001_), .A2(new_n1015_), .A3(new_n704_), .ZN(new_n1016_));
  AND2_X1   g815(.A1(new_n1001_), .A2(new_n694_), .ZN(new_n1017_));
  OAI21_X1  g816(.A(new_n1016_), .B1(new_n1017_), .B2(new_n1015_), .ZN(G1355gat));
endmodule


