//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 0 1 1 0 1 1 0 1 1 0 1 0 1 0 1 1 1 1 0 1 0 0 0 1 1 0 0 0 1 0 1 0 1 0 1 1 1 0 0 0 0 1 0 0 1 0 1 1 0 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n828_, new_n829_, new_n830_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n842_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n895_, new_n896_, new_n897_, new_n899_, new_n900_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_;
  INV_X1    g000(.A(KEYINPUT98), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G127gat), .B(G134gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G113gat), .B(G120gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT31), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G15gat), .B(G43gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT82), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT83), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G227gat), .A2(G233gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT81), .ZN(new_n211_));
  XOR2_X1   g010(.A(G71gat), .B(G99gat), .Z(new_n212_));
  XNOR2_X1  g011(.A(new_n211_), .B(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n209_), .B(new_n213_), .ZN(new_n214_));
  AND2_X1   g013(.A1(KEYINPUT77), .A2(G169gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(KEYINPUT77), .A2(G169gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT22), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(KEYINPUT78), .ZN(new_n218_));
  XOR2_X1   g017(.A(KEYINPUT79), .B(KEYINPUT22), .Z(new_n219_));
  AOI21_X1  g018(.A(G176gat), .B1(new_n219_), .B2(G169gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G183gat), .A2(G190gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n222_), .B(KEYINPUT23), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n223_), .B1(G183gat), .B2(G190gat), .ZN(new_n224_));
  INV_X1    g023(.A(G169gat), .ZN(new_n225_));
  INV_X1    g024(.A(G176gat), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n221_), .B(new_n224_), .C1(new_n225_), .C2(new_n226_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT24), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n223_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(KEYINPUT76), .A2(G183gat), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n232_), .A2(KEYINPUT25), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT26), .B(G190gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n232_), .A2(KEYINPUT25), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n233_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n225_), .A2(new_n226_), .ZN(new_n237_));
  NOR3_X1   g036(.A1(new_n237_), .A2(new_n229_), .A3(new_n228_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n231_), .A2(new_n236_), .A3(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n227_), .A2(new_n240_), .ZN(new_n241_));
  XOR2_X1   g040(.A(KEYINPUT80), .B(KEYINPUT30), .Z(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n242_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n227_), .A2(new_n240_), .A3(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n214_), .A2(new_n243_), .A3(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT84), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n214_), .A2(new_n243_), .A3(KEYINPUT84), .A4(new_n245_), .ZN(new_n249_));
  AND2_X1   g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n214_), .B1(new_n245_), .B2(new_n243_), .ZN(new_n251_));
  OAI211_X1 g050(.A(KEYINPUT85), .B(new_n206_), .C1(new_n250_), .C2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT89), .B(G197gat), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n253_), .A2(KEYINPUT90), .A3(G204gat), .ZN(new_n254_));
  INV_X1    g053(.A(G197gat), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n254_), .B1(new_n255_), .B2(G204gat), .ZN(new_n256_));
  AOI21_X1  g055(.A(KEYINPUT90), .B1(new_n253_), .B2(G204gat), .ZN(new_n257_));
  XOR2_X1   g056(.A(KEYINPUT91), .B(KEYINPUT21), .Z(new_n258_));
  OR3_X1    g057(.A1(new_n256_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G211gat), .B(G218gat), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(G204gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n253_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT21), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n264_), .B1(G197gat), .B2(G204gat), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n261_), .B1(new_n263_), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n259_), .A2(new_n266_), .ZN(new_n267_));
  OR2_X1    g066(.A1(new_n256_), .A2(new_n257_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n260_), .A2(new_n264_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n267_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G228gat), .A2(G233gat), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT29), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G141gat), .A2(G148gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT2), .ZN(new_n275_));
  OAI22_X1  g074(.A1(KEYINPUT87), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(KEYINPUT87), .A2(KEYINPUT3), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  OR2_X1    g077(.A1(G141gat), .A2(G148gat), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n279_), .A2(KEYINPUT87), .A3(KEYINPUT3), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n275_), .A2(new_n278_), .A3(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G155gat), .A2(G162gat), .ZN(new_n282_));
  NOR2_X1   g081(.A1(G155gat), .A2(G162gat), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n281_), .A2(new_n282_), .A3(new_n284_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n282_), .A2(KEYINPUT1), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n282_), .B1(new_n283_), .B2(KEYINPUT1), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n286_), .B1(new_n287_), .B2(KEYINPUT86), .ZN(new_n288_));
  AND2_X1   g087(.A1(new_n286_), .A2(KEYINPUT86), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n274_), .B(new_n279_), .C1(new_n288_), .C2(new_n289_), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n285_), .A2(new_n290_), .ZN(new_n291_));
  OAI211_X1 g090(.A(new_n271_), .B(new_n272_), .C1(new_n273_), .C2(new_n291_), .ZN(new_n292_));
  AOI22_X1  g091(.A1(new_n259_), .A2(new_n266_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n291_), .A2(new_n273_), .ZN(new_n294_));
  OAI211_X1 g093(.A(G228gat), .B(G233gat), .C1(new_n293_), .C2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G78gat), .B(G106gat), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n292_), .A2(new_n295_), .A3(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n291_), .A2(new_n273_), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n299_), .A2(KEYINPUT28), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(KEYINPUT28), .ZN(new_n301_));
  XOR2_X1   g100(.A(G22gat), .B(G50gat), .Z(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n300_), .A2(new_n301_), .A3(new_n303_), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n299_), .A2(KEYINPUT28), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n299_), .A2(KEYINPUT28), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n302_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n298_), .A2(new_n304_), .A3(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n297_), .B1(new_n292_), .B2(new_n295_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(KEYINPUT92), .ZN(new_n312_));
  AOI211_X1 g111(.A(KEYINPUT92), .B(new_n297_), .C1(new_n292_), .C2(new_n295_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n309_), .A2(new_n312_), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n206_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n251_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT85), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n316_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT88), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n307_), .A2(new_n304_), .A3(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n320_), .B1(new_n307_), .B2(new_n304_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n298_), .ZN(new_n324_));
  OAI22_X1  g123(.A1(new_n322_), .A2(new_n323_), .B1(new_n310_), .B2(new_n324_), .ZN(new_n325_));
  NAND4_X1  g124(.A1(new_n252_), .A2(new_n315_), .A3(new_n319_), .A4(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G226gat), .A2(G233gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n271_), .A2(new_n241_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT25), .B(G183gat), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n238_), .B1(new_n234_), .B2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT22), .B(G169gat), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n237_), .B1(new_n334_), .B2(new_n226_), .ZN(new_n335_));
  AOI22_X1  g134(.A1(new_n333_), .A2(new_n231_), .B1(new_n224_), .B2(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(KEYINPUT20), .B1(new_n293_), .B2(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n330_), .B1(new_n331_), .B2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n271_), .A2(new_n241_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n293_), .A2(new_n336_), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n339_), .A2(KEYINPUT20), .A3(new_n329_), .A4(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n338_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G8gat), .B(G36gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(KEYINPUT18), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G64gat), .B(G92gat), .ZN(new_n345_));
  XOR2_X1   g144(.A(new_n344_), .B(new_n345_), .Z(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n342_), .A2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n338_), .A2(new_n346_), .A3(new_n341_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G1gat), .B(G29gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT0), .ZN(new_n353_));
  INV_X1    g152(.A(G57gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(G85gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n285_), .A2(new_n290_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(new_n205_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G225gat), .A2(G233gat), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n356_), .B1(new_n358_), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n358_), .A2(KEYINPUT4), .ZN(new_n362_));
  OR3_X1    g161(.A1(new_n291_), .A2(KEYINPUT4), .A3(new_n205_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n362_), .A2(new_n359_), .A3(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n361_), .A2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT94), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n362_), .A2(new_n360_), .A3(new_n363_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n358_), .A2(new_n359_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n367_), .A2(new_n368_), .A3(new_n356_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT33), .ZN(new_n370_));
  OR2_X1    g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n369_), .A2(new_n370_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n351_), .A2(new_n366_), .A3(new_n371_), .A4(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n367_), .A2(new_n368_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n356_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(new_n369_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n329_), .B1(new_n331_), .B2(new_n337_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n339_), .A2(KEYINPUT20), .A3(new_n330_), .A4(new_n340_), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n346_), .A2(KEYINPUT32), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n378_), .A2(new_n379_), .A3(new_n380_), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n377_), .B(new_n381_), .C1(new_n342_), .C2(new_n380_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n326_), .B1(new_n373_), .B2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n252_), .A2(new_n319_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT92), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n310_), .A2(new_n385_), .ZN(new_n386_));
  NOR3_X1   g185(.A1(new_n386_), .A2(new_n308_), .A3(new_n313_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n307_), .A2(new_n304_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT88), .ZN(new_n389_));
  AOI22_X1  g188(.A1(new_n389_), .A2(new_n321_), .B1(new_n311_), .B2(new_n298_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n387_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n384_), .A2(new_n391_), .ZN(new_n392_));
  OAI211_X1 g191(.A(new_n252_), .B(new_n319_), .C1(new_n387_), .C2(new_n390_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n377_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n378_), .A2(new_n347_), .A3(new_n379_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n395_), .A2(new_n349_), .A3(KEYINPUT27), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT95), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT27), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n350_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT96), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT96), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n350_), .A2(new_n401_), .A3(new_n398_), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n397_), .A2(new_n400_), .A3(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n383_), .B1(new_n394_), .B2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G57gat), .B(G64gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(KEYINPUT11), .ZN(new_n406_));
  XOR2_X1   g205(.A(G71gat), .B(G78gat), .Z(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n405_), .A2(KEYINPUT11), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n406_), .A2(new_n407_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT12), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(KEYINPUT66), .ZN(new_n414_));
  INV_X1    g213(.A(G106gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n418_));
  NOR3_X1   g217(.A1(new_n417_), .A2(new_n418_), .A3(KEYINPUT64), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT64), .ZN(new_n420_));
  OR2_X1    g219(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n420_), .B1(new_n421_), .B2(new_n416_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n415_), .B1(new_n419_), .B2(new_n422_), .ZN(new_n423_));
  AND2_X1   g222(.A1(G85gat), .A2(G92gat), .ZN(new_n424_));
  NOR2_X1   g223(.A1(G85gat), .A2(G92gat), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT9), .ZN(new_n426_));
  NOR3_X1   g225(.A1(new_n424_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G99gat), .A2(G106gat), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT6), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n426_), .A2(G85gat), .A3(G92gat), .ZN(new_n431_));
  NAND3_X1  g230(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n430_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n427_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n423_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT7), .ZN(new_n436_));
  INV_X1    g235(.A(G99gat), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n436_), .A2(new_n437_), .A3(new_n415_), .ZN(new_n438_));
  OAI21_X1  g237(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n438_), .A2(new_n430_), .A3(new_n432_), .A4(new_n439_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n424_), .A2(new_n425_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n440_), .A2(KEYINPUT65), .A3(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT8), .ZN(new_n443_));
  AOI21_X1  g242(.A(KEYINPUT65), .B1(new_n440_), .B2(new_n441_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n435_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  AOI211_X1 g244(.A(KEYINPUT65), .B(KEYINPUT8), .C1(new_n440_), .C2(new_n441_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n412_), .B(new_n414_), .C1(new_n445_), .C2(new_n446_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n413_), .A2(KEYINPUT66), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G230gat), .A2(G233gat), .ZN(new_n451_));
  INV_X1    g250(.A(new_n411_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n452_), .B1(new_n409_), .B2(new_n408_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n440_), .A2(new_n441_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT65), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n456_), .A2(KEYINPUT8), .A3(new_n442_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n446_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n453_), .A2(new_n457_), .A3(new_n458_), .A4(new_n435_), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n412_), .B(new_n448_), .C1(new_n445_), .C2(new_n446_), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n450_), .A2(new_n451_), .A3(new_n459_), .A4(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n457_), .A2(new_n458_), .A3(new_n435_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(new_n412_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n459_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n451_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n461_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G120gat), .B(G148gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n469_), .B(KEYINPUT5), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G176gat), .B(G204gat), .ZN(new_n471_));
  XOR2_X1   g270(.A(new_n470_), .B(new_n471_), .Z(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT67), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n468_), .A2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n467_), .A2(KEYINPUT67), .A3(new_n472_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT68), .ZN(new_n477_));
  OR2_X1    g276(.A1(new_n477_), .A2(KEYINPUT13), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(KEYINPUT13), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n476_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n474_), .A2(new_n477_), .A3(KEYINPUT13), .A4(new_n475_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G113gat), .B(G141gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G169gat), .B(G197gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G1gat), .B(G8gat), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G15gat), .B(G22gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT71), .B(G1gat), .ZN(new_n490_));
  INV_X1    g289(.A(G8gat), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT14), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n489_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT72), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT72), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n496_), .B(new_n489_), .C1(new_n492_), .C2(new_n493_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n488_), .B1(new_n495_), .B2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n495_), .A2(new_n497_), .A3(new_n488_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G29gat), .B(G36gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G43gat), .B(G50gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n502_), .B(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n501_), .A2(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n499_), .A2(new_n500_), .A3(new_n504_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G229gat), .A2(G233gat), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n509_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n504_), .B(KEYINPUT15), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n501_), .A2(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n511_), .B1(new_n513_), .B2(new_n507_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n486_), .B1(new_n510_), .B2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(new_n507_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(new_n509_), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n517_), .B(new_n485_), .C1(new_n508_), .C2(new_n509_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n515_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n482_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G232gat), .A2(G233gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT34), .ZN(new_n524_));
  OAI22_X1  g323(.A1(new_n462_), .A2(new_n505_), .B1(KEYINPUT35), .B2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n462_), .A2(new_n512_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT69), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n462_), .A2(new_n512_), .A3(KEYINPUT69), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n525_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n524_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT35), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n530_), .A2(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n533_), .B1(new_n462_), .B2(new_n512_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT70), .ZN(new_n538_));
  NOR3_X1   g337(.A1(new_n537_), .A2(new_n525_), .A3(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n445_), .A2(new_n446_), .ZN(new_n540_));
  AOI22_X1  g339(.A1(new_n540_), .A2(new_n504_), .B1(new_n532_), .B2(new_n531_), .ZN(new_n541_));
  AOI21_X1  g340(.A(KEYINPUT70), .B1(new_n541_), .B2(new_n536_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n539_), .A2(new_n542_), .ZN(new_n543_));
  XOR2_X1   g342(.A(G190gat), .B(G218gat), .Z(new_n544_));
  XNOR2_X1  g343(.A(G134gat), .B(G162gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n547_), .A2(KEYINPUT36), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n535_), .A2(new_n543_), .A3(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n538_), .B1(new_n537_), .B2(new_n525_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n541_), .A2(KEYINPUT70), .A3(new_n536_), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n550_), .B(new_n551_), .C1(new_n530_), .C2(new_n534_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n546_), .B(KEYINPUT36), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n549_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT37), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  XOR2_X1   g356(.A(G127gat), .B(G155gat), .Z(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT16), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G183gat), .B(G211gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT17), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT73), .ZN(new_n564_));
  INV_X1    g363(.A(new_n500_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n564_), .B1(new_n565_), .B2(new_n498_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n499_), .A2(KEYINPUT73), .A3(new_n500_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G231gat), .A2(G233gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n412_), .B(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n566_), .A2(new_n567_), .A3(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n569_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n563_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n453_), .B(new_n568_), .ZN(new_n574_));
  AOI21_X1  g373(.A(KEYINPUT73), .B1(new_n499_), .B2(new_n500_), .ZN(new_n575_));
  NOR3_X1   g374(.A1(new_n565_), .A2(new_n564_), .A3(new_n498_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n574_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n561_), .B(KEYINPUT17), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n577_), .A2(new_n570_), .A3(new_n578_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n573_), .B1(new_n579_), .B2(KEYINPUT74), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(KEYINPUT74), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(KEYINPUT75), .B1(new_n580_), .B2(new_n582_), .ZN(new_n583_));
  OR2_X1    g382(.A1(new_n579_), .A2(KEYINPUT74), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT75), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n584_), .A2(new_n585_), .A3(new_n581_), .A4(new_n573_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n549_), .A2(new_n554_), .A3(KEYINPUT37), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n557_), .A2(new_n583_), .A3(new_n586_), .A4(new_n587_), .ZN(new_n588_));
  NOR3_X1   g387(.A1(new_n404_), .A2(new_n522_), .A3(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(KEYINPUT97), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n589_), .A2(KEYINPUT97), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n202_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n592_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n594_), .A2(KEYINPUT98), .A3(new_n590_), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n377_), .A2(new_n490_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n593_), .A2(new_n595_), .A3(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT38), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n583_), .A2(new_n586_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n555_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NOR3_X1   g401(.A1(new_n404_), .A2(new_n602_), .A3(new_n522_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n377_), .ZN(new_n605_));
  OAI21_X1  g404(.A(G1gat), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n598_), .A2(new_n606_), .ZN(G1324gat));
  INV_X1    g406(.A(new_n403_), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n593_), .A2(new_n595_), .A3(new_n491_), .A4(new_n608_), .ZN(new_n609_));
  NOR4_X1   g408(.A1(new_n404_), .A2(new_n602_), .A3(new_n522_), .A4(new_n403_), .ZN(new_n610_));
  OAI21_X1  g409(.A(KEYINPUT99), .B1(new_n610_), .B2(new_n491_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT39), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n394_), .A2(new_n403_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n383_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n615_), .A2(new_n601_), .A3(new_n521_), .A4(new_n608_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT99), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n616_), .A2(new_n617_), .A3(G8gat), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n611_), .A2(new_n612_), .A3(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n612_), .B1(new_n611_), .B2(new_n618_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT100), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n619_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  AOI211_X1 g421(.A(KEYINPUT100), .B(new_n612_), .C1(new_n611_), .C2(new_n618_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n609_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  XOR2_X1   g423(.A(KEYINPUT101), .B(KEYINPUT40), .Z(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n625_), .ZN(new_n627_));
  OAI211_X1 g426(.A(new_n609_), .B(new_n627_), .C1(new_n622_), .C2(new_n623_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(G1325gat));
  NOR2_X1   g428(.A1(new_n591_), .A2(new_n592_), .ZN(new_n630_));
  INV_X1    g429(.A(G15gat), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n630_), .A2(new_n631_), .A3(new_n384_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n631_), .B1(new_n603_), .B2(new_n384_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n634_), .A2(KEYINPUT41), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(KEYINPUT41), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n632_), .A2(new_n635_), .A3(new_n636_), .ZN(G1326gat));
  XOR2_X1   g436(.A(new_n391_), .B(KEYINPUT102), .Z(new_n638_));
  NOR2_X1   g437(.A1(new_n638_), .A2(G22gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT103), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n630_), .A2(new_n640_), .ZN(new_n641_));
  OAI21_X1  g440(.A(G22gat), .B1(new_n604_), .B2(new_n638_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n642_), .A2(KEYINPUT42), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n642_), .A2(KEYINPUT42), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n641_), .B1(new_n643_), .B2(new_n644_), .ZN(G1327gat));
  NOR2_X1   g444(.A1(new_n404_), .A2(new_n522_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n599_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n647_), .A2(new_n555_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(G29gat), .B1(new_n650_), .B2(new_n377_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n599_), .B1(KEYINPUT105), .B2(KEYINPUT44), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n522_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT43), .ZN(new_n654_));
  INV_X1    g453(.A(new_n587_), .ZN(new_n655_));
  AOI21_X1  g454(.A(KEYINPUT37), .B1(new_n549_), .B2(new_n554_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n654_), .B1(new_n615_), .B2(new_n658_), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n404_), .A2(KEYINPUT43), .A3(new_n657_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n653_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(KEYINPUT105), .B1(KEYINPUT104), .B2(KEYINPUT44), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  OAI211_X1 g463(.A(new_n653_), .B(new_n662_), .C1(new_n659_), .C2(new_n660_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n377_), .A2(G29gat), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n651_), .B1(new_n666_), .B2(new_n667_), .ZN(G1328gat));
  INV_X1    g467(.A(G36gat), .ZN(new_n669_));
  NAND4_X1  g468(.A1(new_n646_), .A2(new_n669_), .A3(new_n608_), .A4(new_n648_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT45), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n403_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n671_), .B1(new_n672_), .B2(new_n669_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT106), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n674_), .A2(KEYINPUT46), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n673_), .B(new_n675_), .ZN(G1329gat));
  AOI21_X1  g475(.A(G43gat), .B1(new_n650_), .B2(new_n384_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT107), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n666_), .A2(G43gat), .A3(new_n384_), .ZN(new_n680_));
  XOR2_X1   g479(.A(KEYINPUT108), .B(KEYINPUT47), .Z(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n679_), .A2(new_n680_), .A3(new_n682_), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n666_), .A2(G43gat), .A3(new_n384_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n681_), .B1(new_n684_), .B2(new_n678_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n683_), .A2(new_n685_), .ZN(G1330gat));
  INV_X1    g485(.A(new_n638_), .ZN(new_n687_));
  AOI21_X1  g486(.A(G50gat), .B1(new_n650_), .B2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n391_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n689_), .A2(G50gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n688_), .B1(new_n666_), .B2(new_n690_), .ZN(G1331gat));
  INV_X1    g490(.A(new_n482_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n404_), .A2(new_n519_), .A3(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(new_n601_), .ZN(new_n694_));
  OAI21_X1  g493(.A(G57gat), .B1(new_n694_), .B2(new_n605_), .ZN(new_n695_));
  NOR4_X1   g494(.A1(new_n404_), .A2(new_n519_), .A3(new_n692_), .A4(new_n588_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n696_), .A2(new_n354_), .A3(new_n377_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(G1332gat));
  INV_X1    g497(.A(G64gat), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n696_), .A2(new_n699_), .A3(new_n608_), .ZN(new_n700_));
  OAI21_X1  g499(.A(G64gat), .B1(new_n694_), .B2(new_n403_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n701_), .A2(KEYINPUT48), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n701_), .A2(KEYINPUT48), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n700_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT109), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n704_), .B(new_n705_), .ZN(G1333gat));
  INV_X1    g505(.A(new_n384_), .ZN(new_n707_));
  OAI21_X1  g506(.A(G71gat), .B1(new_n694_), .B2(new_n707_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT49), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n707_), .A2(G71gat), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT110), .Z(new_n711_));
  NAND2_X1  g510(.A1(new_n696_), .A2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n709_), .A2(new_n712_), .ZN(G1334gat));
  OAI21_X1  g512(.A(G78gat), .B1(new_n694_), .B2(new_n638_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT50), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n638_), .A2(G78gat), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT111), .Z(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(new_n696_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n715_), .A2(new_n718_), .ZN(G1335gat));
  AND2_X1   g518(.A1(new_n693_), .A2(new_n648_), .ZN(new_n720_));
  INV_X1    g519(.A(G85gat), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n720_), .A2(new_n721_), .A3(new_n377_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n659_), .A2(new_n660_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n692_), .A2(new_n519_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(new_n599_), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n723_), .A2(new_n605_), .A3(new_n725_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n722_), .B1(new_n726_), .B2(new_n721_), .ZN(G1336gat));
  AOI21_X1  g526(.A(G92gat), .B1(new_n720_), .B2(new_n608_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT112), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n723_), .A2(new_n725_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n608_), .A2(G92gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n729_), .B1(new_n730_), .B2(new_n731_), .ZN(G1337gat));
  OAI211_X1 g531(.A(new_n720_), .B(new_n384_), .C1(new_n419_), .C2(new_n422_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT113), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n733_), .B(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT51), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n723_), .A2(new_n707_), .A3(new_n725_), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n735_), .B(new_n736_), .C1(new_n437_), .C2(new_n737_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n733_), .B(KEYINPUT113), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n737_), .A2(new_n437_), .ZN(new_n740_));
  OAI21_X1  g539(.A(KEYINPUT51), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n738_), .A2(new_n741_), .ZN(G1338gat));
  NAND3_X1  g541(.A1(new_n720_), .A2(new_n415_), .A3(new_n689_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n725_), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n689_), .B(new_n744_), .C1(new_n659_), .C2(new_n660_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT52), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n745_), .A2(new_n746_), .A3(G106gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n745_), .B2(G106gat), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n743_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g549(.A(new_n472_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n468_), .A2(new_n751_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n519_), .A2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n460_), .A2(new_n459_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n754_), .B1(new_n447_), .B2(new_n449_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT115), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n755_), .A2(new_n756_), .A3(KEYINPUT55), .A4(new_n451_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT55), .ZN(new_n758_));
  OAI21_X1  g557(.A(KEYINPUT115), .B1(new_n461_), .B2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n460_), .A2(new_n459_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n451_), .B1(new_n761_), .B2(new_n450_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n762_), .B1(new_n758_), .B2(new_n461_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n760_), .A2(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(KEYINPUT56), .B1(new_n764_), .B2(new_n472_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT56), .ZN(new_n766_));
  AOI211_X1 g565(.A(new_n766_), .B(new_n751_), .C1(new_n760_), .C2(new_n763_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n753_), .B1(new_n765_), .B2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n508_), .A2(new_n509_), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n769_), .B(new_n485_), .C1(new_n509_), .C2(new_n516_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n476_), .A2(new_n515_), .A3(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n600_), .B1(new_n768_), .B2(new_n771_), .ZN(new_n772_));
  OAI21_X1  g571(.A(KEYINPUT57), .B1(new_n772_), .B2(KEYINPUT116), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT116), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT57), .ZN(new_n775_));
  INV_X1    g574(.A(new_n771_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n761_), .A2(new_n450_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(new_n465_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n461_), .A2(new_n758_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n780_), .B1(new_n759_), .B2(new_n757_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n766_), .B1(new_n781_), .B2(new_n751_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n764_), .A2(KEYINPUT56), .A3(new_n472_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n776_), .B1(new_n784_), .B2(new_n753_), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n774_), .B(new_n775_), .C1(new_n785_), .C2(new_n600_), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n752_), .A2(new_n515_), .A3(new_n770_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n787_), .B1(new_n765_), .B2(new_n767_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT58), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n657_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  OAI211_X1 g589(.A(KEYINPUT58), .B(new_n787_), .C1(new_n765_), .C2(new_n767_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT117), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n784_), .A2(KEYINPUT117), .A3(KEYINPUT58), .A4(new_n787_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n790_), .A2(new_n793_), .A3(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n773_), .A2(new_n786_), .A3(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(new_n599_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n480_), .A2(new_n520_), .A3(new_n481_), .ZN(new_n798_));
  OAI21_X1  g597(.A(KEYINPUT54), .B1(new_n588_), .B2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT114), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT114), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n801_), .B(KEYINPUT54), .C1(new_n588_), .C2(new_n798_), .ZN(new_n802_));
  OR3_X1    g601(.A1(new_n588_), .A2(new_n798_), .A3(KEYINPUT54), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n800_), .A2(new_n802_), .A3(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n797_), .A2(new_n805_), .ZN(new_n806_));
  NOR3_X1   g605(.A1(new_n608_), .A2(new_n605_), .A3(new_n392_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(G113gat), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n809_), .A2(new_n810_), .A3(new_n519_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n809_), .A2(KEYINPUT118), .A3(KEYINPUT59), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT59), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT118), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n813_), .B1(new_n808_), .B2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n520_), .B1(new_n812_), .B2(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n811_), .B1(new_n816_), .B2(new_n810_), .ZN(G1340gat));
  XNOR2_X1  g616(.A(KEYINPUT119), .B(G120gat), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT60), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n819_), .B1(new_n482_), .B2(new_n820_), .ZN(new_n821_));
  OR2_X1    g620(.A1(new_n821_), .A2(KEYINPUT120), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(KEYINPUT120), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n819_), .A2(new_n820_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n809_), .A2(new_n822_), .A3(new_n823_), .A4(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n692_), .B1(new_n812_), .B2(new_n815_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n825_), .B1(new_n826_), .B2(new_n818_), .ZN(G1341gat));
  INV_X1    g626(.A(G127gat), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n809_), .A2(new_n828_), .A3(new_n647_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n599_), .B1(new_n812_), .B2(new_n815_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n829_), .B1(new_n830_), .B2(new_n828_), .ZN(G1342gat));
  AOI21_X1  g630(.A(G134gat), .B1(new_n809_), .B2(new_n600_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n812_), .A2(new_n815_), .ZN(new_n833_));
  XOR2_X1   g632(.A(KEYINPUT121), .B(G134gat), .Z(new_n834_));
  NOR2_X1   g633(.A1(new_n657_), .A2(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n832_), .B1(new_n833_), .B2(new_n835_), .ZN(G1343gat));
  INV_X1    g635(.A(new_n393_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n403_), .A2(new_n377_), .A3(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n838_), .B1(new_n797_), .B2(new_n805_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n519_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g640(.A1(new_n839_), .A2(new_n482_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(G148gat), .ZN(G1345gat));
  XOR2_X1   g642(.A(KEYINPUT61), .B(G155gat), .Z(new_n844_));
  INV_X1    g643(.A(KEYINPUT123), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n839_), .A2(new_n647_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(KEYINPUT122), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT122), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n839_), .A2(new_n848_), .A3(new_n647_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n845_), .B1(new_n847_), .B2(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n848_), .B1(new_n839_), .B2(new_n647_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n804_), .B1(new_n796_), .B2(new_n599_), .ZN(new_n852_));
  NOR4_X1   g651(.A1(new_n852_), .A2(KEYINPUT122), .A3(new_n599_), .A4(new_n838_), .ZN(new_n853_));
  NOR3_X1   g652(.A1(new_n851_), .A2(new_n853_), .A3(KEYINPUT123), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n844_), .B1(new_n850_), .B2(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n847_), .A2(new_n845_), .A3(new_n849_), .ZN(new_n856_));
  OAI21_X1  g655(.A(KEYINPUT123), .B1(new_n851_), .B2(new_n853_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n844_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n856_), .A2(new_n857_), .A3(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n855_), .A2(new_n859_), .ZN(G1346gat));
  INV_X1    g659(.A(new_n839_), .ZN(new_n861_));
  OR3_X1    g660(.A1(new_n861_), .A2(G162gat), .A3(new_n555_), .ZN(new_n862_));
  OAI21_X1  g661(.A(G162gat), .B1(new_n861_), .B2(new_n657_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(G1347gat));
  AOI21_X1  g663(.A(new_n687_), .B1(new_n797_), .B2(new_n805_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n608_), .A2(new_n605_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n866_), .A2(new_n707_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n868_), .A2(new_n520_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n865_), .A2(new_n334_), .A3(new_n869_), .ZN(new_n870_));
  AOI211_X1 g669(.A(KEYINPUT62), .B(new_n225_), .C1(new_n865_), .C2(new_n869_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT62), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n806_), .A2(new_n638_), .A3(new_n869_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n872_), .B1(new_n873_), .B2(G169gat), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n870_), .B1(new_n871_), .B2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(KEYINPUT124), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT124), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n877_), .B(new_n870_), .C1(new_n871_), .C2(new_n874_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n878_), .ZN(G1348gat));
  INV_X1    g678(.A(new_n865_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n880_), .A2(new_n868_), .ZN(new_n881_));
  AOI21_X1  g680(.A(G176gat), .B1(new_n881_), .B2(new_n482_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n852_), .A2(new_n689_), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n868_), .A2(new_n226_), .A3(new_n692_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n882_), .B1(new_n883_), .B2(new_n884_), .ZN(G1349gat));
  INV_X1    g684(.A(new_n332_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n881_), .A2(new_n647_), .A3(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT125), .ZN(new_n888_));
  NOR4_X1   g687(.A1(new_n852_), .A2(new_n599_), .A3(new_n689_), .A4(new_n868_), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n887_), .B(new_n888_), .C1(G183gat), .C2(new_n889_), .ZN(new_n890_));
  NOR4_X1   g689(.A1(new_n880_), .A2(new_n599_), .A3(new_n332_), .A4(new_n868_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n889_), .A2(G183gat), .ZN(new_n892_));
  OAI21_X1  g691(.A(KEYINPUT125), .B1(new_n891_), .B2(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n890_), .A2(new_n893_), .ZN(G1350gat));
  NAND3_X1  g693(.A1(new_n881_), .A2(new_n600_), .A3(new_n234_), .ZN(new_n895_));
  NOR3_X1   g694(.A1(new_n880_), .A2(new_n657_), .A3(new_n868_), .ZN(new_n896_));
  INV_X1    g695(.A(G190gat), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n895_), .B1(new_n896_), .B2(new_n897_), .ZN(G1351gat));
  NOR3_X1   g697(.A1(new_n852_), .A2(new_n393_), .A3(new_n866_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(new_n519_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g700(.A1(new_n899_), .A2(new_n482_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(G204gat), .ZN(G1353gat));
  NOR4_X1   g702(.A1(new_n852_), .A2(new_n599_), .A3(new_n393_), .A4(new_n866_), .ZN(new_n904_));
  XOR2_X1   g703(.A(KEYINPUT63), .B(G211gat), .Z(new_n905_));
  AND3_X1   g704(.A1(new_n904_), .A2(KEYINPUT126), .A3(new_n905_), .ZN(new_n906_));
  NOR3_X1   g705(.A1(new_n904_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n907_));
  AOI21_X1  g706(.A(KEYINPUT126), .B1(new_n904_), .B2(new_n905_), .ZN(new_n908_));
  NOR3_X1   g707(.A1(new_n906_), .A2(new_n907_), .A3(new_n908_), .ZN(G1354gat));
  NAND2_X1  g708(.A1(new_n899_), .A2(new_n600_), .ZN(new_n910_));
  XOR2_X1   g709(.A(KEYINPUT127), .B(G218gat), .Z(new_n911_));
  NOR2_X1   g710(.A1(new_n657_), .A2(new_n911_), .ZN(new_n912_));
  AOI22_X1  g711(.A1(new_n910_), .A2(new_n911_), .B1(new_n899_), .B2(new_n912_), .ZN(G1355gat));
endmodule


