//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 1 0 0 0 1 1 0 0 0 1 0 1 0 0 1 0 0 1 1 0 1 0 0 1 0 0 1 0 1 0 0 1 1 0 1 0 0 0 1 0 0 0 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n694_, new_n695_, new_n696_, new_n698_, new_n699_, new_n700_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n738_, new_n739_, new_n740_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n822_, new_n823_, new_n824_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n836_, new_n837_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n856_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n864_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G134gat), .B(G162gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n204_), .B(KEYINPUT36), .Z(new_n205_));
  XOR2_X1   g004(.A(G85gat), .B(G92gat), .Z(new_n206_));
  NOR3_X1   g005(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT66), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G99gat), .A2(G106gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT6), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n206_), .B1(new_n208_), .B2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n213_), .B(KEYINPUT8), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT64), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G85gat), .A2(G92gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT9), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n215_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n218_), .B1(new_n206_), .B2(new_n217_), .ZN(new_n219_));
  XOR2_X1   g018(.A(KEYINPUT10), .B(G99gat), .Z(new_n220_));
  INV_X1    g019(.A(G106gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n215_), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n219_), .A2(new_n222_), .A3(new_n223_), .A4(new_n210_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT65), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n214_), .A2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G29gat), .B(G36gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G43gat), .B(G50gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(KEYINPUT15), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n227_), .A2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n214_), .A2(new_n226_), .A3(new_n230_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G232gat), .A2(G233gat), .ZN(new_n234_));
  XOR2_X1   g033(.A(new_n234_), .B(KEYINPUT34), .Z(new_n235_));
  XOR2_X1   g034(.A(KEYINPUT69), .B(KEYINPUT35), .Z(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n233_), .A2(new_n237_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n232_), .A2(new_n238_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n235_), .A2(new_n236_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n239_), .A2(new_n241_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n205_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n244_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n204_), .A2(KEYINPUT36), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n246_), .A2(new_n247_), .A3(new_n242_), .ZN(new_n248_));
  AND2_X1   g047(.A1(new_n245_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT37), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n245_), .A2(new_n248_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT37), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n250_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(G1gat), .ZN(new_n256_));
  INV_X1    g055(.A(G8gat), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT14), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT70), .ZN(new_n259_));
  OR2_X1    g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G15gat), .B(G22gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n258_), .A2(new_n259_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n260_), .A2(new_n261_), .A3(new_n262_), .ZN(new_n263_));
  XOR2_X1   g062(.A(G1gat), .B(G8gat), .Z(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  AND2_X1   g064(.A1(G231gat), .A2(G233gat), .ZN(new_n266_));
  XOR2_X1   g065(.A(new_n265_), .B(new_n266_), .Z(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G71gat), .B(G78gat), .ZN(new_n269_));
  XOR2_X1   g068(.A(G57gat), .B(G64gat), .Z(new_n270_));
  INV_X1    g069(.A(KEYINPUT11), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n269_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G57gat), .B(G64gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT11), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n273_), .A2(new_n269_), .A3(KEYINPUT11), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n268_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT17), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G127gat), .B(G155gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT16), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(G183gat), .ZN(new_n282_));
  INV_X1    g081(.A(G211gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  NOR3_X1   g083(.A1(new_n278_), .A2(new_n279_), .A3(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n277_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n285_), .B1(new_n267_), .B2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n284_), .B(KEYINPUT17), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n277_), .B(KEYINPUT67), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n268_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n267_), .A2(new_n289_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n288_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n287_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n255_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT71), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G225gat), .A2(G233gat), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT79), .ZN(new_n300_));
  INV_X1    g099(.A(G134gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(G127gat), .ZN(new_n302_));
  INV_X1    g101(.A(G127gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(G134gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(G120gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(G113gat), .ZN(new_n307_));
  INV_X1    g106(.A(G113gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(G120gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n305_), .A2(new_n310_), .ZN(new_n311_));
  AOI22_X1  g110(.A1(new_n302_), .A2(new_n304_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n300_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n305_), .A2(new_n310_), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n302_), .A2(new_n304_), .A3(new_n307_), .A4(new_n309_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n314_), .A2(new_n315_), .A3(KEYINPUT79), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n313_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(G155gat), .ZN(new_n318_));
  INV_X1    g117(.A(G162gat), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n318_), .A2(new_n319_), .A3(KEYINPUT81), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT81), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n321_), .B1(G155gat), .B2(G162gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G155gat), .A2(G162gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(KEYINPUT1), .ZN(new_n325_));
  OR2_X1    g124(.A1(new_n324_), .A2(KEYINPUT1), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n323_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  XOR2_X1   g126(.A(G141gat), .B(G148gat), .Z(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  AOI22_X1  g128(.A1(new_n320_), .A2(new_n322_), .B1(G155gat), .B2(G162gat), .ZN(new_n330_));
  NOR2_X1   g129(.A1(G141gat), .A2(G148gat), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT82), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT3), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n331_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G141gat), .A2(G148gat), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT2), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n334_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n333_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n330_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n329_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n317_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n314_), .A2(new_n315_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n329_), .A2(new_n341_), .A3(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n299_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(KEYINPUT4), .B1(new_n317_), .B2(new_n342_), .ZN(new_n347_));
  NOR3_X1   g146(.A1(new_n311_), .A2(new_n312_), .A3(new_n300_), .ZN(new_n348_));
  AOI21_X1  g147(.A(KEYINPUT79), .B1(new_n314_), .B2(new_n315_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n340_), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n351_), .A2(new_n334_), .A3(new_n337_), .A4(new_n338_), .ZN(new_n352_));
  AOI22_X1  g151(.A1(new_n352_), .A2(new_n330_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n345_), .B1(new_n350_), .B2(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n347_), .B1(new_n354_), .B2(KEYINPUT4), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n346_), .B1(new_n355_), .B2(new_n299_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G57gat), .B(G85gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G1gat), .B(G29gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n356_), .A2(new_n361_), .ZN(new_n362_));
  AOI22_X1  g161(.A1(new_n316_), .A2(new_n313_), .B1(new_n329_), .B2(new_n341_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n345_), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT4), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n347_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n365_), .A2(new_n299_), .A3(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n346_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n361_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n362_), .A2(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n227_), .A2(KEYINPUT12), .A3(new_n286_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n289_), .A2(new_n226_), .A3(new_n214_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n289_), .B1(new_n226_), .B2(new_n214_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT68), .B(KEYINPUT12), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n373_), .B(new_n374_), .C1(new_n375_), .C2(new_n376_), .ZN(new_n377_));
  AND2_X1   g176(.A1(G230gat), .A2(G233gat), .ZN(new_n378_));
  OR2_X1    g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n374_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n378_), .B1(new_n380_), .B2(new_n375_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n379_), .A2(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G120gat), .B(G148gat), .ZN(new_n383_));
  INV_X1    g182(.A(G204gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT5), .B(G176gat), .ZN(new_n386_));
  XOR2_X1   g185(.A(new_n385_), .B(new_n386_), .Z(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n382_), .A2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n379_), .A2(new_n381_), .A3(new_n387_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT13), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n389_), .A2(KEYINPUT13), .A3(new_n390_), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n230_), .B(KEYINPUT72), .ZN(new_n396_));
  XOR2_X1   g195(.A(new_n396_), .B(new_n265_), .Z(new_n397_));
  NAND2_X1  g196(.A1(G229gat), .A2(G233gat), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n265_), .ZN(new_n401_));
  OR2_X1    g200(.A1(new_n401_), .A2(new_n396_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n231_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n402_), .A2(new_n398_), .A3(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n400_), .A2(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G113gat), .B(G141gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(G169gat), .ZN(new_n407_));
  INV_X1    g206(.A(G197gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT73), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n405_), .B(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n395_), .A2(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(KEYINPUT78), .A2(G183gat), .A3(G190gat), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(KEYINPUT78), .B1(G183gat), .B2(G190gat), .ZN(new_n417_));
  OAI21_X1  g216(.A(KEYINPUT23), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(G183gat), .ZN(new_n419_));
  INV_X1    g218(.A(G190gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G183gat), .A2(G190gat), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT23), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n418_), .A2(new_n421_), .A3(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G169gat), .A2(G176gat), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(KEYINPUT22), .B(G169gat), .ZN(new_n428_));
  INV_X1    g227(.A(G176gat), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n427_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n425_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(G169gat), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n432_), .A2(new_n429_), .A3(KEYINPUT75), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT75), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n434_), .B1(G169gat), .B2(G176gat), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n433_), .A2(new_n435_), .A3(KEYINPUT24), .A4(new_n426_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT76), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n433_), .A2(new_n435_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT24), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT74), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT26), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n442_), .B1(new_n443_), .B2(G190gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(KEYINPUT25), .B(G183gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(KEYINPUT26), .B(G190gat), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n444_), .B(new_n445_), .C1(new_n446_), .C2(new_n442_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n438_), .A2(new_n441_), .A3(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n422_), .A2(KEYINPUT23), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT77), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n422_), .A2(KEYINPUT77), .A3(KEYINPUT23), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n417_), .ZN(new_n454_));
  AOI21_X1  g253(.A(KEYINPUT23), .B1(new_n454_), .B2(new_n415_), .ZN(new_n455_));
  OAI22_X1  g254(.A1(new_n453_), .A2(new_n455_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n431_), .B1(new_n448_), .B2(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(KEYINPUT30), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(KEYINPUT80), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n317_), .B(KEYINPUT31), .ZN(new_n461_));
  AND2_X1   g260(.A1(G227gat), .A2(G233gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G71gat), .B(G99gat), .ZN(new_n464_));
  OR2_X1    g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G15gat), .B(G43gat), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n463_), .A2(new_n464_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n465_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n467_), .B1(new_n465_), .B2(new_n468_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n460_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n471_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n473_), .A2(new_n459_), .A3(new_n469_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n457_), .ZN(new_n476_));
  OAI21_X1  g275(.A(KEYINPUT87), .B1(new_n408_), .B2(G204gat), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT87), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n478_), .A2(new_n384_), .A3(G197gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n408_), .A2(G204gat), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n477_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT21), .ZN(new_n482_));
  INV_X1    g281(.A(G218gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(G211gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n283_), .A2(G218gat), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n482_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n481_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT89), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n481_), .A2(new_n486_), .A3(KEYINPUT89), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n408_), .A2(G204gat), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n384_), .A2(G197gat), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT21), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  AND2_X1   g293(.A1(new_n484_), .A2(new_n485_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(KEYINPUT88), .B(KEYINPUT21), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n494_), .B(new_n495_), .C1(new_n481_), .C2(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(KEYINPUT90), .B1(new_n491_), .B2(new_n497_), .ZN(new_n498_));
  AND3_X1   g297(.A1(new_n481_), .A2(KEYINPUT89), .A3(new_n486_), .ZN(new_n499_));
  AOI21_X1  g298(.A(KEYINPUT89), .B1(new_n481_), .B2(new_n486_), .ZN(new_n500_));
  OAI211_X1 g299(.A(KEYINPUT90), .B(new_n497_), .C1(new_n499_), .C2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n476_), .B1(new_n498_), .B2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT93), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n503_), .A2(new_n504_), .A3(KEYINPUT20), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n497_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT90), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n457_), .B1(new_n508_), .B2(new_n501_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT20), .ZN(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT93), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G226gat), .A2(G233gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT19), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n421_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(new_n430_), .ZN(new_n515_));
  NOR3_X1   g314(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n516_), .B1(new_n446_), .B2(new_n445_), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n517_), .A2(new_n424_), .A3(new_n418_), .A4(new_n436_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n515_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(new_n506_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n505_), .A2(new_n511_), .A3(new_n513_), .A4(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G8gat), .B(G36gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(KEYINPUT18), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(G64gat), .ZN(new_n524_));
  INV_X1    g323(.A(G92gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n513_), .ZN(new_n528_));
  OAI21_X1  g327(.A(KEYINPUT94), .B1(new_n519_), .B2(new_n506_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n506_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT94), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n530_), .A2(new_n531_), .A3(new_n515_), .A4(new_n518_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n529_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n508_), .A2(new_n457_), .A3(new_n501_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(KEYINPUT20), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n528_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n521_), .A2(new_n527_), .A3(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT95), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT95), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n521_), .A2(new_n539_), .A3(new_n527_), .A4(new_n536_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n521_), .A2(new_n536_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(new_n526_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n538_), .A2(new_n540_), .A3(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT27), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT92), .ZN(new_n546_));
  INV_X1    g345(.A(G233gat), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT85), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n548_), .A2(G228gat), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(G228gat), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n547_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  XOR2_X1   g350(.A(new_n551_), .B(KEYINPUT86), .Z(new_n552_));
  XNOR2_X1  g351(.A(new_n506_), .B(KEYINPUT91), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n342_), .A2(KEYINPUT29), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n552_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n554_), .A2(new_n552_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n556_), .A2(new_n508_), .A3(new_n501_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G78gat), .B(G106gat), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n546_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT83), .ZN(new_n561_));
  OR3_X1    g360(.A1(new_n342_), .A2(new_n561_), .A3(KEYINPUT29), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n561_), .B1(new_n342_), .B2(KEYINPUT29), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G22gat), .B(G50gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(KEYINPUT84), .B(KEYINPUT28), .ZN(new_n566_));
  XOR2_X1   g365(.A(new_n565_), .B(new_n566_), .Z(new_n567_));
  XNOR2_X1  g366(.A(new_n564_), .B(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n559_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n555_), .A2(new_n570_), .A3(new_n557_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n570_), .B1(new_n555_), .B2(new_n557_), .ZN(new_n573_));
  OAI22_X1  g372(.A1(new_n560_), .A2(new_n569_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n573_), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n575_), .A2(new_n568_), .A3(new_n546_), .A4(new_n571_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n372_), .B1(new_n574_), .B2(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n544_), .B1(new_n541_), .B2(new_n526_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n505_), .A2(new_n511_), .A3(new_n528_), .A4(new_n520_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT91), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n506_), .B(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n581_), .A2(new_n519_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n513_), .B1(new_n582_), .B2(new_n535_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n579_), .A2(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(KEYINPUT98), .B1(new_n584_), .B2(new_n527_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT98), .ZN(new_n586_));
  AOI211_X1 g385(.A(new_n586_), .B(new_n526_), .C1(new_n579_), .C2(new_n583_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n578_), .B1(new_n585_), .B2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n545_), .A2(new_n577_), .A3(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n574_), .A2(new_n576_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n355_), .A2(new_n299_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n361_), .B1(new_n354_), .B2(new_n298_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(KEYINPUT33), .B1(new_n356_), .B2(new_n361_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT33), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n369_), .A2(new_n595_), .A3(new_n370_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n593_), .B1(new_n594_), .B2(new_n596_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n538_), .A2(new_n597_), .A3(new_n542_), .A4(new_n540_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n584_), .A2(KEYINPUT32), .A3(new_n526_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n526_), .A2(KEYINPUT32), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n541_), .A2(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n599_), .A2(new_n601_), .A3(new_n372_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n590_), .B1(new_n598_), .B2(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n589_), .B1(KEYINPUT97), .B2(new_n603_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n603_), .A2(KEYINPUT97), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n475_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n372_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n472_), .A2(new_n474_), .A3(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n608_), .A2(new_n590_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n545_), .A2(new_n588_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n414_), .B1(new_n606_), .B2(new_n612_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n297_), .A2(new_n256_), .A3(new_n372_), .A4(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT38), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n249_), .B1(new_n606_), .B2(new_n612_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n414_), .A2(new_n294_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  OAI21_X1  g418(.A(G1gat), .B1(new_n619_), .B2(new_n607_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n614_), .A2(new_n615_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n616_), .A2(new_n620_), .A3(new_n621_), .ZN(G1324gat));
  NAND2_X1  g421(.A1(new_n297_), .A2(new_n613_), .ZN(new_n623_));
  NOR3_X1   g422(.A1(new_n623_), .A2(G8gat), .A3(new_n611_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n617_), .A2(new_n618_), .A3(new_n610_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(G8gat), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(KEYINPUT99), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT99), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n625_), .A2(new_n628_), .A3(G8gat), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n627_), .A2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT39), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT39), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n627_), .A2(new_n632_), .A3(new_n629_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n624_), .B1(new_n631_), .B2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n634_), .B(new_n635_), .Z(G1325gat));
  INV_X1    g435(.A(new_n475_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n617_), .A2(new_n618_), .A3(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(G15gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT41), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n623_), .A2(G15gat), .A3(new_n475_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT101), .ZN(G1326gat));
  INV_X1    g442(.A(new_n590_), .ZN(new_n644_));
  OAI21_X1  g443(.A(G22gat), .B1(new_n619_), .B2(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n645_), .B(new_n646_), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n644_), .A2(G22gat), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n647_), .B1(new_n623_), .B2(new_n648_), .ZN(G1327gat));
  NOR2_X1   g448(.A1(new_n414_), .A2(new_n295_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT43), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n606_), .A2(new_n612_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT103), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n254_), .A2(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n250_), .A2(KEYINPUT103), .A3(new_n253_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n651_), .B1(new_n652_), .B2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n254_), .A2(new_n651_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n658_), .B1(new_n606_), .B2(new_n612_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n650_), .B1(new_n657_), .B2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT44), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  OAI211_X1 g461(.A(KEYINPUT44), .B(new_n650_), .C1(new_n657_), .C2(new_n659_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n372_), .A2(G29gat), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n295_), .A2(new_n251_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n613_), .A2(new_n666_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n667_), .A2(new_n607_), .ZN(new_n668_));
  OAI22_X1  g467(.A1(new_n664_), .A2(new_n665_), .B1(G29gat), .B2(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT104), .ZN(G1328gat));
  INV_X1    g469(.A(KEYINPUT107), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT46), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n667_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT45), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n610_), .B(KEYINPUT106), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n676_), .A2(G36gat), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n674_), .A2(new_n675_), .A3(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n677_), .ZN(new_n679_));
  OAI21_X1  g478(.A(KEYINPUT45), .B1(new_n667_), .B2(new_n679_), .ZN(new_n680_));
  AOI22_X1  g479(.A1(new_n678_), .A2(new_n680_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(G36gat), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n662_), .A2(new_n610_), .A3(new_n663_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT105), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n683_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n662_), .A2(KEYINPUT105), .A3(new_n610_), .A4(new_n663_), .ZN(new_n687_));
  AOI211_X1 g486(.A(new_n673_), .B(new_n682_), .C1(new_n686_), .C2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n673_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n684_), .A2(new_n685_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n690_), .A2(G36gat), .A3(new_n687_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n689_), .B1(new_n691_), .B2(new_n681_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n688_), .A2(new_n692_), .ZN(G1329gat));
  NOR3_X1   g492(.A1(new_n667_), .A2(G43gat), .A3(new_n475_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n662_), .A2(new_n637_), .A3(new_n663_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n695_), .B2(G43gat), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g496(.A(G50gat), .B1(new_n674_), .B2(new_n590_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n664_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n590_), .A2(G50gat), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n698_), .B1(new_n699_), .B2(new_n700_), .ZN(G1331gat));
  NAND2_X1  g500(.A1(new_n393_), .A2(new_n394_), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n617_), .A2(new_n295_), .A3(new_n702_), .A4(new_n412_), .ZN(new_n703_));
  INV_X1    g502(.A(G57gat), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n703_), .A2(new_n704_), .A3(new_n607_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n395_), .A2(new_n413_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n652_), .A2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n297_), .A2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n607_), .B1(new_n709_), .B2(KEYINPUT108), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n710_), .B1(KEYINPUT108), .B2(new_n709_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n705_), .B1(new_n711_), .B2(new_n704_), .ZN(G1332gat));
  OAI21_X1  g511(.A(G64gat), .B1(new_n703_), .B2(new_n676_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT48), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n676_), .A2(G64gat), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT109), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n714_), .B1(new_n708_), .B2(new_n716_), .ZN(G1333gat));
  OAI21_X1  g516(.A(G71gat), .B1(new_n703_), .B2(new_n475_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT49), .ZN(new_n719_));
  OR2_X1    g518(.A1(new_n475_), .A2(G71gat), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n719_), .B1(new_n708_), .B2(new_n720_), .ZN(G1334gat));
  OAI21_X1  g520(.A(G78gat), .B1(new_n703_), .B2(new_n644_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n722_), .B(new_n723_), .ZN(new_n724_));
  OR2_X1    g523(.A1(new_n644_), .A2(G78gat), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n724_), .B1(new_n708_), .B2(new_n725_), .ZN(G1335gat));
  NAND2_X1  g525(.A1(new_n707_), .A2(new_n666_), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n727_), .A2(G85gat), .A3(new_n607_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n652_), .A2(new_n656_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(KEYINPUT43), .ZN(new_n730_));
  INV_X1    g529(.A(new_n659_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  AND3_X1   g531(.A1(new_n732_), .A2(new_n294_), .A3(new_n706_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(new_n372_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n728_), .B1(new_n734_), .B2(G85gat), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT111), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n735_), .B(new_n736_), .ZN(G1336gat));
  OAI21_X1  g536(.A(new_n525_), .B1(new_n727_), .B2(new_n611_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT112), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n676_), .A2(new_n525_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n733_), .B2(new_n740_), .ZN(G1337gat));
  INV_X1    g540(.A(new_n220_), .ZN(new_n742_));
  NOR3_X1   g541(.A1(new_n727_), .A2(new_n742_), .A3(new_n475_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n733_), .A2(new_n637_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n744_), .B2(G99gat), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT51), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n745_), .B(new_n746_), .ZN(G1338gat));
  NAND4_X1  g546(.A1(new_n707_), .A2(new_n221_), .A3(new_n590_), .A4(new_n666_), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n732_), .A2(new_n294_), .A3(new_n590_), .A4(new_n706_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT52), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n749_), .A2(new_n750_), .A3(G106gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(new_n749_), .B2(G106gat), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n748_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g553(.A1(new_n702_), .A2(new_n413_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  OAI21_X1  g555(.A(KEYINPUT54), .B1(new_n756_), .B2(new_n296_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT54), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n755_), .A2(new_n758_), .A3(new_n295_), .A4(new_n255_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(KEYINPUT113), .B1(new_n377_), .B2(new_n378_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(KEYINPUT55), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT55), .ZN(new_n764_));
  OAI211_X1 g563(.A(KEYINPUT113), .B(new_n764_), .C1(new_n377_), .C2(new_n378_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n377_), .A2(new_n378_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n763_), .A2(new_n765_), .A3(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(new_n388_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT56), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT115), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n767_), .A2(KEYINPUT56), .A3(new_n388_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n770_), .A2(new_n771_), .A3(new_n772_), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n397_), .A2(new_n398_), .ZN(new_n774_));
  AND3_X1   g573(.A1(new_n402_), .A2(new_n399_), .A3(new_n403_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n410_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n405_), .A2(new_n409_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n390_), .A2(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(KEYINPUT56), .B1(new_n767_), .B2(new_n388_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n779_), .B1(new_n780_), .B2(KEYINPUT115), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n773_), .A2(KEYINPUT58), .A3(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n773_), .A2(new_n781_), .A3(KEYINPUT116), .A4(KEYINPUT58), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(KEYINPUT58), .B1(new_n773_), .B2(new_n781_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n787_), .A2(new_n255_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n788_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n413_), .A2(new_n390_), .ZN(new_n790_));
  AOI22_X1  g589(.A1(new_n762_), .A2(KEYINPUT55), .B1(new_n378_), .B2(new_n377_), .ZN(new_n791_));
  AOI211_X1 g590(.A(new_n769_), .B(new_n387_), .C1(new_n791_), .C2(new_n765_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n790_), .B1(new_n792_), .B2(new_n780_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n391_), .A2(new_n778_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n249_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(KEYINPUT117), .B1(new_n795_), .B2(KEYINPUT114), .ZN(new_n796_));
  OAI21_X1  g595(.A(KEYINPUT57), .B1(new_n795_), .B2(KEYINPUT117), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  OAI211_X1 g597(.A(KEYINPUT117), .B(KEYINPUT57), .C1(new_n795_), .C2(KEYINPUT114), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n789_), .A2(new_n798_), .A3(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n761_), .B1(new_n800_), .B2(new_n294_), .ZN(new_n801_));
  NOR4_X1   g600(.A1(new_n475_), .A2(new_n610_), .A3(new_n590_), .A4(new_n607_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n801_), .A2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT59), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(KEYINPUT59), .B1(new_n801_), .B2(new_n803_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n806_), .A2(new_n413_), .A3(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(G113gat), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n804_), .A2(new_n308_), .A3(new_n413_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(G1340gat));
  NAND3_X1  g610(.A1(new_n806_), .A2(new_n702_), .A3(new_n807_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(G120gat), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n800_), .A2(new_n294_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n760_), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT60), .B1(new_n702_), .B2(new_n306_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n816_), .B1(KEYINPUT60), .B2(new_n306_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n815_), .A2(new_n802_), .A3(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT118), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n818_), .B(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n813_), .A2(new_n820_), .ZN(G1341gat));
  NAND3_X1  g620(.A1(new_n806_), .A2(new_n295_), .A3(new_n807_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(G127gat), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n804_), .A2(new_n303_), .A3(new_n295_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(G1342gat));
  AOI21_X1  g624(.A(G134gat), .B1(new_n804_), .B2(new_n249_), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n806_), .A2(new_n807_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n254_), .A2(G134gat), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n828_), .B(KEYINPUT119), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n826_), .B1(new_n827_), .B2(new_n829_), .ZN(G1343gat));
  INV_X1    g629(.A(new_n676_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n475_), .A2(new_n590_), .A3(new_n372_), .ZN(new_n832_));
  NOR3_X1   g631(.A1(new_n801_), .A2(new_n831_), .A3(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n413_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n702_), .ZN(new_n836_));
  XOR2_X1   g635(.A(KEYINPUT120), .B(G148gat), .Z(new_n837_));
  XNOR2_X1  g636(.A(new_n836_), .B(new_n837_), .ZN(G1345gat));
  NAND2_X1  g637(.A1(new_n833_), .A2(new_n295_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(KEYINPUT61), .B(G155gat), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(KEYINPUT121), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n839_), .B(new_n842_), .ZN(G1346gat));
  AOI21_X1  g642(.A(G162gat), .B1(new_n833_), .B2(new_n249_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n319_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n844_), .B1(new_n833_), .B2(new_n845_), .ZN(G1347gat));
  NOR2_X1   g645(.A1(new_n801_), .A2(new_n676_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n609_), .ZN(new_n848_));
  OAI211_X1 g647(.A(KEYINPUT62), .B(G169gat), .C1(new_n848_), .C2(new_n412_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n609_), .ZN(new_n850_));
  NOR4_X1   g649(.A1(new_n801_), .A2(new_n850_), .A3(new_n412_), .A4(new_n676_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n428_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT62), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n853_), .B1(new_n851_), .B2(new_n432_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n849_), .A2(new_n852_), .A3(new_n854_), .ZN(G1348gat));
  NAND3_X1  g654(.A1(new_n847_), .A2(new_n609_), .A3(new_n702_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(G176gat), .ZN(G1349gat));
  INV_X1    g656(.A(new_n445_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n858_), .B1(KEYINPUT122), .B2(new_n419_), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n847_), .A2(new_n295_), .A3(new_n609_), .A4(new_n859_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n848_), .A2(new_n294_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(KEYINPUT122), .A2(G183gat), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n860_), .B1(new_n861_), .B2(new_n862_), .ZN(G1350gat));
  NAND2_X1  g662(.A1(new_n249_), .A2(new_n446_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(KEYINPUT123), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n815_), .A2(new_n609_), .A3(new_n831_), .A4(new_n865_), .ZN(new_n866_));
  NOR4_X1   g665(.A1(new_n801_), .A2(new_n255_), .A3(new_n850_), .A4(new_n676_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n866_), .B1(new_n867_), .B2(new_n420_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT124), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  OAI211_X1 g669(.A(KEYINPUT124), .B(new_n866_), .C1(new_n867_), .C2(new_n420_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(G1351gat));
  NAND2_X1  g671(.A1(new_n475_), .A2(new_n577_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n847_), .A2(G197gat), .A3(new_n413_), .A4(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT125), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n801_), .A2(new_n676_), .A3(new_n873_), .ZN(new_n878_));
  NAND4_X1  g677(.A1(new_n878_), .A2(KEYINPUT125), .A3(G197gat), .A4(new_n413_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n847_), .A2(new_n413_), .A3(new_n874_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n408_), .ZN(new_n881_));
  AND3_X1   g680(.A1(new_n877_), .A2(new_n879_), .A3(new_n881_), .ZN(G1352gat));
  NAND2_X1  g681(.A1(new_n878_), .A2(new_n702_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(KEYINPUT126), .B(G204gat), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n883_), .B(new_n884_), .ZN(G1353gat));
  INV_X1    g684(.A(new_n878_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT63), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n283_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(KEYINPUT127), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n295_), .B1(new_n887_), .B2(new_n283_), .ZN(new_n890_));
  OR3_X1    g689(.A1(new_n886_), .A2(new_n889_), .A3(new_n890_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n889_), .B1(new_n886_), .B2(new_n890_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(G1354gat));
  OAI21_X1  g692(.A(G218gat), .B1(new_n886_), .B2(new_n255_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n878_), .A2(new_n483_), .A3(new_n249_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1355gat));
endmodule


