//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1 0 0 0 1 1 1 0 1 0 0 0 1 1 0 0 1 0 0 0 1 1 0 0 0 1 1 0 1 1 0 1 1 1 0 1 0 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n584_, new_n586_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n659_, new_n660_,
    new_n661_, new_n663_, new_n664_, new_n665_, new_n667_, new_n668_,
    new_n669_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n799_, new_n800_, new_n802_, new_n803_,
    new_n805_, new_n807_, new_n808_, new_n810_, new_n811_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n848_, new_n849_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n857_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_;
  XOR2_X1   g000(.A(G127gat), .B(G134gat), .Z(new_n202_));
  XOR2_X1   g001(.A(G113gat), .B(G120gat), .Z(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT25), .B(G183gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT26), .B(G190gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT82), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT23), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT23), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(G183gat), .A3(G190gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT24), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT24), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n214_), .B(new_n217_), .C1(new_n215_), .C2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT83), .ZN(new_n221_));
  INV_X1    g020(.A(G169gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT22), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(G176gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT22), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n225_), .A2(KEYINPUT83), .A3(G169gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n223_), .A2(new_n224_), .A3(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(KEYINPUT84), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT85), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n229_), .B1(new_n210_), .B2(KEYINPUT23), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n230_), .B1(new_n214_), .B2(new_n229_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(G183gat), .A2(G190gat), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n218_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  OAI22_X1  g032(.A1(new_n209_), .A2(new_n220_), .B1(new_n228_), .B2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT30), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G15gat), .B(G43gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT86), .ZN(new_n237_));
  INV_X1    g036(.A(G99gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G227gat), .A2(G233gat), .ZN(new_n240_));
  INV_X1    g039(.A(G71gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n239_), .B(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n235_), .A2(new_n243_), .ZN(new_n244_));
  XOR2_X1   g043(.A(new_n244_), .B(KEYINPUT87), .Z(new_n245_));
  INV_X1    g044(.A(KEYINPUT31), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n235_), .A2(new_n243_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT88), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n245_), .A2(new_n246_), .A3(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n246_), .B1(new_n245_), .B2(new_n248_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n205_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n251_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n253_), .A2(new_n204_), .A3(new_n249_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G155gat), .A2(G162gat), .ZN(new_n255_));
  NOR2_X1   g054(.A1(G155gat), .A2(G162gat), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(G141gat), .A2(G148gat), .ZN(new_n258_));
  XOR2_X1   g057(.A(new_n258_), .B(KEYINPUT3), .Z(new_n259_));
  NAND2_X1  g058(.A1(G141gat), .A2(G148gat), .ZN(new_n260_));
  XOR2_X1   g059(.A(new_n260_), .B(KEYINPUT2), .Z(new_n261_));
  OAI211_X1 g060(.A(new_n255_), .B(new_n257_), .C1(new_n259_), .C2(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n256_), .B1(KEYINPUT1), .B2(new_n255_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n263_), .B1(KEYINPUT1), .B2(new_n255_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n258_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n264_), .A2(new_n265_), .A3(new_n260_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n262_), .A2(new_n266_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n267_), .A2(KEYINPUT29), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT28), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G211gat), .B(G218gat), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  XOR2_X1   g070(.A(G197gat), .B(G204gat), .Z(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(KEYINPUT21), .A3(new_n272_), .ZN(new_n273_));
  XOR2_X1   g072(.A(new_n273_), .B(KEYINPUT90), .Z(new_n274_));
  INV_X1    g073(.A(G197gat), .ZN(new_n275_));
  OR3_X1    g074(.A1(new_n275_), .A2(KEYINPUT89), .A3(G204gat), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT89), .ZN(new_n277_));
  OAI211_X1 g076(.A(KEYINPUT21), .B(new_n276_), .C1(new_n272_), .C2(new_n277_), .ZN(new_n278_));
  OAI211_X1 g077(.A(new_n278_), .B(new_n270_), .C1(KEYINPUT21), .C2(new_n272_), .ZN(new_n279_));
  AOI22_X1  g078(.A1(new_n274_), .A2(new_n279_), .B1(KEYINPUT29), .B2(new_n267_), .ZN(new_n280_));
  XOR2_X1   g079(.A(new_n269_), .B(new_n280_), .Z(new_n281_));
  NAND2_X1  g080(.A1(G228gat), .A2(G233gat), .ZN(new_n282_));
  INV_X1    g081(.A(G78gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(G106gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G22gat), .B(G50gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n281_), .B(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n252_), .A2(new_n254_), .A3(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n290_), .B1(new_n252_), .B2(new_n254_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT27), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT20), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT22), .B(G169gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(new_n224_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n214_), .ZN(new_n299_));
  OAI211_X1 g098(.A(new_n218_), .B(new_n298_), .C1(new_n299_), .C2(new_n232_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n231_), .B1(new_n216_), .B2(new_n215_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT92), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n215_), .B1(new_n219_), .B2(KEYINPUT91), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n303_), .B1(KEYINPUT91), .B2(new_n219_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(new_n208_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n300_), .B1(new_n302_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n274_), .A2(new_n279_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  AOI211_X1 g107(.A(new_n296_), .B(new_n308_), .C1(new_n307_), .C2(new_n234_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G226gat), .A2(G233gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT19), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n309_), .A2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G8gat), .B(G36gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT18), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G64gat), .B(G92gat), .ZN(new_n316_));
  XOR2_X1   g115(.A(new_n315_), .B(new_n316_), .Z(new_n317_));
  NAND2_X1  g116(.A1(new_n306_), .A2(new_n307_), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n318_), .B(KEYINPUT20), .C1(new_n307_), .C2(new_n234_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(new_n311_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n313_), .A2(new_n317_), .A3(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n317_), .B1(new_n313_), .B2(new_n320_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n295_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  AOI211_X1 g123(.A(KEYINPUT4), .B(new_n205_), .C1(new_n266_), .C2(new_n262_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n267_), .B(new_n205_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n325_), .B1(new_n326_), .B2(KEYINPUT4), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G225gat), .A2(G233gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT94), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G1gat), .B(G29gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(G85gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT0), .B(G57gat), .ZN(new_n333_));
  XOR2_X1   g132(.A(new_n332_), .B(new_n333_), .Z(new_n334_));
  INV_X1    g133(.A(new_n329_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n326_), .A2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n330_), .A2(new_n334_), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  OR2_X1    g137(.A1(new_n338_), .A2(KEYINPUT99), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n334_), .B1(new_n330_), .B2(new_n336_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n340_), .B1(new_n338_), .B2(KEYINPUT99), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  MUX2_X1   g142(.A(new_n319_), .B(new_n309_), .S(new_n311_), .Z(new_n344_));
  OAI211_X1 g143(.A(KEYINPUT27), .B(new_n321_), .C1(new_n344_), .C2(new_n317_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n324_), .A2(new_n343_), .A3(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT93), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n347_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n323_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n349_), .A2(KEYINPUT93), .A3(new_n321_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT95), .ZN(new_n351_));
  OAI21_X1  g150(.A(KEYINPUT96), .B1(new_n337_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT33), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  AND2_X1   g153(.A1(KEYINPUT96), .A2(KEYINPUT33), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n337_), .B1(new_n351_), .B2(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n326_), .A2(KEYINPUT97), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n357_), .A2(new_n335_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n326_), .A2(KEYINPUT97), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n334_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  OR2_X1    g159(.A1(new_n360_), .A2(KEYINPUT98), .ZN(new_n361_));
  AOI22_X1  g160(.A1(new_n360_), .A2(KEYINPUT98), .B1(new_n335_), .B2(new_n327_), .ZN(new_n362_));
  AOI22_X1  g161(.A1(new_n354_), .A2(new_n356_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n348_), .A2(new_n350_), .A3(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n317_), .A2(KEYINPUT32), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n313_), .A2(new_n320_), .A3(new_n365_), .ZN(new_n366_));
  OAI211_X1 g165(.A(new_n342_), .B(new_n366_), .C1(new_n344_), .C2(new_n365_), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n364_), .A2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n252_), .A2(new_n254_), .A3(new_n289_), .ZN(new_n369_));
  OAI22_X1  g168(.A1(new_n294_), .A2(new_n346_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT80), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G29gat), .B(G36gat), .ZN(new_n372_));
  AND2_X1   g171(.A1(new_n372_), .A2(KEYINPUT73), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n372_), .A2(KEYINPUT73), .ZN(new_n374_));
  XOR2_X1   g173(.A(G43gat), .B(G50gat), .Z(new_n375_));
  OR3_X1    g174(.A1(new_n373_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n375_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT15), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G15gat), .B(G22gat), .ZN(new_n380_));
  INV_X1    g179(.A(G1gat), .ZN(new_n381_));
  INV_X1    g180(.A(G8gat), .ZN(new_n382_));
  OAI21_X1  g181(.A(KEYINPUT14), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n380_), .A2(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G1gat), .B(G8gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n379_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G229gat), .A2(G233gat), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n386_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n389_), .B1(new_n378_), .B2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n387_), .A2(new_n391_), .ZN(new_n392_));
  XOR2_X1   g191(.A(new_n378_), .B(new_n386_), .Z(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(new_n389_), .ZN(new_n394_));
  XOR2_X1   g193(.A(G113gat), .B(G141gat), .Z(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(KEYINPUT79), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G169gat), .B(G197gat), .ZN(new_n397_));
  XOR2_X1   g196(.A(new_n396_), .B(new_n397_), .Z(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n392_), .A2(new_n394_), .A3(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n399_), .B1(new_n392_), .B2(new_n394_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n371_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n402_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n404_), .A2(KEYINPUT80), .A3(new_n400_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(KEYINPUT81), .ZN(new_n407_));
  AND2_X1   g206(.A1(new_n370_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G230gat), .A2(G233gat), .ZN(new_n409_));
  XOR2_X1   g208(.A(new_n409_), .B(KEYINPUT64), .Z(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n241_), .A2(KEYINPUT69), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT69), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(G71gat), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n412_), .A2(new_n414_), .A3(new_n283_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G57gat), .B(G64gat), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n415_), .B1(new_n416_), .B2(KEYINPUT11), .ZN(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT69), .B(G71gat), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n418_), .A2(new_n283_), .ZN(new_n419_));
  OAI21_X1  g218(.A(KEYINPUT70), .B1(new_n417_), .B2(new_n419_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n413_), .A2(G71gat), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n241_), .A2(KEYINPUT69), .ZN(new_n422_));
  OAI21_X1  g221(.A(G78gat), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT11), .ZN(new_n424_));
  INV_X1    g223(.A(G57gat), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n425_), .A2(G64gat), .ZN(new_n426_));
  INV_X1    g225(.A(G64gat), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n427_), .A2(G57gat), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n424_), .B1(new_n426_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT70), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n423_), .A2(new_n429_), .A3(new_n430_), .A4(new_n415_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n427_), .A2(G57gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n425_), .A2(G64gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n434_), .A2(new_n424_), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n420_), .A2(new_n431_), .A3(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n435_), .B1(new_n420_), .B2(new_n431_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  OR2_X1    g237(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n439_), .A2(new_n285_), .A3(new_n440_), .ZN(new_n441_));
  OR2_X1    g240(.A1(new_n441_), .A2(KEYINPUT65), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G99gat), .A2(G106gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(KEYINPUT6), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT6), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n445_), .A2(G99gat), .A3(G106gat), .ZN(new_n446_));
  AOI22_X1  g245(.A1(new_n441_), .A2(KEYINPUT65), .B1(new_n444_), .B2(new_n446_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(G85gat), .A2(G92gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G85gat), .A2(G92gat), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n448_), .B1(new_n450_), .B2(KEYINPUT9), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT9), .ZN(new_n452_));
  AND3_X1   g251(.A1(new_n449_), .A2(KEYINPUT66), .A3(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(KEYINPUT66), .B1(new_n449_), .B2(new_n452_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n451_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n442_), .A2(new_n447_), .A3(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT68), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT7), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n238_), .B(new_n285_), .C1(new_n459_), .C2(KEYINPUT67), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT67), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n461_), .A2(KEYINPUT7), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n458_), .B1(new_n460_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n238_), .A2(new_n285_), .ZN(new_n464_));
  AOI22_X1  g263(.A1(new_n444_), .A2(new_n446_), .B1(new_n464_), .B2(KEYINPUT7), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n459_), .A2(KEYINPUT67), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n461_), .A2(KEYINPUT7), .ZN(new_n467_));
  NOR2_X1   g266(.A1(G99gat), .A2(G106gat), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n466_), .A2(new_n467_), .A3(KEYINPUT68), .A4(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n463_), .A2(new_n465_), .A3(new_n469_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n450_), .A2(new_n448_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT8), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT8), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n470_), .A2(new_n474_), .A3(new_n471_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n457_), .B1(new_n473_), .B2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n411_), .B1(new_n438_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n435_), .ZN(new_n478_));
  AOI22_X1  g277(.A1(new_n424_), .A2(new_n434_), .B1(new_n418_), .B2(new_n283_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n430_), .B1(new_n479_), .B2(new_n423_), .ZN(new_n480_));
  AND4_X1   g279(.A1(new_n430_), .A2(new_n423_), .A3(new_n429_), .A4(new_n415_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n478_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n420_), .A2(new_n431_), .A3(new_n435_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT12), .ZN(new_n485_));
  AND3_X1   g284(.A1(new_n470_), .A2(new_n474_), .A3(new_n471_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n474_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n456_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n484_), .A2(new_n485_), .A3(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n485_), .B1(new_n484_), .B2(new_n488_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n477_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n438_), .A2(new_n476_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n484_), .A2(new_n488_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n411_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n491_), .A2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G120gat), .B(G148gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT5), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G176gat), .B(G204gat), .ZN(new_n498_));
  XOR2_X1   g297(.A(new_n497_), .B(new_n498_), .Z(new_n499_));
  NAND2_X1  g298(.A1(new_n495_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n499_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n491_), .A2(new_n494_), .A3(new_n501_), .ZN(new_n502_));
  AND3_X1   g301(.A1(new_n500_), .A2(KEYINPUT71), .A3(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(KEYINPUT71), .B1(new_n500_), .B2(new_n502_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  OR2_X1    g304(.A1(new_n505_), .A2(KEYINPUT13), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(KEYINPUT13), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G231gat), .A2(G233gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n386_), .B(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n438_), .B(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G127gat), .B(G155gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G183gat), .B(G211gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT17), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  AND2_X1   g319(.A1(new_n518_), .A2(new_n519_), .ZN(new_n521_));
  OR3_X1    g320(.A1(new_n513_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n513_), .A2(new_n520_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G190gat), .B(G218gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT76), .ZN(new_n526_));
  XOR2_X1   g325(.A(G134gat), .B(G162gat), .Z(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT36), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n476_), .A2(new_n378_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G232gat), .A2(G233gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT34), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  XOR2_X1   g332(.A(KEYINPUT72), .B(KEYINPUT35), .Z(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT75), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n530_), .A2(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n537_), .B1(new_n379_), .B2(new_n488_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n533_), .A2(new_n534_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n539_), .B1(new_n537_), .B2(KEYINPUT74), .ZN(new_n540_));
  OR2_X1    g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n528_), .A2(KEYINPUT36), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n538_), .A2(new_n540_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n541_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n542_), .B1(new_n541_), .B2(new_n543_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n529_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT37), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT77), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n548_), .B1(new_n544_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n547_), .A2(new_n551_), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n550_), .B(new_n529_), .C1(new_n545_), .C2(new_n546_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n524_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n408_), .A2(new_n509_), .A3(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n555_), .A2(new_n381_), .A3(new_n342_), .ZN(new_n556_));
  XOR2_X1   g355(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n547_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n524_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n508_), .A2(new_n406_), .ZN(new_n561_));
  AND4_X1   g360(.A1(new_n559_), .A2(new_n370_), .A3(new_n560_), .A4(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT101), .ZN(new_n563_));
  OAI21_X1  g362(.A(G1gat), .B1(new_n563_), .B2(new_n343_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n558_), .A2(new_n564_), .ZN(G1324gat));
  AND2_X1   g364(.A1(new_n324_), .A2(new_n345_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n382_), .B1(new_n562_), .B2(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n568_), .B(KEYINPUT39), .Z(new_n569_));
  NAND3_X1  g368(.A1(new_n555_), .A2(new_n382_), .A3(new_n567_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT40), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n569_), .A2(KEYINPUT40), .A3(new_n570_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(G1325gat));
  INV_X1    g374(.A(new_n252_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n254_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(G15gat), .B1(new_n563_), .B2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT41), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(G15gat), .ZN(new_n582_));
  INV_X1    g381(.A(new_n578_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n555_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n581_), .A2(new_n584_), .ZN(G1326gat));
  OAI21_X1  g384(.A(G22gat), .B1(new_n563_), .B2(new_n289_), .ZN(new_n586_));
  XOR2_X1   g385(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(G22gat), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n555_), .A2(new_n589_), .A3(new_n290_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(new_n590_), .ZN(G1327gat));
  NAND2_X1  g390(.A1(new_n547_), .A2(new_n524_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT104), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n593_), .A2(new_n508_), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n408_), .A2(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(G29gat), .B1(new_n595_), .B2(new_n342_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n552_), .A2(new_n553_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT43), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT103), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n599_), .B1(new_n598_), .B2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n370_), .A2(new_n598_), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n293_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n346_), .B1(new_n604_), .B2(new_n291_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n369_), .B1(new_n364_), .B2(new_n367_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n598_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(new_n601_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n603_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n561_), .A2(new_n524_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  AOI21_X1  g410(.A(KEYINPUT44), .B1(new_n609_), .B2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT44), .ZN(new_n613_));
  AOI211_X1 g412(.A(new_n613_), .B(new_n610_), .C1(new_n603_), .C2(new_n608_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n342_), .A2(G29gat), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n596_), .B1(new_n615_), .B2(new_n616_), .ZN(G1328gat));
  INV_X1    g416(.A(KEYINPUT106), .ZN(new_n618_));
  INV_X1    g417(.A(G36gat), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n408_), .A2(new_n619_), .A3(new_n567_), .A4(new_n594_), .ZN(new_n620_));
  XOR2_X1   g419(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  NOR3_X1   g421(.A1(new_n612_), .A2(new_n614_), .A3(new_n566_), .ZN(new_n623_));
  OAI211_X1 g422(.A(new_n618_), .B(new_n622_), .C1(new_n623_), .C2(new_n619_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT107), .ZN(new_n625_));
  AOI21_X1  g424(.A(KEYINPUT46), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(KEYINPUT106), .B1(new_n625_), .B2(KEYINPUT46), .ZN(new_n627_));
  INV_X1    g426(.A(new_n612_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n614_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n628_), .A2(new_n629_), .A3(new_n567_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(G36gat), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n627_), .B1(new_n631_), .B2(new_n622_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n626_), .A2(new_n632_), .ZN(G1329gat));
  AND2_X1   g432(.A1(new_n583_), .A2(G43gat), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n615_), .A2(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(G43gat), .B1(new_n595_), .B2(new_n583_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT108), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  AOI211_X1 g437(.A(KEYINPUT108), .B(G43gat), .C1(new_n595_), .C2(new_n583_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n635_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g440(.A(G50gat), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n595_), .A2(new_n642_), .A3(new_n290_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT109), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n615_), .A2(new_n290_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n644_), .B1(new_n645_), .B2(G50gat), .ZN(new_n646_));
  AOI211_X1 g445(.A(KEYINPUT109), .B(new_n642_), .C1(new_n615_), .C2(new_n290_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n643_), .B1(new_n646_), .B2(new_n647_), .ZN(G1331gat));
  NOR3_X1   g447(.A1(new_n509_), .A2(new_n524_), .A3(new_n407_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n370_), .A2(new_n559_), .A3(new_n649_), .ZN(new_n650_));
  NOR3_X1   g449(.A1(new_n650_), .A2(new_n425_), .A3(new_n343_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n370_), .A2(new_n406_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n652_), .A2(KEYINPUT110), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n652_), .A2(KEYINPUT110), .ZN(new_n654_));
  OAI211_X1 g453(.A(new_n508_), .B(new_n554_), .C1(new_n653_), .C2(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n343_), .B1(new_n655_), .B2(KEYINPUT111), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n656_), .B1(KEYINPUT111), .B2(new_n655_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n651_), .B1(new_n657_), .B2(new_n425_), .ZN(G1332gat));
  OAI21_X1  g457(.A(G64gat), .B1(new_n650_), .B2(new_n566_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT48), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n567_), .A2(new_n427_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n660_), .B1(new_n655_), .B2(new_n661_), .ZN(G1333gat));
  OAI21_X1  g461(.A(G71gat), .B1(new_n650_), .B2(new_n578_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT49), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n583_), .A2(new_n241_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n664_), .B1(new_n655_), .B2(new_n665_), .ZN(G1334gat));
  OAI21_X1  g465(.A(G78gat), .B1(new_n650_), .B2(new_n289_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT50), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n290_), .A2(new_n283_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n668_), .B1(new_n655_), .B2(new_n669_), .ZN(G1335gat));
  NOR2_X1   g469(.A1(new_n653_), .A2(new_n654_), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n671_), .A2(new_n509_), .A3(new_n593_), .ZN(new_n672_));
  AOI21_X1  g471(.A(G85gat), .B1(new_n672_), .B2(new_n342_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n508_), .A2(new_n524_), .A3(new_n406_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT112), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n675_), .B1(new_n603_), .B2(new_n608_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT113), .Z(new_n677_));
  AND2_X1   g476(.A1(new_n342_), .A2(G85gat), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n673_), .B1(new_n677_), .B2(new_n678_), .ZN(G1336gat));
  AOI21_X1  g478(.A(G92gat), .B1(new_n672_), .B2(new_n567_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n567_), .A2(G92gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n680_), .B1(new_n677_), .B2(new_n681_), .ZN(G1337gat));
  INV_X1    g481(.A(KEYINPUT114), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n583_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n683_), .B1(new_n672_), .B2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n676_), .A2(new_n583_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(G99gat), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n685_), .A2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(KEYINPUT51), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT51), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n685_), .A2(new_n690_), .A3(new_n687_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n691_), .ZN(G1338gat));
  NAND3_X1  g491(.A1(new_n672_), .A2(new_n285_), .A3(new_n290_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT52), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n676_), .A2(new_n290_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n695_), .B2(G106gat), .ZN(new_n696_));
  AOI211_X1 g495(.A(KEYINPUT52), .B(new_n285_), .C1(new_n676_), .C2(new_n290_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n693_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT53), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT53), .ZN(new_n700_));
  OAI211_X1 g499(.A(new_n693_), .B(new_n700_), .C1(new_n696_), .C2(new_n697_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(G1339gat));
  INV_X1    g501(.A(KEYINPUT59), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n567_), .A2(new_n343_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(new_n293_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT119), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT118), .ZN(new_n708_));
  OAI211_X1 g507(.A(KEYINPUT55), .B(new_n477_), .C1(new_n489_), .C2(new_n490_), .ZN(new_n709_));
  OAI21_X1  g508(.A(KEYINPUT12), .B1(new_n438_), .B2(new_n476_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n484_), .A2(new_n488_), .A3(new_n485_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n493_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n709_), .B1(new_n712_), .B2(new_n410_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT55), .ZN(new_n714_));
  AOI21_X1  g513(.A(KEYINPUT115), .B1(new_n491_), .B2(new_n714_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n713_), .A2(new_n715_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n491_), .A2(KEYINPUT115), .A3(new_n714_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n501_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n708_), .B1(new_n718_), .B2(KEYINPUT56), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT115), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n410_), .B1(new_n484_), .B2(new_n488_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n721_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n720_), .B1(new_n722_), .B2(KEYINPUT55), .ZN(new_n723_));
  OAI22_X1  g522(.A1(new_n489_), .A2(new_n490_), .B1(new_n488_), .B2(new_n484_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(new_n411_), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n723_), .A2(new_n717_), .A3(new_n709_), .A4(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n726_), .A2(KEYINPUT56), .A3(new_n499_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(KEYINPUT117), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT117), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n726_), .A2(new_n729_), .A3(KEYINPUT56), .A4(new_n499_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n726_), .A2(new_n499_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT56), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n731_), .A2(KEYINPUT118), .A3(new_n732_), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n719_), .A2(new_n728_), .A3(new_n730_), .A4(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n388_), .B1(new_n378_), .B2(new_n390_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n387_), .A2(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n399_), .B1(new_n393_), .B2(new_n388_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n401_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(new_n502_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(KEYINPUT58), .B1(new_n734_), .B2(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n707_), .B1(new_n741_), .B2(new_n597_), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n728_), .A2(new_n730_), .ZN(new_n743_));
  AOI21_X1  g542(.A(KEYINPUT118), .B1(new_n731_), .B2(new_n732_), .ZN(new_n744_));
  AOI211_X1 g543(.A(new_n708_), .B(KEYINPUT56), .C1(new_n726_), .C2(new_n499_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n739_), .B1(new_n743_), .B2(new_n746_), .ZN(new_n747_));
  OAI211_X1 g546(.A(new_n598_), .B(KEYINPUT119), .C1(new_n747_), .C2(KEYINPUT58), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(KEYINPUT58), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n742_), .A2(new_n748_), .A3(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n502_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n731_), .A2(new_n732_), .ZN(new_n752_));
  AOI211_X1 g551(.A(new_n751_), .B(new_n406_), .C1(new_n752_), .C2(new_n727_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n738_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT116), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  OAI211_X1 g555(.A(KEYINPUT116), .B(new_n738_), .C1(new_n503_), .C2(new_n504_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  OAI211_X1 g557(.A(KEYINPUT57), .B(new_n559_), .C1(new_n753_), .C2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n752_), .A2(new_n727_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n406_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n761_), .A2(new_n762_), .A3(new_n502_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n763_), .A2(new_n757_), .A3(new_n756_), .ZN(new_n764_));
  AOI21_X1  g563(.A(KEYINPUT57), .B1(new_n764_), .B2(new_n559_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n760_), .A2(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n560_), .B1(new_n750_), .B2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n407_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n509_), .A2(new_n768_), .A3(new_n554_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT54), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT54), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n509_), .A2(new_n554_), .A3(new_n771_), .A4(new_n768_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n703_), .B(new_n706_), .C1(new_n767_), .C2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n750_), .A2(new_n766_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n524_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT120), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n777_), .A2(new_n778_), .A3(new_n773_), .ZN(new_n779_));
  OAI21_X1  g578(.A(KEYINPUT120), .B1(new_n767_), .B2(new_n774_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(new_n706_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n775_), .B1(new_n783_), .B2(new_n703_), .ZN(new_n784_));
  OAI21_X1  g583(.A(G113gat), .B1(new_n784_), .B2(new_n768_), .ZN(new_n785_));
  OR2_X1    g584(.A1(new_n406_), .A2(G113gat), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n785_), .B1(new_n782_), .B2(new_n786_), .ZN(G1340gat));
  OAI21_X1  g586(.A(G120gat), .B1(new_n784_), .B2(new_n509_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT60), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n508_), .A2(new_n789_), .ZN(new_n790_));
  MUX2_X1   g589(.A(new_n790_), .B(new_n789_), .S(G120gat), .Z(new_n791_));
  OAI21_X1  g590(.A(new_n788_), .B1(new_n782_), .B2(new_n791_), .ZN(G1341gat));
  NAND2_X1  g591(.A1(new_n560_), .A2(G127gat), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT121), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n775_), .B(new_n794_), .C1(new_n783_), .C2(new_n703_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(G127gat), .B1(new_n783_), .B2(new_n560_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n796_), .A2(new_n797_), .ZN(G1342gat));
  OAI21_X1  g597(.A(G134gat), .B1(new_n784_), .B2(new_n597_), .ZN(new_n799_));
  OR2_X1    g598(.A1(new_n559_), .A2(G134gat), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n799_), .B1(new_n782_), .B2(new_n800_), .ZN(G1343gat));
  NAND3_X1  g600(.A1(new_n781_), .A2(new_n292_), .A3(new_n704_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n802_), .A2(new_n406_), .ZN(new_n803_));
  XOR2_X1   g602(.A(new_n803_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g603(.A1(new_n802_), .A2(new_n509_), .ZN(new_n805_));
  XOR2_X1   g604(.A(new_n805_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g605(.A1(new_n802_), .A2(new_n524_), .ZN(new_n807_));
  XOR2_X1   g606(.A(KEYINPUT61), .B(G155gat), .Z(new_n808_));
  XNOR2_X1  g607(.A(new_n807_), .B(new_n808_), .ZN(G1346gat));
  OAI21_X1  g608(.A(G162gat), .B1(new_n802_), .B2(new_n597_), .ZN(new_n810_));
  OR2_X1    g609(.A1(new_n559_), .A2(G162gat), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n810_), .B1(new_n802_), .B2(new_n811_), .ZN(G1347gat));
  INV_X1    g611(.A(KEYINPUT62), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n290_), .B1(new_n777_), .B2(new_n773_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n566_), .A2(new_n342_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n583_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(KEYINPUT122), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n814_), .A2(new_n817_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n818_), .A2(new_n406_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n813_), .B1(new_n819_), .B2(new_n222_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n297_), .ZN(new_n821_));
  OAI211_X1 g620(.A(KEYINPUT62), .B(G169gat), .C1(new_n818_), .C2(new_n406_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n820_), .A2(new_n821_), .A3(new_n822_), .ZN(G1348gat));
  INV_X1    g622(.A(new_n818_), .ZN(new_n824_));
  AOI21_X1  g623(.A(G176gat), .B1(new_n824_), .B2(new_n508_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n778_), .B1(new_n777_), .B2(new_n773_), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n767_), .A2(KEYINPUT120), .A3(new_n774_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n289_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT123), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT123), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n781_), .A2(new_n830_), .A3(new_n289_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n829_), .A2(new_n831_), .ZN(new_n832_));
  AND3_X1   g631(.A1(new_n817_), .A2(G176gat), .A3(new_n508_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n825_), .B1(new_n832_), .B2(new_n833_), .ZN(G1349gat));
  NAND2_X1  g633(.A1(new_n817_), .A2(new_n560_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n206_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n836_), .A2(new_n814_), .A3(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n835_), .B1(new_n829_), .B2(new_n831_), .ZN(new_n840_));
  AOI21_X1  g639(.A(G183gat), .B1(new_n840_), .B2(KEYINPUT124), .ZN(new_n841_));
  INV_X1    g640(.A(new_n831_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n830_), .B1(new_n781_), .B2(new_n289_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n836_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT124), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n839_), .B1(new_n841_), .B2(new_n846_), .ZN(G1350gat));
  OAI21_X1  g646(.A(G190gat), .B1(new_n818_), .B2(new_n597_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n547_), .A2(new_n207_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n848_), .B1(new_n818_), .B2(new_n849_), .ZN(G1351gat));
  NOR2_X1   g649(.A1(new_n275_), .A2(KEYINPUT125), .ZN(new_n851_));
  AND3_X1   g650(.A1(new_n781_), .A2(new_n292_), .A3(new_n815_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n851_), .B1(new_n852_), .B2(new_n762_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n275_), .A2(KEYINPUT125), .ZN(new_n854_));
  XOR2_X1   g653(.A(new_n854_), .B(KEYINPUT126), .Z(new_n855_));
  XNOR2_X1  g654(.A(new_n853_), .B(new_n855_), .ZN(G1352gat));
  NAND2_X1  g655(.A1(new_n852_), .A2(new_n508_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g657(.A1(new_n852_), .A2(new_n560_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n859_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n860_));
  XOR2_X1   g659(.A(KEYINPUT63), .B(G211gat), .Z(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(new_n859_), .B2(new_n861_), .ZN(G1354gat));
  AOI21_X1  g661(.A(G218gat), .B1(new_n852_), .B2(new_n547_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n598_), .A2(G218gat), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(KEYINPUT127), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n863_), .B1(new_n852_), .B2(new_n865_), .ZN(G1355gat));
endmodule


