//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 0 0 0 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 0 0 0 0 0 1 1 1 1 1 0 1 1 0 0 1 1 0 1 0 1 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n834_, new_n835_, new_n837_, new_n838_, new_n840_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n881_, new_n882_,
    new_n883_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n901_, new_n902_, new_n903_;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G85gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT0), .ZN(new_n204_));
  INV_X1    g003(.A(G57gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XOR2_X1   g005(.A(G127gat), .B(G134gat), .Z(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(G113gat), .ZN(new_n208_));
  XOR2_X1   g007(.A(new_n208_), .B(G120gat), .Z(new_n209_));
  NAND2_X1  g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G141gat), .A2(G148gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n214_), .B(KEYINPUT1), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n213_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT88), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT87), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT83), .ZN(new_n220_));
  INV_X1    g019(.A(G141gat), .ZN(new_n221_));
  INV_X1    g020(.A(G148gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n220_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT83), .B1(G141gat), .B2(G148gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  OR2_X1    g024(.A1(KEYINPUT84), .A2(KEYINPUT3), .ZN(new_n226_));
  NAND2_X1  g025(.A1(KEYINPUT84), .A2(KEYINPUT3), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT86), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT2), .ZN(new_n230_));
  AND3_X1   g029(.A1(new_n210_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n229_), .B1(new_n210_), .B2(new_n230_), .ZN(new_n232_));
  OAI22_X1  g031(.A1(new_n225_), .A2(new_n228_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT85), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  OAI211_X1 g035(.A(KEYINPUT85), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n211_), .A2(KEYINPUT2), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n219_), .B1(new_n233_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n232_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n210_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  AOI22_X1  g043(.A1(new_n236_), .A2(new_n237_), .B1(new_n211_), .B2(KEYINPUT2), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n223_), .A2(new_n224_), .A3(new_n226_), .A4(new_n227_), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n244_), .A2(new_n245_), .A3(KEYINPUT87), .A4(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n241_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n214_), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n249_), .A2(new_n216_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n218_), .B1(new_n248_), .B2(new_n251_), .ZN(new_n252_));
  AOI211_X1 g051(.A(KEYINPUT88), .B(new_n250_), .C1(new_n241_), .C2(new_n247_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n217_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT89), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  OAI211_X1 g055(.A(KEYINPUT89), .B(new_n217_), .C1(new_n252_), .C2(new_n253_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n209_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  AND2_X1   g057(.A1(new_n223_), .A2(new_n224_), .ZN(new_n259_));
  AND2_X1   g058(.A1(new_n226_), .A2(new_n227_), .ZN(new_n260_));
  AOI22_X1  g059(.A1(new_n259_), .A2(new_n260_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n261_));
  AOI21_X1  g060(.A(KEYINPUT87), .B1(new_n261_), .B2(new_n245_), .ZN(new_n262_));
  AND4_X1   g061(.A1(KEYINPUT87), .A2(new_n244_), .A3(new_n245_), .A4(new_n246_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n251_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT88), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n248_), .A2(new_n218_), .A3(new_n251_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n267_), .A2(new_n217_), .A3(new_n209_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT4), .B1(new_n258_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n209_), .ZN(new_n271_));
  AOI21_X1  g070(.A(KEYINPUT89), .B1(new_n267_), .B2(new_n217_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n257_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n271_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n270_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G225gat), .A2(G233gat), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n274_), .A2(new_n278_), .A3(new_n268_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n206_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n278_), .B1(new_n270_), .B2(new_n276_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n281_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n206_), .ZN(new_n285_));
  NOR3_X1   g084(.A1(new_n283_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n282_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G183gat), .A2(G190gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT23), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n290_), .B1(G183gat), .B2(G190gat), .ZN(new_n291_));
  OAI21_X1  g090(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n292_));
  OR3_X1    g091(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n291_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  XOR2_X1   g093(.A(G169gat), .B(G176gat), .Z(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT25), .B(G183gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT26), .B(G190gat), .ZN(new_n297_));
  AOI22_X1  g096(.A1(new_n295_), .A2(KEYINPUT24), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  OR3_X1    g097(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n298_), .A2(new_n290_), .A3(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n294_), .A2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G71gat), .B(G99gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT30), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n301_), .B(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G227gat), .A2(G233gat), .ZN(new_n305_));
  INV_X1    g104(.A(G15gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(G43gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n304_), .B(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT81), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT82), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n209_), .B(KEYINPUT31), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n312_), .B1(new_n309_), .B2(KEYINPUT81), .ZN(new_n313_));
  OR2_X1    g112(.A1(new_n311_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n311_), .A2(new_n313_), .ZN(new_n315_));
  AND2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n288_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(G204gat), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n318_), .A2(G197gat), .ZN(new_n319_));
  INV_X1    g118(.A(G197gat), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n320_), .A2(G204gat), .ZN(new_n321_));
  OAI21_X1  g120(.A(KEYINPUT21), .B1(new_n319_), .B2(new_n321_), .ZN(new_n322_));
  XOR2_X1   g121(.A(G211gat), .B(G218gat), .Z(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT93), .B1(new_n320_), .B2(G204gat), .ZN(new_n325_));
  MUX2_X1   g124(.A(new_n325_), .B(KEYINPUT93), .S(new_n319_), .Z(new_n326_));
  OAI211_X1 g125(.A(new_n322_), .B(new_n324_), .C1(new_n326_), .C2(KEYINPUT21), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n326_), .A2(KEYINPUT21), .A3(new_n323_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n330_), .B1(new_n254_), .B2(KEYINPUT29), .ZN(new_n331_));
  INV_X1    g130(.A(G228gat), .ZN(new_n332_));
  AND2_X1   g131(.A1(new_n332_), .A2(KEYINPUT92), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n332_), .A2(KEYINPUT92), .ZN(new_n334_));
  OAI21_X1  g133(.A(G233gat), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n331_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n256_), .A2(new_n257_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT29), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n329_), .A2(new_n335_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n336_), .B1(new_n338_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT90), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n342_), .B1(new_n337_), .B2(KEYINPUT29), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT29), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n256_), .A2(KEYINPUT90), .A3(new_n344_), .A4(new_n257_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G22gat), .B(G50gat), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n343_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n346_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n341_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n343_), .A2(new_n345_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n346_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n341_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n353_), .A2(new_n354_), .A3(new_n347_), .ZN(new_n355_));
  XOR2_X1   g154(.A(G78gat), .B(G106gat), .Z(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(KEYINPUT91), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT28), .ZN(new_n358_));
  AND3_X1   g157(.A1(new_n350_), .A2(new_n355_), .A3(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n358_), .B1(new_n350_), .B2(new_n355_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n290_), .A2(new_n299_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT94), .ZN(new_n363_));
  XOR2_X1   g162(.A(KEYINPUT22), .B(G169gat), .Z(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT95), .ZN(new_n365_));
  INV_X1    g164(.A(G176gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G169gat), .A2(G176gat), .ZN(new_n368_));
  AND2_X1   g167(.A1(new_n291_), .A2(new_n368_), .ZN(new_n369_));
  AOI22_X1  g168(.A1(new_n363_), .A2(new_n298_), .B1(new_n367_), .B2(new_n369_), .ZN(new_n370_));
  AND2_X1   g169(.A1(new_n370_), .A2(new_n330_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT20), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G226gat), .A2(G233gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT19), .ZN(new_n374_));
  NOR3_X1   g173(.A1(new_n371_), .A2(new_n372_), .A3(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n329_), .A2(new_n301_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT96), .ZN(new_n377_));
  OR2_X1    g176(.A1(new_n301_), .A2(new_n329_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n378_), .B(KEYINPUT20), .C1(new_n330_), .C2(new_n370_), .ZN(new_n379_));
  AOI22_X1  g178(.A1(new_n375_), .A2(new_n377_), .B1(new_n374_), .B2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G8gat), .B(G36gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT18), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(G64gat), .ZN(new_n383_));
  INV_X1    g182(.A(G92gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n380_), .B(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT27), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n380_), .A2(new_n385_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n379_), .A2(new_n374_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT98), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n371_), .B1(new_n391_), .B2(new_n372_), .ZN(new_n392_));
  OAI211_X1 g191(.A(new_n392_), .B(new_n377_), .C1(new_n391_), .C2(new_n372_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n390_), .B1(new_n393_), .B2(new_n374_), .ZN(new_n394_));
  OAI211_X1 g193(.A(KEYINPUT27), .B(new_n389_), .C1(new_n394_), .C2(new_n385_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n388_), .A2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n317_), .A2(new_n361_), .A3(new_n396_), .ZN(new_n397_));
  OAI211_X1 g196(.A(new_n396_), .B(new_n287_), .C1(new_n359_), .C2(new_n360_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(KEYINPUT4), .B1(new_n337_), .B2(new_n271_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n274_), .A2(new_n268_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n400_), .B1(new_n401_), .B2(KEYINPUT4), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n281_), .B(new_n206_), .C1(new_n402_), .C2(new_n278_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT33), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n206_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n274_), .A2(new_n279_), .A3(new_n268_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n386_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n280_), .A2(KEYINPUT33), .A3(new_n281_), .A4(new_n206_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n405_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT97), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n385_), .A2(KEYINPUT32), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n394_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT99), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NOR3_X1   g214(.A1(new_n394_), .A2(KEYINPUT99), .A3(new_n412_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n380_), .A2(new_n412_), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n417_), .B(new_n418_), .C1(new_n282_), .C2(new_n286_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT97), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n405_), .A2(new_n408_), .A3(new_n420_), .A4(new_n409_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n411_), .A2(new_n419_), .A3(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n399_), .B1(new_n422_), .B2(new_n361_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n316_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n397_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G99gat), .A2(G106gat), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT6), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n426_), .B(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT7), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n428_), .B1(KEYINPUT64), .B2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT64), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n431_), .B1(KEYINPUT65), .B2(KEYINPUT7), .ZN(new_n432_));
  INV_X1    g231(.A(G99gat), .ZN(new_n433_));
  INV_X1    g232(.A(G106gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n432_), .B(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n430_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT8), .ZN(new_n438_));
  XOR2_X1   g237(.A(G85gat), .B(G92gat), .Z(new_n439_));
  NAND3_X1  g238(.A1(new_n437_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n438_), .B1(new_n437_), .B2(new_n439_), .ZN(new_n442_));
  INV_X1    g241(.A(G85gat), .ZN(new_n443_));
  NOR3_X1   g242(.A1(new_n443_), .A2(new_n384_), .A3(KEYINPUT9), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n428_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n439_), .A2(KEYINPUT9), .ZN(new_n446_));
  XOR2_X1   g245(.A(KEYINPUT10), .B(G99gat), .Z(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(new_n434_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n445_), .A2(new_n446_), .A3(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n450_), .A2(KEYINPUT69), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT69), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n449_), .A2(new_n452_), .ZN(new_n453_));
  OAI22_X1  g252(.A1(new_n441_), .A2(new_n442_), .B1(new_n451_), .B2(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G57gat), .B(G64gat), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT67), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n455_), .B(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT11), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT68), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n457_), .A2(new_n458_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(KEYINPUT66), .B(G78gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(G71gat), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n460_), .B1(new_n461_), .B2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n461_), .A2(new_n460_), .A3(new_n463_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n459_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n466_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n459_), .ZN(new_n469_));
  NOR3_X1   g268(.A1(new_n468_), .A2(new_n464_), .A3(new_n469_), .ZN(new_n470_));
  OAI211_X1 g269(.A(KEYINPUT12), .B(new_n454_), .C1(new_n467_), .C2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n437_), .A2(new_n439_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT8), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n450_), .B1(new_n473_), .B2(new_n440_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n469_), .B1(new_n468_), .B2(new_n464_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n465_), .A2(new_n466_), .A3(new_n459_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n474_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n471_), .B1(new_n477_), .B2(KEYINPUT12), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n474_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G230gat), .A2(G233gat), .ZN(new_n480_));
  AOI21_X1  g279(.A(KEYINPUT70), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n479_), .A2(KEYINPUT70), .A3(new_n480_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n478_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n479_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n485_), .A2(new_n477_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n486_), .A2(new_n480_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G120gat), .B(G148gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(KEYINPUT5), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(G176gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(new_n318_), .ZN(new_n491_));
  OR3_X1    g290(.A1(new_n484_), .A2(new_n487_), .A3(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n491_), .B1(new_n484_), .B2(new_n487_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT13), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT15), .ZN(new_n497_));
  INV_X1    g296(.A(G50gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G29gat), .B(G36gat), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT71), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(G43gat), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n499_), .B(KEYINPUT71), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n504_), .A2(G43gat), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n498_), .B1(new_n503_), .B2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT72), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n504_), .A2(G43gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n501_), .A2(new_n502_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n508_), .A2(new_n509_), .A3(G50gat), .ZN(new_n510_));
  AND3_X1   g309(.A1(new_n506_), .A2(new_n507_), .A3(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n507_), .B1(new_n506_), .B2(new_n510_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n497_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  XOR2_X1   g312(.A(G1gat), .B(G8gat), .Z(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT74), .ZN(new_n515_));
  INV_X1    g314(.A(G22gat), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n306_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G15gat), .A2(G22gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G1gat), .A2(G8gat), .ZN(new_n519_));
  AOI22_X1  g318(.A1(new_n517_), .A2(new_n518_), .B1(KEYINPUT14), .B2(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n515_), .B(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n510_), .ZN(new_n522_));
  AOI21_X1  g321(.A(G50gat), .B1(new_n508_), .B2(new_n509_), .ZN(new_n523_));
  OAI21_X1  g322(.A(KEYINPUT72), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n506_), .A2(new_n507_), .A3(new_n510_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n524_), .A2(KEYINPUT15), .A3(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n513_), .A2(new_n521_), .A3(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(KEYINPUT79), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G229gat), .A2(G233gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n506_), .A2(new_n510_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT78), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT78), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n530_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n521_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n532_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT79), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n513_), .A2(new_n526_), .A3(new_n537_), .A4(new_n521_), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n528_), .A2(new_n529_), .A3(new_n536_), .A4(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT80), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G113gat), .B(G141gat), .ZN(new_n542_));
  INV_X1    g341(.A(G169gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(new_n320_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n529_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n536_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n535_), .B1(new_n532_), .B2(new_n534_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n547_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n539_), .A2(new_n550_), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n541_), .B(new_n546_), .C1(new_n551_), .C2(new_n540_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n541_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n540_), .B1(new_n539_), .B2(new_n550_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n545_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n552_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n496_), .A2(new_n557_), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n425_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G190gat), .B(G218gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(G134gat), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n561_), .B(G162gat), .Z(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n563_), .A2(KEYINPUT36), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(KEYINPUT36), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n513_), .A2(new_n526_), .A3(new_n454_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G232gat), .A2(G233gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT34), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT35), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n531_), .A2(new_n474_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n567_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n570_), .A2(new_n571_), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n574_), .A2(new_n575_), .ZN(new_n577_));
  OAI211_X1 g376(.A(new_n565_), .B(new_n566_), .C1(new_n576_), .C2(new_n577_), .ZN(new_n578_));
  OR2_X1    g377(.A1(new_n574_), .A2(new_n575_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n574_), .A2(new_n575_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n579_), .A2(new_n564_), .A3(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n578_), .A2(KEYINPUT37), .A3(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT73), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n578_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n579_), .A2(new_n580_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n585_), .A2(KEYINPUT73), .A3(new_n565_), .A4(new_n566_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n584_), .A2(new_n586_), .A3(new_n581_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n582_), .B1(new_n588_), .B2(KEYINPUT37), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n475_), .A2(new_n476_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G231gat), .A2(G233gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(new_n521_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G127gat), .B(G155gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT16), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(G183gat), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n596_), .B(G211gat), .Z(new_n597_));
  XNOR2_X1  g396(.A(KEYINPUT75), .B(KEYINPUT17), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n599_), .B(KEYINPUT76), .Z(new_n600_));
  NAND2_X1  g399(.A1(new_n593_), .A2(new_n600_), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n601_), .A2(KEYINPUT77), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n597_), .B(KEYINPUT17), .Z(new_n603_));
  OR2_X1    g402(.A1(new_n593_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n601_), .A2(KEYINPUT77), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n602_), .A2(new_n604_), .A3(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n589_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n559_), .A2(new_n607_), .ZN(new_n608_));
  OR2_X1    g407(.A1(new_n608_), .A2(KEYINPUT100), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(KEYINPUT100), .ZN(new_n610_));
  AOI211_X1 g409(.A(G1gat), .B(new_n287_), .C1(new_n609_), .C2(new_n610_), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT38), .Z(new_n612_));
  NOR2_X1   g411(.A1(new_n588_), .A2(new_n606_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n559_), .A2(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(G1gat), .B1(new_n614_), .B2(new_n287_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n612_), .A2(new_n615_), .ZN(G1324gat));
  INV_X1    g415(.A(new_n396_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n559_), .A2(new_n617_), .A3(new_n613_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(G8gat), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT39), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n396_), .A2(G8gat), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n623_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n624_));
  OAI21_X1  g423(.A(KEYINPUT101), .B1(new_n621_), .B2(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n619_), .B(KEYINPUT39), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n609_), .A2(new_n610_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(new_n622_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT101), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n626_), .A2(new_n628_), .A3(new_n629_), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n625_), .A2(new_n630_), .A3(KEYINPUT40), .ZN(new_n631_));
  AOI21_X1  g430(.A(KEYINPUT40), .B1(new_n625_), .B2(new_n630_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n631_), .A2(new_n632_), .ZN(G1325gat));
  OAI21_X1  g432(.A(G15gat), .B1(new_n614_), .B2(new_n316_), .ZN(new_n634_));
  XOR2_X1   g433(.A(new_n634_), .B(KEYINPUT41), .Z(new_n635_));
  INV_X1    g434(.A(new_n608_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n636_), .A2(new_n306_), .A3(new_n424_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n637_), .ZN(G1326gat));
  XOR2_X1   g437(.A(new_n361_), .B(KEYINPUT102), .Z(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n636_), .A2(new_n516_), .A3(new_n640_), .ZN(new_n641_));
  OAI21_X1  g440(.A(G22gat), .B1(new_n614_), .B2(new_n639_), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n642_), .B(KEYINPUT103), .Z(new_n643_));
  AND2_X1   g442(.A1(new_n643_), .A2(KEYINPUT42), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n643_), .A2(KEYINPUT42), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n641_), .B1(new_n644_), .B2(new_n645_), .ZN(G1327gat));
  INV_X1    g445(.A(new_n606_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n647_), .A2(new_n587_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n559_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(G29gat), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n649_), .A2(new_n650_), .A3(new_n288_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n425_), .A2(new_n589_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT43), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n425_), .A2(KEYINPUT43), .A3(new_n589_), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n654_), .A2(new_n558_), .A3(new_n606_), .A4(new_n655_), .ZN(new_n656_));
  XOR2_X1   g455(.A(KEYINPUT104), .B(KEYINPUT44), .Z(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT105), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n654_), .A2(new_n655_), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n661_), .A2(KEYINPUT44), .A3(new_n558_), .A4(new_n606_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n656_), .A2(KEYINPUT105), .A3(new_n657_), .ZN(new_n663_));
  AND4_X1   g462(.A1(new_n288_), .A2(new_n660_), .A3(new_n662_), .A4(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n651_), .B1(new_n664_), .B2(new_n650_), .ZN(G1328gat));
  NAND4_X1  g464(.A1(new_n660_), .A2(new_n617_), .A3(new_n662_), .A4(new_n663_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(G36gat), .ZN(new_n667_));
  INV_X1    g466(.A(G36gat), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n649_), .A2(new_n668_), .A3(new_n617_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT45), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n667_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT46), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n667_), .A2(KEYINPUT46), .A3(new_n670_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(G1329gat));
  AND3_X1   g474(.A1(new_n649_), .A2(new_n502_), .A3(new_n424_), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n660_), .A2(new_n424_), .A3(new_n662_), .A4(new_n663_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n676_), .B1(new_n677_), .B2(G43gat), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT47), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  AOI211_X1 g479(.A(KEYINPUT47), .B(new_n676_), .C1(new_n677_), .C2(G43gat), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n680_), .A2(new_n681_), .ZN(G1330gat));
  NOR2_X1   g481(.A1(new_n639_), .A2(G50gat), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT106), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n649_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n361_), .ZN(new_n686_));
  AND4_X1   g485(.A1(new_n686_), .A2(new_n660_), .A3(new_n662_), .A4(new_n663_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n685_), .B1(new_n687_), .B2(new_n498_), .ZN(G1331gat));
  INV_X1    g487(.A(KEYINPUT107), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n425_), .A2(new_n689_), .A3(new_n557_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n689_), .B1(new_n425_), .B2(new_n557_), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n690_), .A2(new_n691_), .A3(new_n495_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n692_), .A2(new_n607_), .ZN(new_n693_));
  AOI21_X1  g492(.A(G57gat), .B1(new_n693_), .B2(new_n288_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n495_), .A2(new_n556_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n425_), .A2(new_n613_), .A3(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT108), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n696_), .B(new_n697_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n287_), .A2(new_n205_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n694_), .B1(new_n698_), .B2(new_n699_), .ZN(G1332gat));
  INV_X1    g499(.A(G64gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n701_), .B1(new_n698_), .B2(new_n617_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT48), .Z(new_n703_));
  NAND3_X1  g502(.A1(new_n693_), .A2(new_n701_), .A3(new_n617_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(G1333gat));
  INV_X1    g504(.A(G71gat), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n693_), .A2(new_n706_), .A3(new_n424_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n698_), .B2(new_n424_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT109), .ZN(new_n709_));
  OR2_X1    g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(new_n709_), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n710_), .A2(KEYINPUT49), .A3(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(KEYINPUT49), .B1(new_n710_), .B2(new_n711_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n707_), .B1(new_n712_), .B2(new_n713_), .ZN(G1334gat));
  INV_X1    g513(.A(G78gat), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n693_), .A2(new_n715_), .A3(new_n640_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT50), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n698_), .A2(new_n640_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n718_), .B2(G78gat), .ZN(new_n719_));
  AOI211_X1 g518(.A(KEYINPUT50), .B(new_n715_), .C1(new_n698_), .C2(new_n640_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n716_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT110), .ZN(G1335gat));
  AOI21_X1  g521(.A(KEYINPUT111), .B1(new_n692_), .B2(new_n648_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n692_), .A2(KEYINPUT111), .A3(new_n648_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(G85gat), .B1(new_n726_), .B2(new_n288_), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n654_), .A2(new_n606_), .A3(new_n655_), .A4(new_n695_), .ZN(new_n728_));
  OR2_X1    g527(.A1(new_n728_), .A2(KEYINPUT112), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(KEYINPUT112), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n287_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n727_), .B1(G85gat), .B2(new_n731_), .ZN(G1336gat));
  AOI21_X1  g531(.A(G92gat), .B1(new_n726_), .B2(new_n617_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n729_), .A2(new_n730_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n617_), .A2(G92gat), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT113), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n733_), .B1(new_n734_), .B2(new_n736_), .ZN(G1337gat));
  NAND2_X1  g536(.A1(new_n424_), .A2(new_n447_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n738_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n728_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n433_), .B1(new_n740_), .B2(new_n424_), .ZN(new_n741_));
  OR3_X1    g540(.A1(new_n739_), .A2(KEYINPUT51), .A3(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(KEYINPUT51), .B1(new_n739_), .B2(new_n741_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(G1338gat));
  INV_X1    g543(.A(new_n725_), .ZN(new_n745_));
  OAI211_X1 g544(.A(new_n434_), .B(new_n686_), .C1(new_n745_), .C2(new_n723_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT52), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n740_), .A2(new_n686_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n748_), .B2(G106gat), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n747_), .B(G106gat), .C1(new_n728_), .C2(new_n361_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n746_), .B1(new_n749_), .B2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT53), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT53), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n746_), .B(new_n754_), .C1(new_n749_), .C2(new_n751_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(G1339gat));
  INV_X1    g555(.A(KEYINPUT114), .ZN(new_n757_));
  OAI21_X1  g556(.A(KEYINPUT55), .B1(new_n484_), .B2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT55), .ZN(new_n759_));
  INV_X1    g558(.A(new_n483_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n760_), .A2(new_n481_), .ZN(new_n761_));
  OAI211_X1 g560(.A(KEYINPUT114), .B(new_n759_), .C1(new_n761_), .C2(new_n478_), .ZN(new_n762_));
  OAI211_X1 g561(.A(G230gat), .B(G233gat), .C1(new_n478_), .C2(new_n485_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n758_), .A2(new_n762_), .A3(new_n763_), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n764_), .A2(KEYINPUT56), .A3(new_n491_), .ZN(new_n765_));
  AOI21_X1  g564(.A(KEYINPUT56), .B1(new_n764_), .B2(new_n491_), .ZN(new_n766_));
  OAI211_X1 g565(.A(new_n556_), .B(new_n492_), .C1(new_n765_), .C2(new_n766_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n528_), .A2(new_n547_), .A3(new_n536_), .A4(new_n538_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n529_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n768_), .A2(new_n545_), .A3(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n553_), .A2(new_n554_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n771_), .B1(new_n772_), .B2(new_n546_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n773_), .A2(KEYINPUT115), .A3(new_n494_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n552_), .A2(new_n494_), .A3(new_n770_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT115), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n767_), .A2(new_n774_), .A3(new_n777_), .ZN(new_n778_));
  AND3_X1   g577(.A1(new_n778_), .A2(KEYINPUT57), .A3(new_n587_), .ZN(new_n779_));
  AOI21_X1  g578(.A(KEYINPUT57), .B1(new_n778_), .B2(new_n587_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n773_), .B(new_n492_), .C1(new_n765_), .C2(new_n766_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT58), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(new_n589_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT116), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n782_), .A2(new_n783_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n784_), .A2(KEYINPUT116), .A3(new_n589_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n787_), .A2(new_n789_), .A3(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n647_), .B1(new_n781_), .B2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n607_), .A2(new_n557_), .A3(new_n495_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT54), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n793_), .B(new_n794_), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n288_), .B(new_n396_), .C1(new_n792_), .C2(new_n795_), .ZN(new_n796_));
  NOR3_X1   g595(.A1(new_n796_), .A2(new_n686_), .A3(new_n316_), .ZN(new_n797_));
  AOI21_X1  g596(.A(G113gat), .B1(new_n797_), .B2(new_n556_), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n784_), .A2(KEYINPUT116), .A3(new_n589_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT116), .B1(new_n784_), .B2(new_n589_), .ZN(new_n800_));
  NOR3_X1   g599(.A1(new_n799_), .A2(new_n800_), .A3(new_n788_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n778_), .A2(new_n587_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT57), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n778_), .A2(KEYINPUT57), .A3(new_n587_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n606_), .B1(new_n801_), .B2(new_n806_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n793_), .B(KEYINPUT54), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n617_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n809_), .A2(new_n288_), .A3(new_n424_), .A4(new_n361_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(KEYINPUT59), .ZN(new_n811_));
  INV_X1    g610(.A(new_n796_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT59), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n812_), .A2(new_n813_), .A3(new_n424_), .A4(new_n361_), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n811_), .A2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n556_), .A2(G113gat), .ZN(new_n816_));
  XOR2_X1   g615(.A(new_n816_), .B(KEYINPUT117), .Z(new_n817_));
  AOI21_X1  g616(.A(new_n798_), .B1(new_n815_), .B2(new_n817_), .ZN(G1340gat));
  NOR2_X1   g617(.A1(new_n495_), .A2(G120gat), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n797_), .B1(KEYINPUT60), .B2(new_n819_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n820_), .A2(new_n496_), .A3(new_n811_), .A4(new_n814_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(G120gat), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n822_), .B1(KEYINPUT60), .B2(new_n820_), .ZN(G1341gat));
  OR2_X1    g622(.A1(KEYINPUT118), .A2(G127gat), .ZN(new_n824_));
  OAI21_X1  g623(.A(G127gat), .B1(new_n606_), .B2(KEYINPUT118), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n811_), .A2(new_n814_), .A3(new_n824_), .A4(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(G127gat), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(new_n810_), .B2(new_n606_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT119), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n826_), .A2(KEYINPUT119), .A3(new_n828_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(G1342gat));
  AOI21_X1  g632(.A(G134gat), .B1(new_n797_), .B2(new_n588_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n589_), .A2(G134gat), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n834_), .B1(new_n815_), .B2(new_n835_), .ZN(G1343gat));
  NOR3_X1   g635(.A1(new_n796_), .A2(new_n424_), .A3(new_n361_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n556_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n496_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g640(.A1(new_n837_), .A2(new_n647_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(KEYINPUT61), .B(G155gat), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n842_), .B(new_n843_), .ZN(G1346gat));
  AOI21_X1  g643(.A(G162gat), .B1(new_n837_), .B2(new_n588_), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n589_), .A2(G162gat), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n845_), .B1(new_n837_), .B2(new_n846_), .ZN(G1347gat));
  AOI21_X1  g646(.A(new_n396_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n848_), .A2(new_n317_), .A3(new_n639_), .ZN(new_n849_));
  OAI21_X1  g648(.A(G169gat), .B1(new_n849_), .B2(new_n557_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT120), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  OAI211_X1 g651(.A(KEYINPUT120), .B(G169gat), .C1(new_n849_), .C2(new_n557_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n852_), .A2(KEYINPUT62), .A3(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT62), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n850_), .A2(new_n851_), .A3(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n849_), .A2(KEYINPUT121), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT121), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n848_), .A2(new_n858_), .A3(new_n317_), .A4(new_n639_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n556_), .A2(new_n365_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(KEYINPUT122), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n854_), .B(new_n856_), .C1(new_n860_), .C2(new_n862_), .ZN(G1348gat));
  OAI211_X1 g662(.A(new_n617_), .B(new_n317_), .C1(new_n792_), .C2(new_n795_), .ZN(new_n864_));
  NOR4_X1   g663(.A1(new_n864_), .A2(new_n366_), .A3(new_n495_), .A4(new_n686_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n857_), .A2(new_n496_), .A3(new_n859_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n366_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(KEYINPUT123), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT123), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n866_), .A2(new_n869_), .A3(new_n366_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n865_), .B1(new_n868_), .B2(new_n870_), .ZN(G1349gat));
  NOR3_X1   g670(.A1(new_n864_), .A2(new_n686_), .A3(new_n606_), .ZN(new_n872_));
  OR2_X1    g671(.A1(new_n872_), .A2(G183gat), .ZN(new_n873_));
  OR2_X1    g672(.A1(new_n606_), .A2(new_n296_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n873_), .B1(new_n860_), .B2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(KEYINPUT124), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT124), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n873_), .B(new_n877_), .C1(new_n860_), .C2(new_n874_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n878_), .ZN(G1350gat));
  NAND3_X1  g678(.A1(new_n857_), .A2(new_n589_), .A3(new_n859_), .ZN(new_n880_));
  AND3_X1   g679(.A1(new_n880_), .A2(KEYINPUT125), .A3(G190gat), .ZN(new_n881_));
  AOI21_X1  g680(.A(KEYINPUT125), .B1(new_n880_), .B2(G190gat), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n588_), .A2(new_n297_), .ZN(new_n883_));
  OAI22_X1  g682(.A1(new_n881_), .A2(new_n882_), .B1(new_n860_), .B2(new_n883_), .ZN(G1351gat));
  NAND2_X1  g683(.A1(new_n848_), .A2(new_n287_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n885_), .A2(new_n424_), .A3(new_n361_), .ZN(new_n886_));
  AOI211_X1 g685(.A(KEYINPUT126), .B(G197gat), .C1(new_n886_), .C2(new_n556_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT126), .ZN(new_n888_));
  INV_X1    g687(.A(new_n885_), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n889_), .A2(new_n556_), .A3(new_n316_), .A4(new_n686_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n888_), .B1(new_n890_), .B2(new_n320_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n890_), .A2(new_n320_), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n887_), .A2(new_n891_), .A3(new_n892_), .ZN(G1352gat));
  NAND2_X1  g692(.A1(new_n886_), .A2(new_n496_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g694(.A1(new_n886_), .A2(new_n647_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(KEYINPUT63), .B(G211gat), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n898_), .B1(new_n896_), .B2(new_n899_), .ZN(G1354gat));
  AOI21_X1  g699(.A(G218gat), .B1(new_n886_), .B2(new_n588_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n589_), .A2(G218gat), .ZN(new_n902_));
  XOR2_X1   g701(.A(new_n902_), .B(KEYINPUT127), .Z(new_n903_));
  AOI21_X1  g702(.A(new_n901_), .B1(new_n886_), .B2(new_n903_), .ZN(G1355gat));
endmodule


