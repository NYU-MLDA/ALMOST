//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 1 1 1 0 0 1 0 0 1 0 0 1 0 0 1 0 0 1 0 0 1 0 1 0 0 0 0 0 0 1 1 0 0 0 1 1 0 1 0 1 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n704_,
    new_n705_, new_n706_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n820_, new_n821_, new_n822_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n838_, new_n840_, new_n841_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n871_, new_n872_, new_n874_, new_n875_, new_n876_,
    new_n878_, new_n879_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n889_, new_n890_;
  XOR2_X1   g000(.A(G1gat), .B(G29gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G57gat), .B(G85gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G225gat), .A2(G233gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT1), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT1), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(G155gat), .A3(G162gat), .ZN(new_n213_));
  OR2_X1    g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT85), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n211_), .A2(new_n213_), .A3(new_n214_), .A4(new_n215_), .ZN(new_n216_));
  OR2_X1    g015(.A1(G141gat), .A2(G148gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G141gat), .A2(G148gat), .ZN(new_n218_));
  AND2_X1   g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n216_), .B(new_n219_), .C1(new_n215_), .C2(new_n213_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT86), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n220_), .B(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n217_), .B(KEYINPUT3), .ZN(new_n223_));
  XOR2_X1   g022(.A(new_n218_), .B(KEYINPUT2), .Z(new_n224_));
  OAI211_X1 g023(.A(new_n210_), .B(new_n214_), .C1(new_n223_), .C2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n222_), .A2(new_n225_), .ZN(new_n226_));
  XOR2_X1   g025(.A(G127gat), .B(G134gat), .Z(new_n227_));
  XOR2_X1   g026(.A(G113gat), .B(G120gat), .Z(new_n228_));
  NOR2_X1   g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n229_), .A2(KEYINPUT84), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(KEYINPUT84), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n227_), .A2(new_n228_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n230_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n226_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT4), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n229_), .ZN(new_n238_));
  AND2_X1   g037(.A1(new_n238_), .A2(new_n232_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n235_), .B1(new_n226_), .B2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n209_), .B(new_n237_), .C1(new_n241_), .C2(new_n236_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n240_), .A2(new_n208_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n207_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT33), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT33), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n237_), .B1(new_n241_), .B2(new_n236_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(new_n208_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n206_), .B1(new_n241_), .B2(new_n209_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n246_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n245_), .B1(new_n250_), .B2(new_n244_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G226gat), .A2(G233gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT19), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G183gat), .A2(G190gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT23), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n256_), .B1(G183gat), .B2(G190gat), .ZN(new_n257_));
  NOR2_X1   g056(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(G169gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT25), .ZN(new_n261_));
  OAI21_X1  g060(.A(KEYINPUT78), .B1(new_n261_), .B2(G183gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT25), .B(G183gat), .ZN(new_n263_));
  OAI211_X1 g062(.A(KEYINPUT79), .B(new_n262_), .C1(new_n263_), .C2(KEYINPUT78), .ZN(new_n264_));
  INV_X1    g063(.A(G183gat), .ZN(new_n265_));
  OR4_X1    g064(.A1(KEYINPUT78), .A2(new_n265_), .A3(KEYINPUT79), .A4(KEYINPUT25), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT26), .B(G190gat), .ZN(new_n268_));
  XOR2_X1   g067(.A(G169gat), .B(G176gat), .Z(new_n269_));
  AOI22_X1  g068(.A1(new_n267_), .A2(new_n268_), .B1(KEYINPUT24), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT80), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n256_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT24), .ZN(new_n274_));
  NOR2_X1   g073(.A1(G169gat), .A2(G176gat), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n273_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n272_), .A2(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n270_), .A2(new_n271_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n260_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G197gat), .B(G204gat), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT21), .ZN(new_n281_));
  OR2_X1    g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G211gat), .B(G218gat), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n282_), .B1(KEYINPUT88), .B2(new_n284_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n285_), .B1(KEYINPUT88), .B2(new_n284_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n280_), .A2(new_n281_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n282_), .A2(new_n287_), .A3(new_n283_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT87), .ZN(new_n289_));
  OR2_X1    g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n288_), .A2(new_n289_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n286_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT20), .B1(new_n279_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT91), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n273_), .B1(new_n268_), .B2(new_n263_), .ZN(new_n295_));
  XOR2_X1   g094(.A(KEYINPUT92), .B(KEYINPUT24), .Z(new_n296_));
  NAND2_X1  g095(.A1(new_n269_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n275_), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n295_), .B(new_n297_), .C1(new_n298_), .C2(new_n296_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT93), .ZN(new_n300_));
  XOR2_X1   g099(.A(new_n260_), .B(KEYINPUT94), .Z(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  AOI22_X1  g101(.A1(new_n293_), .A2(new_n294_), .B1(new_n292_), .B2(new_n302_), .ZN(new_n303_));
  OAI211_X1 g102(.A(KEYINPUT91), .B(KEYINPUT20), .C1(new_n279_), .C2(new_n292_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n254_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  OAI211_X1 g104(.A(KEYINPUT20), .B(new_n254_), .C1(new_n302_), .C2(new_n292_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n279_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n292_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n306_), .A2(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n305_), .A2(new_n310_), .ZN(new_n311_));
  XOR2_X1   g110(.A(G8gat), .B(G36gat), .Z(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G64gat), .B(G92gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n311_), .A2(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n316_), .B1(new_n305_), .B2(new_n310_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n251_), .B1(new_n320_), .B2(KEYINPUT96), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT96), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n318_), .A2(new_n319_), .A3(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n317_), .A2(KEYINPUT32), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NOR3_X1   g124(.A1(new_n305_), .A2(new_n310_), .A3(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT98), .ZN(new_n327_));
  AND3_X1   g126(.A1(new_n242_), .A2(new_n207_), .A3(new_n243_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n328_), .A2(new_n244_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n299_), .A2(new_n260_), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT20), .B1(new_n292_), .B2(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n253_), .B1(new_n309_), .B2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT99), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  OAI211_X1 g133(.A(KEYINPUT99), .B(new_n253_), .C1(new_n309_), .C2(new_n331_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n303_), .A2(new_n304_), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n334_), .B(new_n335_), .C1(new_n336_), .C2(new_n253_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n329_), .B1(new_n337_), .B2(new_n325_), .ZN(new_n338_));
  AOI22_X1  g137(.A1(new_n321_), .A2(new_n323_), .B1(new_n327_), .B2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G227gat), .A2(G233gat), .ZN(new_n340_));
  INV_X1    g139(.A(G71gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(G99gat), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT81), .B(KEYINPUT30), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G15gat), .B(G43gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT82), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n279_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n279_), .A2(new_n348_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n346_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n348_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n307_), .A2(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n354_), .A2(new_n345_), .A3(new_n349_), .ZN(new_n355_));
  OR2_X1    g154(.A1(new_n234_), .A2(KEYINPUT31), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT83), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n234_), .A2(KEYINPUT31), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n356_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n352_), .A2(new_n355_), .A3(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n359_), .B1(new_n352_), .B2(new_n355_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n344_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n362_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n364_), .A2(new_n360_), .A3(new_n343_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n226_), .A2(KEYINPUT29), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G228gat), .A2(G233gat), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n367_), .A2(new_n292_), .A3(new_n368_), .ZN(new_n369_));
  XOR2_X1   g168(.A(KEYINPUT89), .B(KEYINPUT29), .Z(new_n370_));
  AOI21_X1  g169(.A(new_n308_), .B1(new_n226_), .B2(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n369_), .B1(new_n371_), .B2(new_n368_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G78gat), .B(G106gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n373_), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n375_), .B(new_n369_), .C1(new_n371_), .C2(new_n368_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n226_), .A2(KEYINPUT29), .ZN(new_n377_));
  XOR2_X1   g176(.A(G22gat), .B(G50gat), .Z(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT28), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n377_), .B(new_n379_), .ZN(new_n380_));
  AND4_X1   g179(.A1(KEYINPUT90), .A2(new_n374_), .A3(new_n376_), .A4(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT90), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n376_), .A2(new_n382_), .ZN(new_n383_));
  AOI22_X1  g182(.A1(new_n383_), .A2(new_n380_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n381_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n366_), .A2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT100), .B(KEYINPUT27), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n320_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n337_), .A2(new_n316_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n389_), .A2(new_n318_), .A3(KEYINPUT27), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n385_), .A2(new_n363_), .A3(new_n365_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n385_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n329_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  OAI22_X1  g193(.A1(new_n339_), .A2(new_n386_), .B1(new_n391_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT70), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G230gat), .A2(G233gat), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  OAI21_X1  g197(.A(KEYINPUT65), .B1(G85gat), .B2(G92gat), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G85gat), .A2(G92gat), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT64), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n400_), .A2(KEYINPUT9), .A3(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n399_), .B1(new_n402_), .B2(new_n401_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT9), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n406_), .B1(new_n399_), .B2(new_n401_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n404_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(KEYINPUT66), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT66), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n404_), .B(new_n410_), .C1(new_n405_), .C2(new_n407_), .ZN(new_n411_));
  OR2_X1    g210(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n412_));
  INV_X1    g211(.A(G106gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n412_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G99gat), .A2(G106gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT6), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT6), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n418_), .A2(G99gat), .A3(G106gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n415_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n409_), .A2(new_n411_), .A3(new_n422_), .ZN(new_n423_));
  AND2_X1   g222(.A1(G85gat), .A2(G92gat), .ZN(new_n424_));
  NOR2_X1   g223(.A1(G85gat), .A2(G92gat), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n417_), .A2(new_n419_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT7), .ZN(new_n428_));
  INV_X1    g227(.A(G99gat), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n428_), .A2(new_n429_), .A3(new_n413_), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n426_), .B1(new_n427_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT8), .ZN(new_n434_));
  OR2_X1    g233(.A1(new_n424_), .A2(new_n425_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n434_), .B1(new_n435_), .B2(KEYINPUT67), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n433_), .A2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n420_), .A2(new_n431_), .A3(new_n430_), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n438_), .A2(KEYINPUT67), .A3(new_n434_), .A4(new_n426_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n341_), .A2(KEYINPUT68), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT68), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(G71gat), .ZN(new_n443_));
  INV_X1    g242(.A(G78gat), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n441_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n442_), .A2(G71gat), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n341_), .A2(KEYINPUT68), .ZN(new_n447_));
  OAI21_X1  g246(.A(G78gat), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(G64gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(G57gat), .ZN(new_n450_));
  INV_X1    g249(.A(G57gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(G64gat), .ZN(new_n452_));
  AND3_X1   g251(.A1(new_n450_), .A2(new_n452_), .A3(KEYINPUT11), .ZN(new_n453_));
  AOI21_X1  g252(.A(KEYINPUT11), .B1(new_n450_), .B2(new_n452_), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n445_), .B(new_n448_), .C1(new_n453_), .C2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n450_), .A2(new_n452_), .A3(KEYINPUT11), .ZN(new_n456_));
  INV_X1    g255(.A(new_n445_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n444_), .B1(new_n441_), .B2(new_n443_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n456_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n455_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n423_), .A2(new_n440_), .A3(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n460_), .B1(new_n423_), .B2(new_n440_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT69), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n461_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n421_), .B1(new_n408_), .B2(KEYINPUT66), .ZN(new_n465_));
  AOI22_X1  g264(.A1(new_n465_), .A2(new_n411_), .B1(new_n437_), .B2(new_n439_), .ZN(new_n466_));
  NOR3_X1   g265(.A1(new_n466_), .A2(KEYINPUT69), .A3(new_n460_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n398_), .B1(new_n464_), .B2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n462_), .A2(KEYINPUT12), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT12), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n470_), .B1(new_n466_), .B2(new_n460_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n469_), .A2(new_n471_), .A3(new_n397_), .A4(new_n461_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G120gat), .B(G148gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT5), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G176gat), .B(G204gat), .ZN(new_n475_));
  XOR2_X1   g274(.A(new_n474_), .B(new_n475_), .Z(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  AND3_X1   g276(.A1(new_n468_), .A2(new_n472_), .A3(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n477_), .B1(new_n468_), .B2(new_n472_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n396_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n468_), .A2(new_n472_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(new_n476_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n468_), .A2(new_n472_), .A3(new_n477_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n482_), .A2(KEYINPUT70), .A3(new_n483_), .ZN(new_n484_));
  AND3_X1   g283(.A1(new_n480_), .A2(new_n484_), .A3(KEYINPUT13), .ZN(new_n485_));
  AOI21_X1  g284(.A(KEYINPUT13), .B1(new_n480_), .B2(new_n484_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G29gat), .B(G36gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G43gat), .B(G50gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT15), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G15gat), .B(G22gat), .ZN(new_n493_));
  INV_X1    g292(.A(G1gat), .ZN(new_n494_));
  INV_X1    g293(.A(G8gat), .ZN(new_n495_));
  OAI21_X1  g294(.A(KEYINPUT14), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n493_), .B1(new_n496_), .B2(KEYINPUT74), .ZN(new_n497_));
  AND2_X1   g296(.A1(new_n496_), .A2(KEYINPUT74), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G1gat), .B(G8gat), .ZN(new_n499_));
  OR3_X1    g298(.A1(new_n497_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n499_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n492_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G229gat), .A2(G233gat), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n500_), .A2(new_n501_), .A3(new_n491_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n503_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n504_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n505_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n491_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n507_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G113gat), .B(G141gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT76), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G169gat), .B(G197gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n506_), .A2(new_n510_), .A3(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT77), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n515_), .B1(new_n506_), .B2(new_n510_), .ZN(new_n519_));
  OR3_X1    g318(.A1(new_n517_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n518_), .B1(new_n517_), .B2(new_n519_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n488_), .A2(new_n523_), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n395_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n466_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(new_n492_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n466_), .A2(new_n491_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G232gat), .A2(G233gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT34), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT35), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n527_), .A2(new_n528_), .A3(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n531_), .A2(new_n532_), .ZN(new_n535_));
  OR2_X1    g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(new_n535_), .ZN(new_n537_));
  XOR2_X1   g336(.A(G190gat), .B(G218gat), .Z(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT71), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G134gat), .B(G162gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n541_), .A2(KEYINPUT36), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n536_), .A2(new_n537_), .A3(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT72), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n536_), .A2(new_n537_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n541_), .B(KEYINPUT36), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n546_), .A2(new_n548_), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n536_), .A2(KEYINPUT72), .A3(new_n537_), .A4(new_n542_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n545_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(KEYINPUT37), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT73), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n549_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT37), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n546_), .A2(KEYINPUT73), .A3(new_n548_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n554_), .A2(new_n555_), .A3(new_n556_), .A4(new_n543_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n552_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n502_), .B1(G231gat), .B2(G233gat), .ZN(new_n560_));
  NAND2_X1  g359(.A1(G231gat), .A2(G233gat), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n561_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n562_));
  OR3_X1    g361(.A1(new_n560_), .A2(new_n460_), .A3(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n460_), .B1(new_n560_), .B2(new_n562_), .ZN(new_n564_));
  XOR2_X1   g363(.A(G127gat), .B(G155gat), .Z(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT16), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G183gat), .B(G211gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT17), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n563_), .A2(new_n564_), .A3(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n568_), .A2(new_n569_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n573_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n574_));
  OAI21_X1  g373(.A(KEYINPUT75), .B1(new_n572_), .B2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT75), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n563_), .A2(new_n564_), .ZN(new_n577_));
  OAI211_X1 g376(.A(new_n576_), .B(new_n571_), .C1(new_n577_), .C2(new_n573_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n575_), .A2(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n559_), .A2(new_n579_), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n525_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n329_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n581_), .A2(new_n494_), .A3(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT38), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n554_), .A2(new_n556_), .A3(new_n543_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(KEYINPUT102), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT102), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n554_), .A2(new_n587_), .A3(new_n556_), .A4(new_n543_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n586_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n579_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n336_), .A2(new_n253_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n310_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n317_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  NOR3_X1   g394(.A1(new_n305_), .A2(new_n316_), .A3(new_n310_), .ZN(new_n596_));
  OAI21_X1  g395(.A(KEYINPUT96), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n250_), .A2(new_n244_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n597_), .A2(new_n323_), .A3(new_n245_), .A4(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n311_), .A2(KEYINPUT98), .A3(new_n324_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(KEYINPUT98), .B1(new_n311_), .B2(new_n324_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n338_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n386_), .B1(new_n599_), .B2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  OR2_X1    g404(.A1(new_n394_), .A2(new_n391_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n592_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n524_), .A2(KEYINPUT101), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n524_), .A2(KEYINPUT101), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n607_), .A2(new_n610_), .ZN(new_n611_));
  OAI21_X1  g410(.A(G1gat), .B1(new_n611_), .B2(new_n329_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n584_), .A2(new_n612_), .ZN(G1324gat));
  XNOR2_X1  g412(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n607_), .A2(new_n610_), .A3(new_n391_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(G8gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT39), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n581_), .A2(new_n495_), .A3(new_n391_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n614_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n616_), .A2(KEYINPUT39), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT39), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n621_), .B1(new_n615_), .B2(G8gat), .ZN(new_n622_));
  OAI211_X1 g421(.A(new_n618_), .B(new_n614_), .C1(new_n620_), .C2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n619_), .A2(new_n624_), .ZN(G1325gat));
  OAI21_X1  g424(.A(G15gat), .B1(new_n611_), .B2(new_n366_), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n626_), .B(KEYINPUT41), .Z(new_n627_));
  INV_X1    g426(.A(G15gat), .ZN(new_n628_));
  INV_X1    g427(.A(new_n366_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n581_), .A2(new_n628_), .A3(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n627_), .A2(new_n630_), .ZN(G1326gat));
  INV_X1    g430(.A(G22gat), .ZN(new_n632_));
  INV_X1    g431(.A(new_n385_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n581_), .A2(new_n632_), .A3(new_n633_), .ZN(new_n634_));
  OAI21_X1  g433(.A(G22gat), .B1(new_n611_), .B2(new_n385_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n635_), .A2(KEYINPUT42), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n635_), .A2(KEYINPUT42), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n634_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT104), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  OAI211_X1 g439(.A(KEYINPUT104), .B(new_n634_), .C1(new_n636_), .C2(new_n637_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(G1327gat));
  NOR2_X1   g441(.A1(KEYINPUT106), .A2(KEYINPUT44), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n558_), .B(KEYINPUT105), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n394_), .A2(new_n391_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n644_), .B1(new_n645_), .B2(new_n604_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n558_), .A2(KEYINPUT43), .ZN(new_n647_));
  AOI22_X1  g446(.A1(new_n646_), .A2(KEYINPUT43), .B1(new_n395_), .B2(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n591_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n643_), .B1(new_n648_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n643_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT43), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n653_), .B1(new_n395_), .B2(new_n644_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n647_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n655_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n649_), .B(new_n652_), .C1(new_n654_), .C2(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n651_), .A2(new_n582_), .A3(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(G29gat), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n590_), .A2(new_n591_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n525_), .A2(new_n660_), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n329_), .A2(G29gat), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n659_), .B1(new_n661_), .B2(new_n662_), .ZN(G1328gat));
  NAND3_X1  g462(.A1(new_n651_), .A2(new_n391_), .A3(new_n657_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(G36gat), .ZN(new_n665_));
  INV_X1    g464(.A(G36gat), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n525_), .A2(new_n666_), .A3(new_n391_), .A4(new_n660_), .ZN(new_n667_));
  XOR2_X1   g466(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n668_));
  XNOR2_X1  g467(.A(new_n667_), .B(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n665_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT46), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n665_), .A2(new_n669_), .A3(KEYINPUT46), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1329gat));
  NAND4_X1  g473(.A1(new_n651_), .A2(new_n657_), .A3(G43gat), .A4(new_n629_), .ZN(new_n675_));
  INV_X1    g474(.A(G43gat), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n676_), .B1(new_n661_), .B2(new_n366_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n678_), .B(new_n679_), .ZN(G1330gat));
  OR3_X1    g479(.A1(new_n661_), .A2(G50gat), .A3(new_n385_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n651_), .A2(new_n633_), .A3(new_n657_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT109), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(G50gat), .B1(new_n682_), .B2(new_n683_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n681_), .B1(new_n684_), .B2(new_n685_), .ZN(G1331gat));
  NOR2_X1   g485(.A1(new_n487_), .A2(new_n522_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n395_), .A2(new_n687_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n688_), .A2(new_n580_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n689_), .A2(new_n451_), .A3(new_n582_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n607_), .A2(new_n687_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n691_), .A2(new_n582_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n690_), .B1(new_n692_), .B2(new_n451_), .ZN(G1332gat));
  AOI21_X1  g492(.A(new_n449_), .B1(new_n691_), .B2(new_n391_), .ZN(new_n694_));
  XOR2_X1   g493(.A(new_n694_), .B(KEYINPUT48), .Z(new_n695_));
  NAND2_X1  g494(.A1(new_n391_), .A2(new_n449_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT110), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n689_), .A2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n695_), .A2(new_n698_), .ZN(G1333gat));
  AOI21_X1  g498(.A(new_n341_), .B1(new_n691_), .B2(new_n629_), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT49), .Z(new_n701_));
  NAND3_X1  g500(.A1(new_n689_), .A2(new_n341_), .A3(new_n629_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(G1334gat));
  AOI21_X1  g502(.A(new_n444_), .B1(new_n691_), .B2(new_n633_), .ZN(new_n704_));
  XOR2_X1   g503(.A(new_n704_), .B(KEYINPUT50), .Z(new_n705_));
  NAND3_X1  g504(.A1(new_n689_), .A2(new_n444_), .A3(new_n633_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(G1335gat));
  NOR3_X1   g506(.A1(new_n487_), .A2(new_n522_), .A3(new_n591_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n708_), .B1(new_n654_), .B2(new_n656_), .ZN(new_n709_));
  OAI21_X1  g508(.A(G85gat), .B1(new_n709_), .B2(new_n329_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n688_), .A2(new_n660_), .ZN(new_n711_));
  INV_X1    g510(.A(G85gat), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n711_), .A2(new_n712_), .A3(new_n582_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n710_), .A2(new_n713_), .ZN(G1336gat));
  INV_X1    g513(.A(G92gat), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n711_), .A2(new_n715_), .A3(new_n391_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n709_), .B1(new_n388_), .B2(new_n390_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n716_), .B1(new_n717_), .B2(new_n715_), .ZN(G1337gat));
  NAND4_X1  g517(.A1(new_n711_), .A2(new_n412_), .A3(new_n414_), .A4(new_n629_), .ZN(new_n719_));
  OAI21_X1  g518(.A(G99gat), .B1(new_n709_), .B2(new_n366_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g521(.A1(new_n711_), .A2(new_n413_), .A3(new_n633_), .ZN(new_n723_));
  OAI211_X1 g522(.A(new_n633_), .B(new_n708_), .C1(new_n654_), .C2(new_n656_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT52), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n724_), .A2(new_n725_), .A3(G106gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n724_), .B2(G106gat), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n723_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(KEYINPUT53), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT53), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n730_), .B(new_n723_), .C1(new_n726_), .C2(new_n727_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(G1339gat));
  NAND3_X1  g531(.A1(new_n503_), .A2(new_n507_), .A3(new_n505_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n504_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n733_), .A2(new_n514_), .A3(new_n734_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n516_), .A2(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(KEYINPUT115), .B1(new_n736_), .B2(new_n483_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n736_), .A2(new_n483_), .A3(KEYINPUT115), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n461_), .B1(new_n462_), .B2(KEYINPUT12), .ZN(new_n741_));
  NOR3_X1   g540(.A1(new_n466_), .A2(new_n470_), .A3(new_n460_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n398_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(KEYINPUT55), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(new_n472_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT55), .ZN(new_n746_));
  NOR4_X1   g545(.A1(new_n741_), .A2(new_n742_), .A3(new_n746_), .A4(new_n398_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n477_), .B1(new_n745_), .B2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT56), .ZN(new_n750_));
  NOR3_X1   g549(.A1(new_n741_), .A2(new_n742_), .A3(new_n398_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(KEYINPUT55), .B2(new_n743_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n476_), .B1(new_n752_), .B2(new_n747_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT56), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n740_), .B1(new_n750_), .B2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT116), .ZN(new_n757_));
  OAI21_X1  g556(.A(KEYINPUT58), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n750_), .A2(new_n755_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n738_), .A2(new_n739_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT58), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n761_), .A2(KEYINPUT116), .A3(new_n762_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n758_), .A2(new_n763_), .A3(new_n559_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT114), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n765_), .B1(new_n749_), .B2(KEYINPUT56), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n754_), .B1(new_n749_), .B2(KEYINPUT113), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT113), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n753_), .A2(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n766_), .B1(new_n767_), .B2(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(KEYINPUT56), .B1(new_n753_), .B2(new_n768_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n749_), .A2(KEYINPUT113), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n771_), .A2(new_n765_), .A3(new_n772_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n523_), .A2(new_n478_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n770_), .A2(new_n773_), .A3(new_n774_), .ZN(new_n775_));
  NOR3_X1   g574(.A1(new_n478_), .A2(new_n479_), .A3(new_n396_), .ZN(new_n776_));
  AOI21_X1  g575(.A(KEYINPUT70), .B1(new_n482_), .B2(new_n483_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n736_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n589_), .B1(new_n775_), .B2(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n764_), .B1(new_n779_), .B2(KEYINPUT57), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT57), .ZN(new_n781_));
  AOI211_X1 g580(.A(new_n781_), .B(new_n589_), .C1(new_n775_), .C2(new_n778_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n579_), .B1(new_n780_), .B2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT111), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n579_), .A2(new_n522_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n784_), .B1(new_n487_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT13), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n787_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n480_), .A2(new_n484_), .A3(KEYINPUT13), .ZN(new_n789_));
  AND4_X1   g588(.A1(new_n784_), .A2(new_n785_), .A3(new_n788_), .A4(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n558_), .B1(new_n786_), .B2(new_n790_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n791_), .B(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n783_), .A2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n388_), .A2(new_n392_), .A3(new_n390_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT59), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n798_), .A2(KEYINPUT117), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  AND4_X1   g599(.A1(new_n582_), .A2(new_n795_), .A3(new_n797_), .A4(new_n800_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(KEYINPUT117), .B(KEYINPUT59), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n329_), .B1(new_n783_), .B2(new_n794_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n802_), .B1(new_n803_), .B2(new_n797_), .ZN(new_n804_));
  OAI21_X1  g603(.A(KEYINPUT118), .B1(new_n801_), .B2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n803_), .A2(new_n797_), .A3(new_n800_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT118), .ZN(new_n807_));
  AOI211_X1 g606(.A(new_n329_), .B(new_n796_), .C1(new_n783_), .C2(new_n794_), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n806_), .B(new_n807_), .C1(new_n808_), .C2(new_n802_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n805_), .A2(new_n522_), .A3(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(G113gat), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n803_), .A2(new_n797_), .ZN(new_n812_));
  OR3_X1    g611(.A1(new_n812_), .A2(G113gat), .A3(new_n523_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n811_), .A2(new_n813_), .ZN(G1340gat));
  INV_X1    g613(.A(G120gat), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n815_), .B1(new_n487_), .B2(KEYINPUT60), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n808_), .B(new_n816_), .C1(KEYINPUT60), .C2(new_n815_), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n801_), .A2(new_n804_), .A3(new_n487_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n817_), .B1(new_n818_), .B2(new_n815_), .ZN(G1341gat));
  NAND3_X1  g618(.A1(new_n805_), .A2(new_n591_), .A3(new_n809_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(G127gat), .ZN(new_n821_));
  OR3_X1    g620(.A1(new_n812_), .A2(G127gat), .A3(new_n579_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(G1342gat));
  AND2_X1   g622(.A1(new_n805_), .A2(new_n809_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n559_), .A2(G134gat), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n825_), .B(KEYINPUT120), .ZN(new_n826_));
  INV_X1    g625(.A(G134gat), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(new_n812_), .B2(new_n590_), .ZN(new_n828_));
  OR2_X1    g627(.A1(new_n828_), .A2(KEYINPUT119), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(KEYINPUT119), .ZN(new_n830_));
  AOI22_X1  g629(.A1(new_n824_), .A2(new_n826_), .B1(new_n829_), .B2(new_n830_), .ZN(G1343gat));
  NOR3_X1   g630(.A1(new_n391_), .A2(new_n385_), .A3(new_n629_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n795_), .A2(new_n582_), .A3(new_n832_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n833_), .A2(KEYINPUT121), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n833_), .A2(KEYINPUT121), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n522_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n836_), .B(G141gat), .ZN(G1344gat));
  OAI21_X1  g636(.A(new_n488_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(G148gat), .ZN(G1345gat));
  OAI21_X1  g638(.A(new_n591_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(KEYINPUT61), .B(G155gat), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n840_), .B(new_n841_), .ZN(G1346gat));
  OR2_X1    g641(.A1(new_n834_), .A2(new_n835_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n644_), .A2(G162gat), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n589_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n845_));
  INV_X1    g644(.A(G162gat), .ZN(new_n846_));
  AOI22_X1  g645(.A1(new_n843_), .A2(new_n844_), .B1(new_n845_), .B2(new_n846_), .ZN(G1347gat));
  AOI21_X1  g646(.A(new_n582_), .B1(new_n388_), .B2(new_n390_), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n795_), .A2(new_n522_), .A3(new_n392_), .A4(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT62), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n849_), .A2(new_n850_), .A3(G169gat), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT122), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n851_), .A2(new_n852_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n849_), .A2(G169gat), .ZN(new_n855_));
  AOI21_X1  g654(.A(KEYINPUT123), .B1(new_n855_), .B2(KEYINPUT62), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT123), .ZN(new_n857_));
  AOI211_X1 g656(.A(new_n857_), .B(new_n850_), .C1(new_n849_), .C2(G169gat), .ZN(new_n858_));
  OAI22_X1  g657(.A1(new_n853_), .A2(new_n854_), .B1(new_n856_), .B2(new_n858_), .ZN(new_n859_));
  AND3_X1   g658(.A1(new_n795_), .A2(new_n392_), .A3(new_n848_), .ZN(new_n860_));
  XOR2_X1   g659(.A(KEYINPUT22), .B(G169gat), .Z(new_n861_));
  NOR2_X1   g660(.A1(new_n523_), .A2(new_n861_), .ZN(new_n862_));
  XOR2_X1   g661(.A(new_n862_), .B(KEYINPUT124), .Z(new_n863_));
  NAND2_X1  g662(.A1(new_n860_), .A2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n859_), .A2(new_n864_), .ZN(G1348gat));
  INV_X1    g664(.A(G176gat), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(KEYINPUT125), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n860_), .A2(new_n488_), .A3(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n866_), .A2(KEYINPUT125), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n868_), .B(new_n869_), .ZN(G1349gat));
  NAND2_X1  g669(.A1(new_n860_), .A2(new_n591_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n871_), .A2(new_n263_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n872_), .B1(new_n265_), .B2(new_n871_), .ZN(G1350gat));
  NAND3_X1  g672(.A1(new_n860_), .A2(new_n268_), .A3(new_n589_), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n860_), .A2(new_n559_), .ZN(new_n875_));
  INV_X1    g674(.A(G190gat), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n874_), .B1(new_n875_), .B2(new_n876_), .ZN(G1351gat));
  NAND3_X1  g676(.A1(new_n795_), .A2(new_n393_), .A3(new_n848_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n878_), .A2(new_n523_), .ZN(new_n879_));
  XOR2_X1   g678(.A(new_n879_), .B(G197gat), .Z(G1352gat));
  NOR2_X1   g679(.A1(new_n878_), .A2(new_n487_), .ZN(new_n881_));
  XOR2_X1   g680(.A(new_n881_), .B(G204gat), .Z(G1353gat));
  NOR2_X1   g681(.A1(new_n878_), .A2(new_n579_), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n883_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n884_));
  XOR2_X1   g683(.A(KEYINPUT63), .B(G211gat), .Z(new_n885_));
  AOI21_X1  g684(.A(new_n884_), .B1(new_n883_), .B2(new_n885_), .ZN(G1354gat));
  OAI21_X1  g685(.A(G218gat), .B1(new_n878_), .B2(new_n558_), .ZN(new_n887_));
  OR2_X1    g686(.A1(new_n590_), .A2(G218gat), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n878_), .B2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT126), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n889_), .B(new_n890_), .ZN(G1355gat));
endmodule


