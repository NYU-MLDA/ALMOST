//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 1 0 0 0 1 1 1 0 0 0 0 1 0 1 1 1 1 0 0 1 1 1 0 1 1 1 0 0 0 0 1 0 0 0 0 0 1 0 0 1 1 0 1 1 1 0 1 0 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n747_, new_n748_,
    new_n749_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n798_, new_n799_, new_n800_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n916_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n959_, new_n960_, new_n961_, new_n963_, new_n964_, new_n966_,
    new_n967_, new_n969_, new_n970_, new_n972_, new_n974_, new_n975_,
    new_n976_, new_n978_, new_n979_;
  XNOR2_X1  g000(.A(G141gat), .B(G148gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT86), .ZN(new_n204_));
  INV_X1    g003(.A(G155gat), .ZN(new_n205_));
  INV_X1    g004(.A(G162gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT86), .B1(G155gat), .B2(G162gat), .ZN(new_n208_));
  AND2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT1), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT1), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(G155gat), .A3(G162gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n203_), .B1(new_n209_), .B2(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G141gat), .A2(G148gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT3), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G141gat), .A2(G148gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT2), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n218_), .A2(new_n221_), .A3(new_n222_), .A4(new_n223_), .ZN(new_n224_));
  AOI22_X1  g023(.A1(new_n207_), .A2(new_n208_), .B1(G155gat), .B2(G162gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n215_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT4), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G127gat), .B(G134gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G113gat), .B(G120gat), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n229_), .A2(new_n230_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n227_), .A2(new_n228_), .A3(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G225gat), .A2(G233gat), .ZN(new_n235_));
  XOR2_X1   g034(.A(new_n235_), .B(KEYINPUT102), .Z(new_n236_));
  NAND2_X1  g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  AND2_X1   g037(.A1(new_n224_), .A2(new_n225_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n214_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n207_), .A2(new_n208_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n202_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n233_), .B1(new_n239_), .B2(new_n242_), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n215_), .B(new_n226_), .C1(new_n231_), .C2(new_n232_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT100), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n243_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n227_), .A2(KEYINPUT100), .A3(new_n233_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(KEYINPUT101), .B1(new_n248_), .B2(KEYINPUT4), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT101), .ZN(new_n250_));
  AOI211_X1 g049(.A(new_n250_), .B(new_n228_), .C1(new_n246_), .C2(new_n247_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n238_), .B1(new_n249_), .B2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n248_), .A2(new_n235_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G1gat), .B(G29gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(G85gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT0), .B(G57gat), .ZN(new_n256_));
  XOR2_X1   g055(.A(new_n255_), .B(new_n256_), .Z(new_n257_));
  NAND3_X1  g056(.A1(new_n252_), .A2(new_n253_), .A3(new_n257_), .ZN(new_n258_));
  XOR2_X1   g057(.A(KEYINPUT103), .B(KEYINPUT33), .Z(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT33), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n252_), .A2(new_n261_), .A3(new_n253_), .A4(new_n257_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G8gat), .B(G36gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT18), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G64gat), .B(G92gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  OR2_X1    g066(.A1(G183gat), .A2(G190gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(KEYINPUT82), .B(KEYINPUT23), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G183gat), .A2(G190gat), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n270_), .A2(KEYINPUT23), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n268_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G169gat), .A2(G176gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT98), .ZN(new_n276_));
  INV_X1    g075(.A(G176gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT22), .B(G169gat), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n276_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n274_), .A2(new_n279_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(G169gat), .A2(G176gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n275_), .A2(KEYINPUT24), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n281_), .B1(new_n282_), .B2(KEYINPUT97), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n283_), .B1(KEYINPUT97), .B2(new_n282_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n271_), .A2(KEYINPUT23), .ZN(new_n285_));
  XOR2_X1   g084(.A(KEYINPUT82), .B(KEYINPUT23), .Z(new_n286_));
  AOI21_X1  g085(.A(new_n285_), .B1(new_n286_), .B2(new_n271_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT24), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n281_), .A2(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n284_), .A2(new_n287_), .A3(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT26), .B(G190gat), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(G183gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(KEYINPUT25), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT25), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(G183gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT96), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n294_), .A2(new_n296_), .A3(KEYINPUT96), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n292_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n280_), .B1(new_n290_), .B2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(G197gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(G204gat), .ZN(new_n304_));
  INV_X1    g103(.A(G204gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(G197gat), .ZN(new_n306_));
  AND2_X1   g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT21), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(G218gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(G211gat), .ZN(new_n311_));
  INV_X1    g110(.A(G211gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(G218gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n311_), .A2(new_n313_), .A3(KEYINPUT91), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT91), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n312_), .A2(G218gat), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n310_), .A2(G211gat), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n315_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n309_), .A2(new_n314_), .A3(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n314_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT89), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n304_), .A2(new_n306_), .A3(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT90), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n303_), .A2(KEYINPUT89), .A3(G204gat), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n322_), .A2(new_n323_), .A3(KEYINPUT21), .A4(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n307_), .A2(new_n308_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n320_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  AND2_X1   g126(.A1(new_n324_), .A2(KEYINPUT21), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n323_), .B1(new_n328_), .B2(new_n322_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n319_), .B1(new_n327_), .B2(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT20), .B1(new_n302_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT80), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n332_), .A2(new_n295_), .A3(G183gat), .ZN(new_n333_));
  OAI21_X1  g132(.A(KEYINPUT80), .B1(new_n293_), .B2(KEYINPUT25), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n291_), .A2(new_n294_), .A3(new_n333_), .A4(new_n334_), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n282_), .A2(new_n281_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT81), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n335_), .A2(KEYINPUT81), .A3(new_n336_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n286_), .A2(new_n270_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n341_), .B1(KEYINPUT23), .B2(new_n270_), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n339_), .A2(new_n340_), .A3(new_n342_), .A4(new_n289_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n287_), .A2(new_n268_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(G169gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n329_), .ZN(new_n348_));
  AOI22_X1  g147(.A1(new_n318_), .A2(new_n314_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n348_), .A2(new_n325_), .A3(new_n349_), .ZN(new_n350_));
  AOI22_X1  g149(.A1(new_n343_), .A2(new_n347_), .B1(new_n350_), .B2(new_n319_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G226gat), .A2(G233gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  NOR3_X1   g153(.A1(new_n331_), .A2(new_n351_), .A3(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n354_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT20), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n357_), .B1(new_n302_), .B2(new_n330_), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n343_), .A2(new_n347_), .A3(new_n350_), .A4(new_n319_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n356_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n267_), .B1(new_n355_), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n358_), .A2(new_n359_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(new_n354_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n267_), .ZN(new_n364_));
  OR2_X1    g163(.A1(new_n302_), .A2(new_n330_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n342_), .A2(new_n340_), .A3(new_n289_), .ZN(new_n366_));
  AOI21_X1  g165(.A(KEYINPUT81), .B1(new_n335_), .B2(new_n336_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n347_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(new_n330_), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n365_), .A2(new_n369_), .A3(KEYINPUT20), .A4(new_n356_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n363_), .A2(new_n364_), .A3(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n361_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT99), .ZN(new_n373_));
  OAI211_X1 g172(.A(new_n235_), .B(new_n234_), .C1(new_n249_), .C2(new_n251_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n257_), .B1(new_n248_), .B2(new_n236_), .ZN(new_n375_));
  AOI22_X1  g174(.A1(new_n372_), .A2(new_n373_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n361_), .A2(KEYINPUT99), .A3(new_n371_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n263_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n257_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n248_), .A2(KEYINPUT4), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(new_n250_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n248_), .A2(KEYINPUT101), .A3(KEYINPUT4), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n237_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n253_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n379_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT104), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(new_n386_), .A3(new_n258_), .ZN(new_n387_));
  OAI211_X1 g186(.A(KEYINPUT104), .B(new_n379_), .C1(new_n383_), .C2(new_n384_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n364_), .A2(KEYINPUT32), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n389_), .B1(new_n355_), .B2(new_n360_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n354_), .B1(new_n331_), .B2(new_n351_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n358_), .A2(new_n359_), .A3(new_n356_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n390_), .B1(new_n393_), .B2(new_n389_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n387_), .A2(new_n388_), .A3(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n378_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n227_), .A2(KEYINPUT29), .ZN(new_n397_));
  INV_X1    g196(.A(G228gat), .ZN(new_n398_));
  NOR2_X1   g197(.A1(KEYINPUT88), .A2(G233gat), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(KEYINPUT88), .A2(G233gat), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n398_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT92), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n330_), .A2(new_n397_), .A3(new_n403_), .ZN(new_n404_));
  AOI22_X1  g203(.A1(new_n350_), .A2(new_n319_), .B1(new_n227_), .B2(KEYINPUT29), .ZN(new_n405_));
  XOR2_X1   g204(.A(new_n402_), .B(KEYINPUT92), .Z(new_n406_));
  OAI21_X1  g205(.A(new_n404_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G78gat), .B(G106gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n408_), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n404_), .B(new_n410_), .C1(new_n405_), .C2(new_n406_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT93), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n411_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT94), .ZN(new_n415_));
  XNOR2_X1  g214(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n417_), .B1(new_n227_), .B2(KEYINPUT29), .ZN(new_n418_));
  XOR2_X1   g217(.A(G22gat), .B(G50gat), .Z(new_n419_));
  INV_X1    g218(.A(KEYINPUT29), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n215_), .A2(new_n420_), .A3(new_n226_), .A4(new_n416_), .ZN(new_n421_));
  AND3_X1   g220(.A1(new_n418_), .A2(new_n419_), .A3(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n419_), .B1(new_n418_), .B2(new_n421_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  AND3_X1   g223(.A1(new_n414_), .A2(new_n415_), .A3(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n415_), .B1(new_n414_), .B2(new_n424_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n412_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n414_), .A2(new_n424_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(KEYINPUT94), .ZN(new_n429_));
  INV_X1    g228(.A(new_n412_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n414_), .A2(new_n415_), .A3(new_n424_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n429_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n427_), .A2(new_n432_), .ZN(new_n433_));
  OAI211_X1 g232(.A(KEYINPUT30), .B(new_n347_), .C1(new_n366_), .C2(new_n367_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(KEYINPUT30), .B1(new_n343_), .B2(new_n347_), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT84), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT30), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n368_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT84), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n439_), .A2(new_n440_), .A3(new_n434_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G227gat), .A2(G233gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(KEYINPUT83), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G71gat), .B(G99gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  XOR2_X1   g244(.A(G15gat), .B(G43gat), .Z(new_n446_));
  XNOR2_X1  g245(.A(new_n445_), .B(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n437_), .A2(new_n441_), .A3(new_n447_), .ZN(new_n448_));
  OR2_X1    g247(.A1(new_n233_), .A2(KEYINPUT31), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n233_), .A2(KEYINPUT31), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n449_), .A2(KEYINPUT85), .A3(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n447_), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n452_), .A2(new_n439_), .A3(new_n440_), .A4(new_n434_), .ZN(new_n453_));
  AND3_X1   g252(.A1(new_n448_), .A2(new_n451_), .A3(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n451_), .B1(new_n448_), .B2(new_n453_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n433_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n448_), .A2(new_n453_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n451_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n448_), .A2(new_n451_), .A3(new_n453_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NOR3_X1   g262(.A1(new_n425_), .A2(new_n426_), .A3(new_n412_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n430_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n463_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n456_), .A2(new_n432_), .A3(new_n427_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT27), .ZN(new_n469_));
  NOR3_X1   g268(.A1(new_n355_), .A2(new_n360_), .A3(new_n267_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n364_), .B1(new_n363_), .B2(new_n370_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n469_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n393_), .A2(new_n267_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n473_), .A2(KEYINPUT27), .A3(new_n371_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n475_), .B1(new_n388_), .B2(new_n387_), .ZN(new_n476_));
  AOI22_X1  g275(.A1(new_n396_), .A2(new_n458_), .B1(new_n468_), .B2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G29gat), .B(G36gat), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  XOR2_X1   g278(.A(G43gat), .B(G50gat), .Z(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G43gat), .B(G50gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n478_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n481_), .A2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G1gat), .B(G8gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT74), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G15gat), .B(G22gat), .ZN(new_n487_));
  INV_X1    g286(.A(G1gat), .ZN(new_n488_));
  INV_X1    g287(.A(G8gat), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT14), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n487_), .A2(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n486_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n491_), .ZN(new_n493_));
  OR2_X1    g292(.A1(new_n485_), .A2(KEYINPUT74), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n485_), .A2(KEYINPUT74), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n493_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n484_), .B1(new_n492_), .B2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT15), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n484_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n486_), .A2(new_n491_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n493_), .A2(new_n494_), .A3(new_n495_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n481_), .A2(KEYINPUT15), .A3(new_n483_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n499_), .A2(new_n500_), .A3(new_n501_), .A4(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G229gat), .A2(G233gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(KEYINPUT76), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n497_), .A2(new_n503_), .A3(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT77), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n504_), .ZN(new_n509_));
  NOR3_X1   g308(.A1(new_n492_), .A2(new_n496_), .A3(new_n484_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n484_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n511_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n509_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n497_), .A2(new_n503_), .A3(KEYINPUT77), .A4(new_n505_), .ZN(new_n514_));
  XOR2_X1   g313(.A(G113gat), .B(G141gat), .Z(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT78), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G169gat), .B(G197gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n508_), .A2(new_n513_), .A3(new_n514_), .A4(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT79), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n513_), .A2(new_n514_), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n522_), .A2(KEYINPUT79), .A3(new_n508_), .A4(new_n518_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n508_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n518_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n524_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n477_), .A2(new_n529_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n492_), .A2(new_n496_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT75), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G231gat), .A2(G233gat), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n532_), .B(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G57gat), .B(G64gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G71gat), .B(G78gat), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n536_), .A2(new_n537_), .A3(KEYINPUT11), .ZN(new_n538_));
  XOR2_X1   g337(.A(G71gat), .B(G78gat), .Z(new_n539_));
  INV_X1    g338(.A(G64gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(G57gat), .ZN(new_n541_));
  INV_X1    g340(.A(G57gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(G64gat), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n541_), .A2(new_n543_), .A3(KEYINPUT11), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n539_), .A2(new_n544_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n536_), .A2(KEYINPUT11), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n538_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n535_), .A2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n532_), .B(new_n533_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n547_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G127gat), .B(G155gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT16), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G183gat), .B(G211gat), .ZN(new_n554_));
  XOR2_X1   g353(.A(new_n553_), .B(new_n554_), .Z(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n548_), .A2(new_n551_), .A3(KEYINPUT17), .A4(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT70), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n547_), .B(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n549_), .A2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n547_), .B(KEYINPUT70), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n535_), .A2(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n555_), .B(KEYINPUT17), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n560_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  AND2_X1   g363(.A1(new_n557_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT13), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G230gat), .A2(G233gat), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G99gat), .A2(G106gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT6), .ZN(new_n570_));
  OAI21_X1  g369(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n571_));
  NOR2_X1   g370(.A1(G99gat), .A2(G106gat), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT7), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n570_), .A2(new_n571_), .A3(new_n574_), .ZN(new_n575_));
  XOR2_X1   g374(.A(G85gat), .B(G92gat), .Z(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(KEYINPUT8), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT68), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT6), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n569_), .B(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n574_), .A2(new_n571_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n579_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n570_), .A2(KEYINPUT68), .A3(new_n571_), .A4(new_n574_), .ZN(new_n584_));
  XOR2_X1   g383(.A(KEYINPUT69), .B(KEYINPUT8), .Z(new_n585_));
  NAND4_X1  g384(.A1(new_n583_), .A2(new_n584_), .A3(new_n576_), .A4(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(G85gat), .A2(G92gat), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(KEYINPUT66), .B(KEYINPUT9), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT67), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G85gat), .A2(G92gat), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n590_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n591_), .B1(new_n590_), .B2(new_n592_), .ZN(new_n595_));
  OAI211_X1 g394(.A(new_n588_), .B(new_n589_), .C1(new_n594_), .C2(new_n595_), .ZN(new_n596_));
  OR2_X1    g395(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n597_));
  NAND2_X1  g396(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(KEYINPUT64), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT64), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n597_), .A2(new_n601_), .A3(new_n598_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(KEYINPUT65), .B(G106gat), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n581_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  AOI22_X1  g404(.A1(new_n578_), .A2(new_n586_), .B1(new_n596_), .B2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(new_n559_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n606_), .A2(new_n559_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n568_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT12), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n611_), .B1(new_n606_), .B2(new_n559_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n550_), .A2(KEYINPUT12), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n596_), .A2(new_n605_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n585_), .A2(new_n576_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n617_), .B1(new_n575_), .B2(new_n579_), .ZN(new_n618_));
  AOI22_X1  g417(.A1(new_n618_), .A2(new_n584_), .B1(new_n577_), .B2(KEYINPUT8), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n614_), .B1(new_n616_), .B2(new_n619_), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n612_), .A2(new_n567_), .A3(new_n620_), .A4(new_n607_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G120gat), .B(G148gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT5), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G176gat), .B(G204gat), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n623_), .B(new_n624_), .Z(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n610_), .A2(new_n621_), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n626_), .B1(new_n610_), .B2(new_n621_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n566_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n629_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n631_), .A2(KEYINPUT13), .A3(new_n627_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(G232gat), .A2(G233gat), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT34), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT35), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT72), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n606_), .A2(new_n639_), .A3(new_n484_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n639_), .B1(new_n606_), .B2(new_n484_), .ZN(new_n641_));
  OAI22_X1  g440(.A1(new_n640_), .A2(new_n641_), .B1(KEYINPUT35), .B2(new_n635_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n578_), .A2(new_n586_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(new_n615_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n499_), .A2(new_n502_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n644_), .A2(KEYINPUT71), .A3(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT71), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n648_), .B1(new_n606_), .B2(new_n645_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n638_), .B1(new_n642_), .B2(new_n650_), .ZN(new_n651_));
  XOR2_X1   g450(.A(G190gat), .B(G218gat), .Z(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT73), .ZN(new_n653_));
  XNOR2_X1  g452(.A(G134gat), .B(G162gat), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n653_), .B(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n655_), .A2(KEYINPUT36), .ZN(new_n656_));
  OAI21_X1  g455(.A(KEYINPUT72), .B1(new_n644_), .B2(new_n511_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n606_), .A2(new_n639_), .A3(new_n484_), .ZN(new_n658_));
  AOI22_X1  g457(.A1(new_n657_), .A2(new_n658_), .B1(new_n637_), .B2(new_n636_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n638_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n647_), .A2(new_n649_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n659_), .A2(new_n660_), .A3(new_n661_), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n651_), .A2(new_n656_), .A3(new_n662_), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n655_), .B(KEYINPUT36), .Z(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n665_), .B1(new_n651_), .B2(new_n662_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n663_), .A2(new_n666_), .A3(KEYINPUT37), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT37), .ZN(new_n668_));
  NOR3_X1   g467(.A1(new_n642_), .A2(new_n650_), .A3(new_n638_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n660_), .B1(new_n659_), .B2(new_n661_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n664_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n651_), .A2(new_n662_), .A3(new_n656_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n668_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  OAI211_X1 g472(.A(new_n565_), .B(new_n633_), .C1(new_n667_), .C2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n530_), .A2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n387_), .A2(new_n388_), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n676_), .A2(G1gat), .A3(new_n677_), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n678_), .A2(KEYINPUT38), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(KEYINPUT38), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n663_), .A2(new_n666_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n477_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n633_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n557_), .A2(new_n564_), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n683_), .A2(new_n529_), .A3(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n682_), .A2(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(G1gat), .B1(new_n686_), .B2(new_n677_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n679_), .A2(new_n680_), .A3(new_n687_), .ZN(G1324gat));
  INV_X1    g487(.A(new_n676_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n689_), .A2(new_n489_), .A3(new_n475_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT39), .ZN(new_n691_));
  INV_X1    g490(.A(new_n686_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(new_n475_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n691_), .B1(new_n693_), .B2(G8gat), .ZN(new_n694_));
  AOI211_X1 g493(.A(KEYINPUT39), .B(new_n489_), .C1(new_n692_), .C2(new_n475_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n690_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT40), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n696_), .B(new_n697_), .ZN(G1325gat));
  OAI21_X1  g497(.A(G15gat), .B1(new_n686_), .B2(new_n456_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT41), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n676_), .A2(G15gat), .A3(new_n456_), .ZN(new_n701_));
  OR2_X1    g500(.A1(new_n700_), .A2(new_n701_), .ZN(G1326gat));
  OAI21_X1  g501(.A(G22gat), .B1(new_n686_), .B2(new_n433_), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT42), .Z(new_n704_));
  NOR3_X1   g503(.A1(new_n676_), .A2(G22gat), .A3(new_n433_), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1327gat));
  INV_X1    g505(.A(new_n681_), .ZN(new_n707_));
  NOR3_X1   g506(.A1(new_n565_), .A2(new_n683_), .A3(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n530_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n677_), .ZN(new_n711_));
  AOI21_X1  g510(.A(G29gat), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(KEYINPUT37), .B1(new_n663_), .B2(new_n666_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n671_), .A2(new_n668_), .A3(new_n672_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  OAI21_X1  g514(.A(KEYINPUT43), .B1(new_n477_), .B2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT43), .ZN(new_n717_));
  INV_X1    g516(.A(new_n715_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n468_), .A2(new_n476_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n457_), .B1(new_n378_), .B2(new_n395_), .ZN(new_n720_));
  OAI211_X1 g519(.A(new_n717_), .B(new_n718_), .C1(new_n719_), .C2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n716_), .A2(new_n721_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n633_), .A2(new_n528_), .A3(new_n684_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT105), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n722_), .A2(KEYINPUT44), .A3(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(KEYINPUT44), .B1(new_n722_), .B2(new_n724_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n711_), .A2(G29gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n712_), .B1(new_n727_), .B2(new_n728_), .ZN(G1328gat));
  INV_X1    g528(.A(G36gat), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n475_), .A2(new_n730_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n709_), .A2(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n732_), .B(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n475_), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n725_), .A2(new_n726_), .A3(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n734_), .B1(new_n736_), .B2(new_n730_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT46), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  OAI211_X1 g538(.A(KEYINPUT46), .B(new_n734_), .C1(new_n736_), .C2(new_n730_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(G1329gat));
  AOI21_X1  g540(.A(G43gat), .B1(new_n710_), .B2(new_n463_), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n463_), .A2(G43gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n727_), .B2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT47), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n744_), .B(new_n745_), .ZN(G1330gat));
  INV_X1    g545(.A(new_n433_), .ZN(new_n747_));
  AOI21_X1  g546(.A(G50gat), .B1(new_n710_), .B2(new_n747_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n747_), .A2(G50gat), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n727_), .B2(new_n749_), .ZN(G1331gat));
  OAI21_X1  g549(.A(KEYINPUT107), .B1(new_n477_), .B2(new_n528_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT107), .ZN(new_n752_));
  OAI211_X1 g551(.A(new_n752_), .B(new_n529_), .C1(new_n719_), .C2(new_n720_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n751_), .A2(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n684_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n755_));
  AND3_X1   g554(.A1(new_n754_), .A2(new_n683_), .A3(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n756_), .A2(new_n542_), .A3(new_n711_), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n633_), .A2(new_n684_), .A3(new_n528_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n682_), .A2(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(G57gat), .B1(new_n759_), .B2(new_n677_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n757_), .A2(new_n760_), .ZN(G1332gat));
  NAND3_X1  g560(.A1(new_n756_), .A2(new_n540_), .A3(new_n475_), .ZN(new_n762_));
  OAI21_X1  g561(.A(G64gat), .B1(new_n759_), .B2(new_n735_), .ZN(new_n763_));
  OR2_X1    g562(.A1(new_n763_), .A2(KEYINPUT109), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(KEYINPUT109), .ZN(new_n765_));
  XNOR2_X1  g564(.A(KEYINPUT108), .B(KEYINPUT48), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n764_), .A2(new_n765_), .A3(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n762_), .B1(new_n767_), .B2(new_n768_), .ZN(G1333gat));
  OAI21_X1  g568(.A(G71gat), .B1(new_n759_), .B2(new_n456_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT49), .ZN(new_n771_));
  INV_X1    g570(.A(G71gat), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n756_), .A2(new_n772_), .A3(new_n463_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(G1334gat));
  NAND3_X1  g573(.A1(new_n682_), .A2(new_n747_), .A3(new_n758_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(G78gat), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT50), .ZN(new_n777_));
  INV_X1    g576(.A(G78gat), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n756_), .A2(new_n778_), .A3(new_n747_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT110), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n780_), .B(new_n781_), .ZN(G1335gat));
  NAND3_X1  g581(.A1(new_n683_), .A2(new_n529_), .A3(new_n684_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n783_), .B1(new_n716_), .B2(new_n721_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT111), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n784_), .A2(new_n785_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n711_), .A2(G85gat), .ZN(new_n788_));
  XOR2_X1   g587(.A(new_n788_), .B(KEYINPUT112), .Z(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  NOR3_X1   g589(.A1(new_n786_), .A2(new_n787_), .A3(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n683_), .A2(new_n684_), .A3(new_n681_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n792_), .B1(new_n751_), .B2(new_n753_), .ZN(new_n793_));
  AOI21_X1  g592(.A(G85gat), .B1(new_n793_), .B2(new_n711_), .ZN(new_n794_));
  OR3_X1    g593(.A1(new_n791_), .A2(KEYINPUT113), .A3(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(KEYINPUT113), .B1(new_n791_), .B2(new_n794_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(G1336gat));
  AOI21_X1  g596(.A(G92gat), .B1(new_n793_), .B2(new_n475_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n786_), .A2(new_n787_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n475_), .A2(G92gat), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n798_), .B1(new_n799_), .B2(new_n800_), .ZN(G1337gat));
  NAND2_X1  g600(.A1(new_n463_), .A2(new_n603_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n793_), .A2(new_n803_), .ZN(new_n804_));
  AOI211_X1 g603(.A(new_n456_), .B(new_n783_), .C1(new_n716_), .C2(new_n721_), .ZN(new_n805_));
  INV_X1    g604(.A(G99gat), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n804_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(KEYINPUT116), .B(KEYINPUT51), .ZN(new_n808_));
  OR2_X1    g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT115), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT51), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT114), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n811_), .B1(new_n807_), .B2(new_n812_), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n804_), .B(KEYINPUT114), .C1(new_n805_), .C2(new_n806_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n810_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n806_), .B1(new_n784_), .B2(new_n463_), .ZN(new_n816_));
  AOI211_X1 g615(.A(new_n792_), .B(new_n802_), .C1(new_n751_), .C2(new_n753_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n812_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  AND4_X1   g617(.A1(new_n810_), .A2(new_n818_), .A3(KEYINPUT51), .A4(new_n814_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n809_), .B1(new_n815_), .B2(new_n819_), .ZN(G1338gat));
  NAND3_X1  g619(.A1(new_n793_), .A2(new_n747_), .A3(new_n604_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n784_), .A2(new_n747_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n823_));
  AND3_X1   g622(.A1(new_n822_), .A2(new_n823_), .A3(G106gat), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n823_), .B1(new_n822_), .B2(G106gat), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n821_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n826_), .B(KEYINPUT53), .ZN(G1339gat));
  OAI21_X1  g626(.A(KEYINPUT54), .B1(new_n674_), .B2(new_n528_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT54), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n755_), .A2(new_n829_), .A3(new_n529_), .A4(new_n633_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n828_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT56), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n832_), .A2(KEYINPUT119), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n612_), .A2(new_n607_), .A3(new_n620_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n568_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT55), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n835_), .B1(new_n836_), .B2(new_n621_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT117), .ZN(new_n838_));
  AND3_X1   g637(.A1(new_n621_), .A2(new_n838_), .A3(new_n836_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n838_), .B1(new_n621_), .B2(new_n836_), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n837_), .A2(new_n839_), .A3(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n833_), .B1(new_n841_), .B2(new_n626_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n621_), .A2(new_n836_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(KEYINPUT117), .ZN(new_n844_));
  OR2_X1    g643(.A1(new_n621_), .A2(new_n836_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n621_), .A2(new_n838_), .A3(new_n836_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n844_), .A2(new_n845_), .A3(new_n846_), .A4(new_n835_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n847_), .A2(new_n625_), .A3(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n505_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n497_), .A2(new_n503_), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n850_), .B(new_n526_), .C1(new_n851_), .C2(new_n505_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n524_), .A2(new_n627_), .A3(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n842_), .A2(new_n849_), .A3(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT58), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n715_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n842_), .A2(KEYINPUT58), .A3(new_n849_), .A4(new_n854_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT120), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n847_), .A2(new_n625_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n853_), .B1(new_n861_), .B2(new_n833_), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n862_), .A2(KEYINPUT120), .A3(KEYINPUT58), .A4(new_n849_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n857_), .A2(new_n860_), .A3(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT57), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n628_), .A2(new_n629_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n524_), .A2(new_n852_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n528_), .A2(new_n627_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n832_), .A2(KEYINPUT118), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n869_), .B1(new_n861_), .B2(new_n870_), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n847_), .A2(KEYINPUT118), .A3(new_n832_), .A4(new_n625_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n868_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n865_), .B1(new_n873_), .B2(new_n681_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n870_), .B1(new_n841_), .B2(new_n626_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n869_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n875_), .A2(new_n876_), .A3(new_n872_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n868_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n879_), .A2(KEYINPUT57), .A3(new_n707_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n864_), .A2(new_n874_), .A3(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n831_), .B1(new_n881_), .B2(new_n684_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n711_), .A2(new_n735_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(new_n466_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(KEYINPUT121), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n883_), .A2(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(G113gat), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n888_), .A2(new_n889_), .A3(new_n528_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT59), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n887_), .A2(new_n891_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n883_), .A2(KEYINPUT59), .A3(new_n886_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n529_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n890_), .B1(new_n894_), .B2(new_n889_), .ZN(G1340gat));
  INV_X1    g694(.A(G120gat), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n896_), .B1(new_n633_), .B2(KEYINPUT60), .ZN(new_n897_));
  OAI211_X1 g696(.A(new_n888_), .B(new_n897_), .C1(KEYINPUT60), .C2(new_n896_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n633_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n899_), .B2(new_n896_), .ZN(G1341gat));
  INV_X1    g699(.A(G127gat), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n888_), .A2(new_n901_), .A3(new_n565_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n684_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n902_), .B1(new_n903_), .B2(new_n901_), .ZN(G1342gat));
  AOI21_X1  g703(.A(G134gat), .B1(new_n888_), .B2(new_n681_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n892_), .A2(new_n893_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(KEYINPUT122), .B(G134gat), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n715_), .A2(new_n907_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n905_), .B1(new_n906_), .B2(new_n908_), .ZN(G1343gat));
  NOR2_X1   g708(.A1(new_n884_), .A2(new_n467_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(KEYINPUT123), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n882_), .A2(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(new_n528_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g714(.A1(new_n913_), .A2(new_n683_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g716(.A(KEYINPUT61), .B(G155gat), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT124), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n913_), .A2(new_n920_), .A3(new_n565_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n921_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n920_), .B1(new_n913_), .B2(new_n565_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n919_), .B1(new_n922_), .B2(new_n923_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n923_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n925_), .A2(new_n921_), .A3(new_n918_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n924_), .A2(new_n926_), .ZN(G1346gat));
  NAND2_X1  g726(.A1(new_n883_), .A2(new_n911_), .ZN(new_n928_));
  NOR3_X1   g727(.A1(new_n928_), .A2(new_n206_), .A3(new_n715_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n206_), .B1(new_n928_), .B2(new_n707_), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT125), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(new_n932_));
  OAI211_X1 g731(.A(KEYINPUT125), .B(new_n206_), .C1(new_n928_), .C2(new_n707_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n929_), .B1(new_n932_), .B2(new_n933_), .ZN(G1347gat));
  NOR2_X1   g733(.A1(new_n711_), .A2(new_n735_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(new_n463_), .ZN(new_n936_));
  NOR3_X1   g735(.A1(new_n882_), .A2(new_n747_), .A3(new_n936_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n937_), .A2(new_n528_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n938_), .A2(G169gat), .ZN(new_n939_));
  INV_X1    g738(.A(KEYINPUT62), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n939_), .A2(new_n940_), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n937_), .A2(new_n278_), .A3(new_n528_), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n938_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n941_), .A2(new_n942_), .A3(new_n943_), .ZN(G1348gat));
  INV_X1    g743(.A(KEYINPUT126), .ZN(new_n945_));
  AOI21_X1  g744(.A(KEYINPUT57), .B1(new_n879_), .B2(new_n707_), .ZN(new_n946_));
  AOI211_X1 g745(.A(new_n865_), .B(new_n681_), .C1(new_n877_), .C2(new_n878_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n946_), .A2(new_n947_), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n565_), .B1(new_n948_), .B2(new_n864_), .ZN(new_n949_));
  OAI211_X1 g748(.A(new_n945_), .B(new_n433_), .C1(new_n949_), .C2(new_n831_), .ZN(new_n950_));
  OAI21_X1  g749(.A(KEYINPUT126), .B1(new_n882_), .B2(new_n747_), .ZN(new_n951_));
  NOR3_X1   g750(.A1(new_n936_), .A2(new_n277_), .A3(new_n633_), .ZN(new_n952_));
  AND3_X1   g751(.A1(new_n950_), .A2(new_n951_), .A3(new_n952_), .ZN(new_n953_));
  AOI21_X1  g752(.A(G176gat), .B1(new_n937_), .B2(new_n683_), .ZN(new_n954_));
  OAI21_X1  g753(.A(KEYINPUT127), .B1(new_n953_), .B2(new_n954_), .ZN(new_n955_));
  INV_X1    g754(.A(new_n936_), .ZN(new_n956_));
  NAND3_X1  g755(.A1(new_n883_), .A2(new_n433_), .A3(new_n956_), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n277_), .B1(new_n957_), .B2(new_n633_), .ZN(new_n958_));
  NAND3_X1  g757(.A1(new_n950_), .A2(new_n951_), .A3(new_n952_), .ZN(new_n959_));
  INV_X1    g758(.A(KEYINPUT127), .ZN(new_n960_));
  NAND3_X1  g759(.A1(new_n958_), .A2(new_n959_), .A3(new_n960_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n955_), .A2(new_n961_), .ZN(G1349gat));
  NAND4_X1  g761(.A1(new_n950_), .A2(new_n951_), .A3(new_n565_), .A4(new_n956_), .ZN(new_n963_));
  AND3_X1   g762(.A1(new_n565_), .A2(new_n300_), .A3(new_n299_), .ZN(new_n964_));
  AOI22_X1  g763(.A1(new_n963_), .A2(new_n293_), .B1(new_n937_), .B2(new_n964_), .ZN(G1350gat));
  OAI21_X1  g764(.A(G190gat), .B1(new_n957_), .B2(new_n715_), .ZN(new_n966_));
  NAND3_X1  g765(.A1(new_n937_), .A2(new_n291_), .A3(new_n681_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n966_), .A2(new_n967_), .ZN(G1351gat));
  NOR4_X1   g767(.A1(new_n882_), .A2(new_n467_), .A3(new_n711_), .A4(new_n735_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n969_), .A2(new_n528_), .ZN(new_n970_));
  XNOR2_X1  g769(.A(new_n970_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g770(.A1(new_n969_), .A2(new_n683_), .ZN(new_n972_));
  XNOR2_X1  g771(.A(new_n972_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g772(.A(KEYINPUT63), .B(G211gat), .C1(new_n969_), .C2(new_n565_), .ZN(new_n974_));
  XOR2_X1   g773(.A(KEYINPUT63), .B(G211gat), .Z(new_n975_));
  AND3_X1   g774(.A1(new_n969_), .A2(new_n565_), .A3(new_n975_), .ZN(new_n976_));
  NOR2_X1   g775(.A1(new_n974_), .A2(new_n976_), .ZN(G1354gat));
  NAND3_X1  g776(.A1(new_n969_), .A2(new_n310_), .A3(new_n681_), .ZN(new_n978_));
  AND2_X1   g777(.A1(new_n969_), .A2(new_n718_), .ZN(new_n979_));
  OAI21_X1  g778(.A(new_n978_), .B1(new_n979_), .B2(new_n310_), .ZN(G1355gat));
endmodule


