//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 1 1 0 1 1 1 0 1 1 1 1 0 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 0 1 0 1 0 1 0 0 1 1 0 0 1 1 1 0 0 0 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n801_, new_n802_,
    new_n803_, new_n805_, new_n806_, new_n807_, new_n808_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n896_, new_n898_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n908_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n927_, new_n928_,
    new_n929_, new_n931_, new_n932_, new_n934_, new_n935_, new_n936_,
    new_n937_, new_n939_, new_n940_, new_n941_, new_n942_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_,
    new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_,
    new_n969_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n978_, new_n979_;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT19), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G183gat), .A2(G190gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT23), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n206_), .A2(G183gat), .A3(G190gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  AND2_X1   g008(.A1(KEYINPUT82), .A2(G190gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(KEYINPUT82), .A2(G190gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT26), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  OR2_X1    g011(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT25), .B(G183gat), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n209_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT24), .ZN(new_n217_));
  INV_X1    g016(.A(G169gat), .ZN(new_n218_));
  INV_X1    g017(.A(G176gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n218_), .A2(new_n219_), .A3(KEYINPUT83), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT83), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n221_), .B1(G169gat), .B2(G176gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT84), .ZN(new_n223_));
  AND3_X1   g022(.A1(new_n220_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n223_), .B1(new_n220_), .B2(new_n222_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n217_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n220_), .A2(new_n222_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT84), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n220_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n217_), .B1(G169gat), .B2(G176gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n228_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n216_), .A2(new_n226_), .A3(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(G197gat), .ZN(new_n233_));
  INV_X1    g032(.A(G204gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G197gat), .A2(G204gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT21), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n235_), .A2(KEYINPUT21), .A3(new_n236_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G211gat), .B(G218gat), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n239_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  OR2_X1    g041(.A1(new_n240_), .A2(new_n241_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G169gat), .A2(G176gat), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT22), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n247_), .A2(KEYINPUT85), .A3(G169gat), .ZN(new_n248_));
  AND2_X1   g047(.A1(KEYINPUT85), .A2(G169gat), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n248_), .B(new_n219_), .C1(new_n247_), .C2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT86), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n251_), .B1(new_n204_), .B2(KEYINPUT23), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n252_), .B1(new_n208_), .B2(new_n251_), .ZN(new_n253_));
  NOR3_X1   g052(.A1(new_n210_), .A2(new_n211_), .A3(G183gat), .ZN(new_n254_));
  OAI211_X1 g053(.A(new_n246_), .B(new_n250_), .C1(new_n253_), .C2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n232_), .A2(new_n245_), .A3(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT20), .ZN(new_n257_));
  AOI21_X1  g056(.A(KEYINPUT24), .B1(new_n220_), .B2(new_n222_), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT97), .B1(new_n253_), .B2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n227_), .A2(new_n217_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT97), .ZN(new_n261_));
  AOI21_X1  g060(.A(KEYINPUT86), .B1(new_n205_), .B2(new_n207_), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n260_), .B(new_n261_), .C1(new_n262_), .C2(new_n252_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT26), .B(G190gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(new_n215_), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n259_), .A2(new_n263_), .A3(new_n231_), .A4(new_n265_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n208_), .B1(G183gat), .B2(G190gat), .ZN(new_n267_));
  XOR2_X1   g066(.A(KEYINPUT22), .B(G169gat), .Z(new_n268_));
  OAI211_X1 g067(.A(new_n267_), .B(new_n246_), .C1(G176gat), .C2(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n245_), .B1(new_n266_), .B2(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n203_), .B1(new_n257_), .B2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n232_), .A2(new_n255_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(new_n244_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n266_), .A2(new_n245_), .A3(new_n269_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n203_), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n273_), .A2(new_n274_), .A3(KEYINPUT20), .A4(new_n275_), .ZN(new_n276_));
  XOR2_X1   g075(.A(G8gat), .B(G36gat), .Z(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  XOR2_X1   g078(.A(G64gat), .B(G92gat), .Z(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  AND3_X1   g080(.A1(new_n271_), .A2(new_n276_), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT27), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n273_), .A2(new_n274_), .A3(KEYINPUT20), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(new_n203_), .ZN(new_n286_));
  NOR3_X1   g085(.A1(new_n257_), .A2(new_n270_), .A3(new_n203_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT102), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n286_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  NOR4_X1   g088(.A1(new_n257_), .A2(new_n270_), .A3(KEYINPUT102), .A4(new_n203_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n284_), .B1(new_n291_), .B2(new_n281_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n281_), .B1(new_n271_), .B2(new_n276_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n283_), .B1(new_n282_), .B2(new_n293_), .ZN(new_n294_));
  AND2_X1   g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G141gat), .A2(G148gat), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT92), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT2), .ZN(new_n299_));
  NAND3_X1  g098(.A1(KEYINPUT92), .A2(G141gat), .A3(G148gat), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n298_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT93), .ZN(new_n302_));
  INV_X1    g101(.A(G141gat), .ZN(new_n303_));
  INV_X1    g102(.A(G148gat), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n302_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT3), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT3), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n302_), .A2(new_n307_), .A3(new_n303_), .A4(new_n304_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n301_), .A2(new_n306_), .A3(new_n308_), .A4(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(G155gat), .ZN(new_n311_));
  INV_X1    g110(.A(G162gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G155gat), .A2(G162gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  OR2_X1    g115(.A1(new_n315_), .A2(KEYINPUT1), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n303_), .A2(new_n304_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n319_));
  AND4_X1   g118(.A1(new_n298_), .A2(new_n318_), .A3(new_n300_), .A4(new_n319_), .ZN(new_n320_));
  AOI22_X1  g119(.A1(new_n310_), .A2(new_n316_), .B1(new_n317_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT29), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n244_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(G228gat), .ZN(new_n324_));
  INV_X1    g123(.A(G233gat), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n323_), .A2(new_n326_), .ZN(new_n327_));
  OAI221_X1 g126(.A(new_n244_), .B1(new_n324_), .B2(new_n325_), .C1(new_n321_), .C2(new_n322_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G78gat), .B(G106gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n310_), .A2(new_n316_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n317_), .A2(new_n320_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(KEYINPUT28), .B1(new_n334_), .B2(KEYINPUT29), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT28), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n321_), .A2(new_n336_), .A3(new_n322_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G22gat), .B(G50gat), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n335_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n335_), .A2(new_n337_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n338_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n330_), .B(KEYINPUT95), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n327_), .A2(new_n328_), .A3(new_n343_), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n331_), .A2(new_n339_), .A3(new_n342_), .A4(new_n344_), .ZN(new_n345_));
  AND3_X1   g144(.A1(new_n342_), .A2(KEYINPUT94), .A3(new_n339_), .ZN(new_n346_));
  AOI21_X1  g145(.A(KEYINPUT94), .B1(new_n342_), .B2(new_n339_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n343_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n329_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT96), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n350_), .A2(new_n351_), .A3(new_n344_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n329_), .A2(KEYINPUT96), .A3(new_n349_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n345_), .B1(new_n348_), .B2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G1gat), .B(G29gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G57gat), .B(G85gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G225gat), .A2(G233gat), .ZN(new_n362_));
  INV_X1    g161(.A(G134gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(G127gat), .ZN(new_n364_));
  INV_X1    g163(.A(G127gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(G134gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n364_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(G120gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(G113gat), .ZN(new_n369_));
  INV_X1    g168(.A(G113gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(G120gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n369_), .A2(new_n371_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n367_), .A2(new_n372_), .ZN(new_n373_));
  AOI22_X1  g172(.A1(new_n364_), .A2(new_n366_), .B1(new_n369_), .B2(new_n371_), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT89), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(KEYINPUT89), .B1(new_n367_), .B2(new_n372_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n378_), .A2(new_n321_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n367_), .A2(new_n372_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G127gat), .B(G134gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G113gat), .B(G120gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n380_), .A2(new_n383_), .ZN(new_n384_));
  AND3_X1   g183(.A1(new_n332_), .A2(new_n333_), .A3(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(KEYINPUT4), .B1(new_n379_), .B2(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n376_), .B1(new_n384_), .B2(KEYINPUT89), .ZN(new_n387_));
  AOI21_X1  g186(.A(KEYINPUT4), .B1(new_n334_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n362_), .B1(new_n386_), .B2(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n332_), .A2(new_n333_), .A3(new_n384_), .ZN(new_n391_));
  OAI211_X1 g190(.A(new_n391_), .B(new_n362_), .C1(new_n321_), .C2(new_n378_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT100), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n334_), .A2(new_n387_), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n395_), .A2(KEYINPUT100), .A3(new_n362_), .A4(new_n391_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n394_), .A2(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n361_), .B1(new_n390_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n362_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT4), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n400_), .B1(new_n395_), .B2(new_n391_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n399_), .B1(new_n401_), .B2(new_n388_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n361_), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n402_), .A2(new_n403_), .A3(new_n394_), .A4(new_n396_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n398_), .A2(new_n404_), .A3(KEYINPUT103), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT103), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n406_), .B(new_n361_), .C1(new_n390_), .C2(new_n397_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n405_), .A2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n295_), .A2(new_n356_), .A3(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n232_), .A2(KEYINPUT30), .A3(new_n255_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(KEYINPUT30), .B1(new_n232_), .B2(new_n255_), .ZN(new_n412_));
  NOR3_X1   g211(.A1(new_n411_), .A2(KEYINPUT87), .A3(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n387_), .B(KEYINPUT31), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT88), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT87), .ZN(new_n418_));
  INV_X1    g217(.A(new_n412_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n418_), .B1(new_n419_), .B2(new_n410_), .ZN(new_n420_));
  XOR2_X1   g219(.A(G71gat), .B(G99gat), .Z(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(G43gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G227gat), .A2(G233gat), .ZN(new_n423_));
  INV_X1    g222(.A(G15gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  XOR2_X1   g224(.A(new_n422_), .B(new_n425_), .Z(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n417_), .B1(new_n420_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT90), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT87), .B1(new_n411_), .B2(new_n412_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n378_), .B(KEYINPUT31), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT88), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n430_), .A2(new_n432_), .A3(new_n426_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n428_), .A2(new_n429_), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n429_), .B1(new_n428_), .B2(new_n433_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n414_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  NOR3_X1   g236(.A1(new_n420_), .A2(new_n417_), .A3(new_n427_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n432_), .B1(new_n430_), .B2(new_n426_), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT90), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n440_), .A2(new_n413_), .A3(new_n434_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n437_), .A2(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n409_), .A2(new_n442_), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n437_), .A2(new_n441_), .A3(KEYINPUT91), .ZN(new_n444_));
  AOI21_X1  g243(.A(KEYINPUT91), .B1(new_n437_), .B2(new_n441_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n292_), .A2(new_n355_), .A3(new_n408_), .A4(new_n294_), .ZN(new_n447_));
  AND2_X1   g246(.A1(new_n281_), .A2(KEYINPUT32), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n448_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n281_), .A2(KEYINPUT32), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n271_), .A2(new_n276_), .A3(new_n450_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n449_), .A2(new_n407_), .A3(new_n405_), .A4(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n282_), .A2(new_n293_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n362_), .B1(new_n401_), .B2(new_n388_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n395_), .A2(new_n399_), .A3(new_n391_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n455_), .A2(KEYINPUT101), .A3(new_n361_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n454_), .A2(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(KEYINPUT101), .B1(new_n455_), .B2(new_n361_), .ZN(new_n458_));
  OR2_X1    g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n390_), .A2(new_n397_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n460_), .A2(KEYINPUT33), .A3(new_n403_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT33), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n404_), .A2(new_n462_), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n453_), .A2(new_n459_), .A3(new_n461_), .A4(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n355_), .B1(new_n452_), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT104), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n447_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  AOI211_X1 g266(.A(KEYINPUT104), .B(new_n355_), .C1(new_n452_), .C2(new_n464_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n446_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT105), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT105), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n446_), .B(new_n471_), .C1(new_n467_), .C2(new_n468_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n443_), .B1(new_n470_), .B2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT6), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(KEYINPUT66), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT66), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT6), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n475_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G99gat), .A2(G106gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT7), .ZN(new_n481_));
  INV_X1    g280(.A(G99gat), .ZN(new_n482_));
  INV_X1    g281(.A(G106gat), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n481_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n485_));
  AND2_X1   g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n475_), .A2(new_n477_), .A3(G99gat), .A4(G106gat), .ZN(new_n487_));
  AND3_X1   g286(.A1(new_n480_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  XOR2_X1   g287(.A(G85gat), .B(G92gat), .Z(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT8), .B1(new_n488_), .B2(new_n490_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n480_), .A2(new_n487_), .A3(new_n485_), .A4(new_n484_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT8), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n492_), .A2(new_n493_), .A3(new_n489_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT64), .ZN(new_n495_));
  INV_X1    g294(.A(G92gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(KEYINPUT64), .A2(G92gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(G85gat), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT9), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n500_), .A2(KEYINPUT65), .A3(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT65), .ZN(new_n503_));
  INV_X1    g302(.A(G85gat), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n504_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n503_), .B1(new_n505_), .B2(KEYINPUT9), .ZN(new_n506_));
  NOR3_X1   g305(.A1(new_n501_), .A2(new_n504_), .A3(new_n496_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n507_), .B1(new_n504_), .B2(new_n496_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n502_), .A2(new_n506_), .A3(new_n508_), .ZN(new_n509_));
  OR2_X1    g308(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n510_), .A2(new_n483_), .A3(new_n511_), .ZN(new_n512_));
  AND3_X1   g311(.A1(new_n480_), .A2(new_n512_), .A3(new_n487_), .ZN(new_n513_));
  AOI22_X1  g312(.A1(new_n491_), .A2(new_n494_), .B1(new_n509_), .B2(new_n513_), .ZN(new_n514_));
  XOR2_X1   g313(.A(G29gat), .B(G36gat), .Z(new_n515_));
  XOR2_X1   g314(.A(G43gat), .B(G50gat), .Z(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n514_), .A2(KEYINPUT71), .A3(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n509_), .A2(new_n513_), .ZN(new_n519_));
  AND3_X1   g318(.A1(new_n492_), .A2(new_n493_), .A3(new_n489_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n493_), .B1(new_n492_), .B2(new_n489_), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n519_), .B(new_n517_), .C1(new_n520_), .C2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT71), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n518_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT70), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n519_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n517_), .B(KEYINPUT15), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT35), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G232gat), .A2(G233gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT34), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  AOI22_X1  g331(.A1(new_n527_), .A2(new_n528_), .B1(new_n529_), .B2(new_n532_), .ZN(new_n533_));
  AND3_X1   g332(.A1(new_n525_), .A2(new_n526_), .A3(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n526_), .B1(new_n525_), .B2(new_n533_), .ZN(new_n535_));
  OAI22_X1  g334(.A1(new_n534_), .A2(new_n535_), .B1(new_n529_), .B2(new_n532_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n525_), .A2(new_n533_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT70), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n532_), .A2(new_n529_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n525_), .A2(new_n526_), .A3(new_n533_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n538_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n536_), .A2(new_n541_), .ZN(new_n542_));
  XOR2_X1   g341(.A(G190gat), .B(G218gat), .Z(new_n543_));
  XNOR2_X1  g342(.A(G134gat), .B(G162gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT36), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  XOR2_X1   g346(.A(new_n547_), .B(KEYINPUT72), .Z(new_n548_));
  NAND2_X1  g347(.A1(new_n542_), .A2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n545_), .B(KEYINPUT36), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n536_), .A2(new_n541_), .A3(new_n550_), .ZN(new_n551_));
  AND3_X1   g350(.A1(new_n549_), .A2(KEYINPUT107), .A3(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(KEYINPUT107), .B1(new_n549_), .B2(new_n551_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n473_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  XOR2_X1   g356(.A(G1gat), .B(G8gat), .Z(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(KEYINPUT76), .B(G1gat), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(G8gat), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(KEYINPUT14), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT77), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT14), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n565_), .B1(new_n560_), .B2(G8gat), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(KEYINPUT77), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n564_), .A2(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(G15gat), .B(G22gat), .Z(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n559_), .B1(new_n568_), .B2(new_n570_), .ZN(new_n571_));
  AOI211_X1 g370(.A(new_n569_), .B(new_n558_), .C1(new_n564_), .C2(new_n567_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(G231gat), .A2(G233gat), .ZN(new_n574_));
  XOR2_X1   g373(.A(new_n574_), .B(KEYINPUT78), .Z(new_n575_));
  XNOR2_X1  g374(.A(new_n573_), .B(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G57gat), .B(G64gat), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(KEYINPUT11), .ZN(new_n578_));
  XOR2_X1   g377(.A(G71gat), .B(G78gat), .Z(new_n579_));
  AND2_X1   g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n580_), .B1(KEYINPUT11), .B2(new_n577_), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n578_), .A2(new_n579_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n576_), .B(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(G127gat), .B(G155gat), .Z(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT16), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G183gat), .B(G211gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT17), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n588_), .A2(new_n589_), .ZN(new_n591_));
  OR3_X1    g390(.A1(new_n584_), .A2(new_n590_), .A3(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT79), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n593_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n584_), .A2(new_n590_), .ZN(new_n596_));
  AND3_X1   g395(.A1(new_n594_), .A2(new_n595_), .A3(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(G230gat), .A2(G233gat), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  OAI211_X1 g398(.A(new_n583_), .B(new_n519_), .C1(new_n520_), .C2(new_n521_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n514_), .A2(new_n583_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n599_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT67), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n600_), .A2(new_n604_), .A3(new_n598_), .ZN(new_n605_));
  NOR3_X1   g404(.A1(new_n514_), .A2(KEYINPUT12), .A3(new_n583_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT12), .ZN(new_n607_));
  INV_X1    g406(.A(new_n583_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n607_), .B1(new_n527_), .B2(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n605_), .B1(new_n606_), .B2(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n599_), .B1(new_n514_), .B2(new_n583_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n611_), .A2(new_n604_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n603_), .B1(new_n610_), .B2(new_n612_), .ZN(new_n613_));
  XOR2_X1   g412(.A(KEYINPUT68), .B(KEYINPUT5), .Z(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT69), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G120gat), .B(G148gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G176gat), .B(G204gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n613_), .B(new_n620_), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n621_), .A2(KEYINPUT13), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(KEYINPUT13), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n517_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n567_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n566_), .A2(KEYINPUT77), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n570_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(new_n558_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n517_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n568_), .A2(new_n570_), .A3(new_n559_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n629_), .A2(new_n630_), .A3(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n625_), .A2(new_n632_), .A3(KEYINPUT80), .ZN(new_n633_));
  NAND2_X1  g432(.A1(G229gat), .A2(G233gat), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT80), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n573_), .A2(new_n636_), .A3(new_n630_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n633_), .A2(new_n635_), .A3(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n573_), .A2(new_n528_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n639_), .A2(new_n634_), .A3(new_n625_), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n638_), .A2(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(G113gat), .B(G141gat), .ZN(new_n642_));
  XNOR2_X1  g441(.A(G169gat), .B(G197gat), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n642_), .B(new_n643_), .Z(new_n644_));
  OR2_X1    g443(.A1(new_n641_), .A2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n638_), .A2(new_n640_), .A3(new_n644_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT81), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n638_), .A2(new_n640_), .A3(KEYINPUT81), .A4(new_n644_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n645_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n624_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n597_), .A2(new_n653_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n557_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(G1gat), .B1(new_n656_), .B2(new_n408_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT38), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n473_), .A2(new_n652_), .ZN(new_n659_));
  XOR2_X1   g458(.A(new_n550_), .B(KEYINPUT73), .Z(new_n660_));
  NAND3_X1  g459(.A1(new_n536_), .A2(new_n541_), .A3(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n549_), .A2(KEYINPUT74), .A3(new_n661_), .ZN(new_n662_));
  OAI211_X1 g461(.A(new_n662_), .B(KEYINPUT37), .C1(KEYINPUT74), .C2(new_n661_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT75), .ZN(new_n664_));
  INV_X1    g463(.A(new_n551_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n548_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n666_), .B1(new_n536_), .B2(new_n541_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n665_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT37), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n664_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n549_), .A2(new_n669_), .A3(new_n551_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n671_), .A2(KEYINPUT75), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n663_), .B1(new_n670_), .B2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(new_n597_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n674_), .A2(new_n624_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n408_), .A2(new_n560_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n659_), .A2(new_n675_), .A3(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT106), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n677_), .B(new_n678_), .ZN(new_n679_));
  AND3_X1   g478(.A1(new_n679_), .A2(KEYINPUT108), .A3(new_n658_), .ZN(new_n680_));
  AOI21_X1  g479(.A(KEYINPUT108), .B1(new_n679_), .B2(new_n658_), .ZN(new_n681_));
  OAI221_X1 g480(.A(new_n657_), .B1(new_n658_), .B2(new_n679_), .C1(new_n680_), .C2(new_n681_), .ZN(G1324gat));
  AND2_X1   g481(.A1(new_n659_), .A2(new_n675_), .ZN(new_n683_));
  INV_X1    g482(.A(G8gat), .ZN(new_n684_));
  INV_X1    g483(.A(new_n295_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n683_), .A2(new_n684_), .A3(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT39), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT109), .ZN(new_n688_));
  INV_X1    g487(.A(new_n654_), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n556_), .A2(new_n688_), .A3(new_n685_), .A4(new_n689_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n690_), .A2(G8gat), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n556_), .A2(new_n685_), .A3(new_n689_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(KEYINPUT109), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n687_), .B1(new_n691_), .B2(new_n693_), .ZN(new_n694_));
  AND4_X1   g493(.A1(new_n687_), .A2(new_n693_), .A3(new_n690_), .A4(G8gat), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n686_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT40), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  OAI211_X1 g497(.A(KEYINPUT40), .B(new_n686_), .C1(new_n694_), .C2(new_n695_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1325gat));
  INV_X1    g499(.A(new_n446_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n424_), .B1(new_n655_), .B2(new_n701_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT41), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n683_), .A2(new_n424_), .A3(new_n701_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(G1326gat));
  INV_X1    g504(.A(G22gat), .ZN(new_n706_));
  XOR2_X1   g505(.A(new_n355_), .B(KEYINPUT110), .Z(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n683_), .A2(new_n706_), .A3(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n655_), .A2(new_n708_), .ZN(new_n710_));
  XOR2_X1   g509(.A(KEYINPUT111), .B(KEYINPUT42), .Z(new_n711_));
  AND3_X1   g510(.A1(new_n710_), .A2(G22gat), .A3(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n711_), .B1(new_n710_), .B2(G22gat), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n709_), .B1(new_n712_), .B2(new_n713_), .ZN(G1327gat));
  INV_X1    g513(.A(new_n443_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n452_), .A2(new_n464_), .ZN(new_n716_));
  OAI21_X1  g515(.A(KEYINPUT104), .B1(new_n716_), .B2(new_n355_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n465_), .A2(new_n466_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n717_), .A2(new_n718_), .A3(new_n447_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n471_), .B1(new_n719_), .B2(new_n446_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n472_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n715_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n624_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n597_), .A2(new_n554_), .ZN(new_n724_));
  AND4_X1   g523(.A1(new_n651_), .A2(new_n722_), .A3(new_n723_), .A4(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n408_), .ZN(new_n726_));
  AOI21_X1  g525(.A(G29gat), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n673_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT43), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n729_), .A2(KEYINPUT112), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n722_), .A2(new_n728_), .A3(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(KEYINPUT112), .B(KEYINPUT43), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n734_), .B1(new_n473_), .B2(new_n673_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n732_), .A2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n597_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(new_n653_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(KEYINPUT44), .B1(new_n736_), .B2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT44), .ZN(new_n741_));
  AOI211_X1 g540(.A(new_n741_), .B(new_n738_), .C1(new_n732_), .C2(new_n735_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n740_), .A2(new_n742_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n726_), .A2(G29gat), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n727_), .B1(new_n743_), .B2(new_n744_), .ZN(G1328gat));
  XNOR2_X1  g544(.A(KEYINPUT114), .B(KEYINPUT46), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(G36gat), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n748_), .B1(new_n743_), .B2(new_n685_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n725_), .A2(new_n748_), .A3(new_n685_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(KEYINPUT113), .B(KEYINPUT45), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n750_), .B(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n747_), .B1(new_n749_), .B2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n751_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n750_), .B(new_n754_), .ZN(new_n755_));
  NOR3_X1   g554(.A1(new_n740_), .A2(new_n742_), .A3(new_n295_), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n755_), .B(new_n746_), .C1(new_n756_), .C2(new_n748_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n753_), .A2(new_n757_), .ZN(G1329gat));
  INV_X1    g557(.A(new_n442_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(G43gat), .ZN(new_n760_));
  NOR3_X1   g559(.A1(new_n740_), .A2(new_n742_), .A3(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(G43gat), .B1(new_n725_), .B2(new_n701_), .ZN(new_n762_));
  OR3_X1    g561(.A1(new_n761_), .A2(KEYINPUT47), .A3(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(KEYINPUT47), .B1(new_n761_), .B2(new_n762_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(G1330gat));
  INV_X1    g564(.A(G50gat), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n725_), .A2(new_n766_), .A3(new_n708_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n743_), .A2(KEYINPUT115), .A3(new_n355_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(G50gat), .ZN(new_n769_));
  AOI21_X1  g568(.A(KEYINPUT115), .B1(new_n743_), .B2(new_n355_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n767_), .B1(new_n769_), .B2(new_n770_), .ZN(G1331gat));
  NOR4_X1   g570(.A1(new_n473_), .A2(new_n674_), .A3(new_n651_), .A4(new_n723_), .ZN(new_n772_));
  INV_X1    g571(.A(G57gat), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n772_), .A2(new_n773_), .A3(new_n726_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n723_), .A2(new_n651_), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n556_), .A2(new_n597_), .A3(new_n775_), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n776_), .A2(new_n726_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n774_), .B1(new_n777_), .B2(new_n773_), .ZN(G1332gat));
  INV_X1    g577(.A(G64gat), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n779_), .B1(new_n776_), .B2(new_n685_), .ZN(new_n780_));
  XOR2_X1   g579(.A(new_n780_), .B(KEYINPUT48), .Z(new_n781_));
  NAND3_X1  g580(.A1(new_n772_), .A2(new_n779_), .A3(new_n685_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(G1333gat));
  INV_X1    g582(.A(G71gat), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n784_), .B1(new_n776_), .B2(new_n701_), .ZN(new_n785_));
  XOR2_X1   g584(.A(new_n785_), .B(KEYINPUT49), .Z(new_n786_));
  NAND3_X1  g585(.A1(new_n772_), .A2(new_n784_), .A3(new_n701_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(G1334gat));
  INV_X1    g587(.A(G78gat), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n789_), .B1(new_n776_), .B2(new_n708_), .ZN(new_n790_));
  XOR2_X1   g589(.A(new_n790_), .B(KEYINPUT50), .Z(new_n791_));
  NAND3_X1  g590(.A1(new_n772_), .A2(new_n789_), .A3(new_n708_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(G1335gat));
  NOR3_X1   g592(.A1(new_n473_), .A2(new_n651_), .A3(new_n723_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(new_n724_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n796_), .A2(new_n504_), .A3(new_n726_), .ZN(new_n797_));
  AND3_X1   g596(.A1(new_n736_), .A2(new_n737_), .A3(new_n775_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n798_), .A2(new_n726_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n797_), .B1(new_n799_), .B2(new_n504_), .ZN(G1336gat));
  AOI21_X1  g599(.A(G92gat), .B1(new_n796_), .B2(new_n685_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n685_), .A2(new_n499_), .ZN(new_n802_));
  XOR2_X1   g601(.A(new_n802_), .B(KEYINPUT116), .Z(new_n803_));
  AOI21_X1  g602(.A(new_n801_), .B1(new_n798_), .B2(new_n803_), .ZN(G1337gat));
  AOI21_X1  g603(.A(new_n482_), .B1(new_n798_), .B2(new_n701_), .ZN(new_n805_));
  AND4_X1   g604(.A1(new_n759_), .A2(new_n796_), .A3(new_n510_), .A4(new_n511_), .ZN(new_n806_));
  OR3_X1    g605(.A1(new_n805_), .A2(new_n806_), .A3(KEYINPUT51), .ZN(new_n807_));
  OAI21_X1  g606(.A(KEYINPUT51), .B1(new_n805_), .B2(new_n806_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(G1338gat));
  NAND3_X1  g608(.A1(new_n796_), .A2(new_n483_), .A3(new_n355_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n736_), .A2(new_n355_), .A3(new_n737_), .A4(new_n775_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT52), .ZN(new_n812_));
  AND3_X1   g611(.A1(new_n811_), .A2(new_n812_), .A3(G106gat), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n812_), .B1(new_n811_), .B2(G106gat), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n810_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n817_), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n810_), .B(new_n816_), .C1(new_n813_), .C2(new_n814_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(G1339gat));
  OAI21_X1  g619(.A(KEYINPUT12), .B1(new_n514_), .B2(new_n583_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n527_), .A2(new_n607_), .A3(new_n608_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n598_), .B1(new_n823_), .B2(new_n600_), .ZN(new_n824_));
  OAI21_X1  g623(.A(KEYINPUT55), .B1(new_n610_), .B2(new_n612_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n600_), .A2(new_n598_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(KEYINPUT67), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT55), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n827_), .A2(new_n823_), .A3(new_n828_), .A4(new_n605_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n824_), .B1(new_n825_), .B2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT118), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n620_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n824_), .ZN(new_n833_));
  AOI22_X1  g632(.A1(new_n821_), .A2(new_n822_), .B1(new_n611_), .B2(new_n604_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n828_), .B1(new_n834_), .B2(new_n827_), .ZN(new_n835_));
  AND4_X1   g634(.A1(new_n828_), .A2(new_n827_), .A3(new_n823_), .A4(new_n605_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n833_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(KEYINPUT118), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n832_), .A2(new_n838_), .A3(KEYINPUT56), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(KEYINPUT119), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT119), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n832_), .A2(new_n838_), .A3(new_n841_), .A4(KEYINPUT56), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT56), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n831_), .B(new_n833_), .C1(new_n835_), .C2(new_n836_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n619_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n830_), .A2(new_n831_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n843_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n840_), .A2(new_n842_), .A3(new_n847_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n633_), .A2(new_n634_), .A3(new_n637_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n625_), .A2(new_n635_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n644_), .B1(new_n850_), .B2(new_n639_), .ZN(new_n851_));
  AOI22_X1  g650(.A1(new_n648_), .A2(new_n649_), .B1(new_n849_), .B2(new_n851_), .ZN(new_n852_));
  OR2_X1    g651(.A1(new_n613_), .A2(new_n619_), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n848_), .A2(KEYINPUT58), .A3(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(KEYINPUT58), .B1(new_n848_), .B2(new_n854_), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n855_), .A2(new_n856_), .A3(new_n673_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n651_), .A2(new_n853_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n858_), .B1(new_n847_), .B2(new_n839_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n621_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n852_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n554_), .B1(new_n859_), .B2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  OAI211_X1 g664(.A(KEYINPUT57), .B(new_n554_), .C1(new_n859_), .C2(new_n862_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n737_), .B1(new_n857_), .B2(new_n867_), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n673_), .A2(new_n652_), .A3(new_n597_), .A4(new_n723_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(KEYINPUT54), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n868_), .A2(new_n870_), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n685_), .A2(new_n408_), .A3(new_n442_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n871_), .A2(new_n356_), .A3(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n874_), .A2(new_n370_), .A3(new_n651_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT120), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n873_), .B1(new_n876_), .B2(KEYINPUT59), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n355_), .B1(new_n868_), .B2(new_n870_), .ZN(new_n878_));
  XOR2_X1   g677(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n879_));
  NAND3_X1  g678(.A1(new_n878_), .A2(new_n872_), .A3(new_n879_), .ZN(new_n880_));
  AND3_X1   g679(.A1(new_n877_), .A2(new_n651_), .A3(new_n880_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n875_), .B1(new_n881_), .B2(new_n370_), .ZN(G1340gat));
  OAI21_X1  g681(.A(new_n368_), .B1(new_n723_), .B2(KEYINPUT60), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n874_), .B(new_n883_), .C1(KEYINPUT60), .C2(new_n368_), .ZN(new_n884_));
  AND3_X1   g683(.A1(new_n877_), .A2(new_n624_), .A3(new_n880_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n885_), .B2(new_n368_), .ZN(G1341gat));
  AND2_X1   g685(.A1(new_n878_), .A2(new_n597_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n887_), .A2(new_n365_), .A3(new_n872_), .ZN(new_n888_));
  AND3_X1   g687(.A1(new_n877_), .A2(new_n597_), .A3(new_n880_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n889_), .B2(new_n365_), .ZN(G1342gat));
  NAND3_X1  g689(.A1(new_n874_), .A2(new_n363_), .A3(new_n555_), .ZN(new_n891_));
  AND3_X1   g690(.A1(new_n877_), .A2(new_n728_), .A3(new_n880_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n892_), .B2(new_n363_), .ZN(G1343gat));
  NOR3_X1   g692(.A1(new_n685_), .A2(new_n356_), .A3(new_n408_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n871_), .A2(new_n446_), .A3(new_n894_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n895_), .A2(new_n652_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(new_n303_), .ZN(G1344gat));
  NOR2_X1   g696(.A1(new_n895_), .A2(new_n723_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(new_n304_), .ZN(G1345gat));
  OAI21_X1  g698(.A(KEYINPUT121), .B1(new_n895_), .B2(new_n737_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n701_), .B1(new_n868_), .B2(new_n870_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT121), .ZN(new_n902_));
  NAND4_X1  g701(.A1(new_n901_), .A2(new_n902_), .A3(new_n597_), .A4(new_n894_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(KEYINPUT61), .B(G155gat), .ZN(new_n904_));
  AND3_X1   g703(.A1(new_n900_), .A2(new_n903_), .A3(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n904_), .B1(new_n900_), .B2(new_n903_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n905_), .A2(new_n906_), .ZN(G1346gat));
  OAI21_X1  g706(.A(G162gat), .B1(new_n895_), .B2(new_n673_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n555_), .A2(new_n312_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n895_), .B2(new_n909_), .ZN(G1347gat));
  NOR3_X1   g709(.A1(new_n446_), .A2(new_n726_), .A3(new_n295_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n707_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n912_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n871_), .A2(new_n651_), .A3(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(G169gat), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(KEYINPUT122), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT122), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n914_), .A2(new_n917_), .A3(G169gat), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n916_), .A2(KEYINPUT62), .A3(new_n918_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n912_), .B1(new_n868_), .B2(new_n870_), .ZN(new_n921_));
  AOI211_X1 g720(.A(KEYINPUT122), .B(new_n218_), .C1(new_n921_), .C2(new_n651_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n917_), .B1(new_n914_), .B2(G169gat), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n920_), .B1(new_n922_), .B2(new_n923_), .ZN(new_n924_));
  OR2_X1    g723(.A1(new_n914_), .A2(new_n268_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n919_), .A2(new_n924_), .A3(new_n925_), .ZN(G1348gat));
  AOI21_X1  g725(.A(G176gat), .B1(new_n921_), .B2(new_n624_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n911_), .A2(G176gat), .A3(new_n624_), .ZN(new_n928_));
  INV_X1    g727(.A(new_n928_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n927_), .B1(new_n878_), .B2(new_n929_), .ZN(G1349gat));
  AOI21_X1  g729(.A(G183gat), .B1(new_n887_), .B2(new_n911_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n737_), .A2(new_n215_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n931_), .B1(new_n921_), .B2(new_n932_), .ZN(G1350gat));
  NAND3_X1  g732(.A1(new_n921_), .A2(new_n264_), .A3(new_n555_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n921_), .A2(new_n728_), .ZN(new_n935_));
  AND3_X1   g734(.A1(new_n935_), .A2(KEYINPUT123), .A3(G190gat), .ZN(new_n936_));
  AOI21_X1  g735(.A(KEYINPUT123), .B1(new_n935_), .B2(G190gat), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n934_), .B1(new_n936_), .B2(new_n937_), .ZN(G1351gat));
  NOR3_X1   g737(.A1(new_n295_), .A2(new_n356_), .A3(new_n726_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n901_), .A2(new_n651_), .A3(new_n939_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n940_), .B1(KEYINPUT124), .B2(new_n233_), .ZN(new_n941_));
  XOR2_X1   g740(.A(KEYINPUT124), .B(G197gat), .Z(new_n942_));
  AOI21_X1  g741(.A(new_n941_), .B1(new_n940_), .B2(new_n942_), .ZN(G1352gat));
  NAND4_X1  g742(.A1(new_n871_), .A2(new_n446_), .A3(new_n624_), .A4(new_n939_), .ZN(new_n944_));
  OAI21_X1  g743(.A(KEYINPUT126), .B1(new_n944_), .B2(G204gat), .ZN(new_n945_));
  INV_X1    g744(.A(KEYINPUT125), .ZN(new_n946_));
  NAND4_X1  g745(.A1(new_n901_), .A2(new_n946_), .A3(new_n624_), .A4(new_n939_), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n234_), .B1(new_n944_), .B2(KEYINPUT125), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n945_), .B1(new_n947_), .B2(new_n948_), .ZN(new_n949_));
  INV_X1    g748(.A(KEYINPUT126), .ZN(new_n950_));
  INV_X1    g749(.A(new_n858_), .ZN(new_n951_));
  NOR3_X1   g750(.A1(new_n845_), .A2(new_n846_), .A3(new_n843_), .ZN(new_n952_));
  AOI21_X1  g751(.A(KEYINPUT56), .B1(new_n832_), .B2(new_n838_), .ZN(new_n953_));
  OAI21_X1  g752(.A(new_n951_), .B1(new_n952_), .B2(new_n953_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n954_), .A2(new_n861_), .ZN(new_n955_));
  AOI21_X1  g754(.A(KEYINPUT57), .B1(new_n955_), .B2(new_n554_), .ZN(new_n956_));
  INV_X1    g755(.A(new_n866_), .ZN(new_n957_));
  NOR2_X1   g756(.A1(new_n956_), .A2(new_n957_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n848_), .A2(new_n854_), .ZN(new_n959_));
  INV_X1    g758(.A(KEYINPUT58), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n959_), .A2(new_n960_), .ZN(new_n961_));
  NAND3_X1  g760(.A1(new_n848_), .A2(KEYINPUT58), .A3(new_n854_), .ZN(new_n962_));
  NAND3_X1  g761(.A1(new_n961_), .A2(new_n728_), .A3(new_n962_), .ZN(new_n963_));
  AOI21_X1  g762(.A(new_n597_), .B1(new_n958_), .B2(new_n963_), .ZN(new_n964_));
  INV_X1    g763(.A(KEYINPUT54), .ZN(new_n965_));
  XNOR2_X1  g764(.A(new_n869_), .B(new_n965_), .ZN(new_n966_));
  OAI211_X1 g765(.A(new_n446_), .B(new_n939_), .C1(new_n964_), .C2(new_n966_), .ZN(new_n967_));
  OAI21_X1  g766(.A(KEYINPUT125), .B1(new_n967_), .B2(new_n723_), .ZN(new_n968_));
  AND4_X1   g767(.A1(new_n950_), .A2(new_n968_), .A3(G204gat), .A4(new_n947_), .ZN(new_n969_));
  NOR2_X1   g768(.A1(new_n949_), .A2(new_n969_), .ZN(G1353gat));
  NOR2_X1   g769(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n971_));
  AND2_X1   g770(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n972_));
  NOR4_X1   g771(.A1(new_n967_), .A2(new_n737_), .A3(new_n971_), .A4(new_n972_), .ZN(new_n973_));
  OAI21_X1  g772(.A(new_n971_), .B1(new_n967_), .B2(new_n737_), .ZN(new_n974_));
  OR2_X1    g773(.A1(new_n974_), .A2(KEYINPUT127), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n974_), .A2(KEYINPUT127), .ZN(new_n976_));
  AOI21_X1  g775(.A(new_n973_), .B1(new_n975_), .B2(new_n976_), .ZN(G1354gat));
  OAI21_X1  g776(.A(G218gat), .B1(new_n967_), .B2(new_n673_), .ZN(new_n978_));
  OR2_X1    g777(.A1(new_n554_), .A2(G218gat), .ZN(new_n979_));
  OAI21_X1  g778(.A(new_n978_), .B1(new_n967_), .B2(new_n979_), .ZN(G1355gat));
endmodule


