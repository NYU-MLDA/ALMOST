//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 1 1 0 0 1 0 0 0 0 1 0 1 0 0 1 0 1 0 1 0 0 0 1 0 1 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n610_, new_n611_,
    new_n612_, new_n614_, new_n615_, new_n616_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n675_, new_n676_, new_n677_, new_n679_,
    new_n680_, new_n681_, new_n683_, new_n684_, new_n685_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n699_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n825_, new_n826_, new_n827_, new_n829_,
    new_n830_, new_n832_, new_n833_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n852_, new_n853_, new_n854_, new_n856_, new_n857_, new_n858_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_;
  XOR2_X1   g000(.A(G127gat), .B(G134gat), .Z(new_n202_));
  XOR2_X1   g001(.A(G113gat), .B(G120gat), .Z(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G127gat), .B(G134gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G113gat), .B(G120gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n204_), .A2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT31), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G227gat), .A2(G233gat), .ZN(new_n210_));
  XOR2_X1   g009(.A(new_n210_), .B(G15gat), .Z(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(G71gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(G99gat), .ZN(new_n213_));
  XOR2_X1   g012(.A(KEYINPUT79), .B(KEYINPUT30), .Z(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  NOR3_X1   g014(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G183gat), .A2(G190gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n218_), .B(KEYINPUT76), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT23), .ZN(new_n220_));
  AND2_X1   g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n220_), .B1(G183gat), .B2(G190gat), .ZN(new_n222_));
  OAI211_X1 g021(.A(KEYINPUT77), .B(new_n217_), .C1(new_n221_), .C2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT77), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n222_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n224_), .B1(new_n225_), .B2(new_n216_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(KEYINPUT75), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(KEYINPUT25), .B(G183gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT26), .B(G190gat), .ZN(new_n232_));
  AOI22_X1  g031(.A1(new_n228_), .A2(new_n230_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n223_), .A2(new_n226_), .A3(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n235_), .B1(new_n219_), .B2(KEYINPUT23), .ZN(new_n236_));
  NOR2_X1   g035(.A1(G183gat), .A2(G190gat), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n236_), .A2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(KEYINPUT22), .B(G169gat), .ZN(new_n240_));
  INV_X1    g039(.A(G176gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(new_n228_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT78), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n242_), .A2(new_n228_), .A3(KEYINPUT78), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n239_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n234_), .A2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT80), .B(G43gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  OR2_X1    g049(.A1(new_n215_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n215_), .A2(new_n250_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n209_), .B1(new_n253_), .B2(KEYINPUT81), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT81), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n251_), .A2(new_n255_), .A3(new_n252_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n254_), .A2(new_n256_), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n251_), .A2(new_n255_), .A3(new_n252_), .A4(new_n209_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT21), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G197gat), .B(G204gat), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT84), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G211gat), .B(G218gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n264_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(new_n261_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n260_), .B1(new_n265_), .B2(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(KEYINPUT21), .B1(new_n263_), .B2(new_n264_), .ZN(new_n269_));
  OR2_X1    g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n230_), .A2(new_n227_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n216_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n236_), .A2(new_n272_), .A3(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT86), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT87), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n228_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n228_), .A2(new_n276_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n277_), .A2(new_n278_), .A3(new_n242_), .ZN(new_n279_));
  OAI211_X1 g078(.A(KEYINPUT88), .B(new_n238_), .C1(new_n221_), .C2(new_n222_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT88), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n281_), .B1(new_n225_), .B2(new_n237_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n279_), .B1(new_n280_), .B2(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n271_), .B1(new_n275_), .B2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n234_), .A2(new_n270_), .A3(new_n247_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n284_), .A2(KEYINPUT20), .A3(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G226gat), .A2(G233gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT19), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n270_), .B1(new_n234_), .B2(new_n247_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n288_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT20), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n275_), .A2(new_n283_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n293_), .B1(new_n294_), .B2(new_n271_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n289_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G64gat), .B(G92gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT90), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G8gat), .B(G36gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n296_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT27), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n289_), .A2(new_n295_), .A3(new_n302_), .ZN(new_n306_));
  AND3_X1   g105(.A1(new_n304_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT96), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n289_), .A2(new_n295_), .A3(KEYINPUT96), .A4(new_n302_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT95), .B(KEYINPUT20), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n270_), .A2(new_n274_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n311_), .B1(new_n312_), .B2(new_n283_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n288_), .B1(new_n313_), .B2(new_n290_), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n284_), .A2(KEYINPUT20), .A3(new_n285_), .A4(new_n291_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(new_n303_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n309_), .A2(new_n310_), .A3(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n307_), .B1(KEYINPUT27), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(G155gat), .ZN(new_n320_));
  INV_X1    g119(.A(G162gat), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n320_), .A2(new_n321_), .A3(KEYINPUT82), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G155gat), .A2(G162gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT1), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT82), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n325_), .B1(G155gat), .B2(G162gat), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n322_), .A2(new_n324_), .A3(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT83), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n322_), .A2(new_n324_), .A3(new_n326_), .A4(KEYINPUT83), .ZN(new_n330_));
  OAI211_X1 g129(.A(new_n329_), .B(new_n330_), .C1(KEYINPUT1), .C2(new_n323_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G141gat), .A2(G148gat), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(G141gat), .A2(G148gat), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(KEYINPUT3), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n332_), .B(KEYINPUT2), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  AND3_X1   g137(.A1(new_n322_), .A2(new_n326_), .A3(new_n323_), .ZN(new_n339_));
  AOI22_X1  g138(.A1(new_n331_), .A2(new_n335_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n270_), .B1(new_n341_), .B2(KEYINPUT29), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G228gat), .A2(G233gat), .ZN(new_n343_));
  OR2_X1    g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n342_), .A2(new_n343_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G78gat), .B(G106gat), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n344_), .A2(new_n345_), .A3(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT85), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n341_), .A2(KEYINPUT29), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G22gat), .B(G50gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT28), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n351_), .B(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n345_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n342_), .A2(new_n343_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n346_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  AOI22_X1  g156(.A1(new_n350_), .A2(new_n354_), .B1(new_n357_), .B2(new_n348_), .ZN(new_n358_));
  AND4_X1   g157(.A1(KEYINPUT85), .A2(new_n357_), .A3(new_n348_), .A4(new_n354_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G1gat), .B(G29gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(G85gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT0), .B(G57gat), .ZN(new_n363_));
  XOR2_X1   g162(.A(new_n362_), .B(new_n363_), .Z(new_n364_));
  INV_X1    g163(.A(KEYINPUT91), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n208_), .B(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n366_), .A2(new_n340_), .A3(KEYINPUT92), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n366_), .A2(new_n340_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT92), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n369_), .B1(new_n340_), .B2(new_n208_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n367_), .B1(new_n368_), .B2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G225gat), .A2(G233gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT93), .ZN(new_n374_));
  OAI211_X1 g173(.A(KEYINPUT4), .B(new_n367_), .C1(new_n368_), .C2(new_n370_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT4), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n376_), .B1(new_n340_), .B2(new_n208_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n372_), .B1(new_n375_), .B2(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n374_), .A2(new_n378_), .ZN(new_n379_));
  AOI211_X1 g178(.A(KEYINPUT93), .B(new_n372_), .C1(new_n375_), .C2(new_n377_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n364_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT93), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n378_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n364_), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n383_), .B(new_n384_), .C1(new_n378_), .C2(new_n374_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n360_), .A2(new_n381_), .A3(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n319_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT33), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n381_), .A2(new_n388_), .ZN(new_n389_));
  OAI211_X1 g188(.A(KEYINPUT33), .B(new_n364_), .C1(new_n379_), .C2(new_n380_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n372_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n364_), .B1(new_n371_), .B2(new_n391_), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n375_), .A2(new_n377_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n392_), .B1(new_n393_), .B2(new_n391_), .ZN(new_n394_));
  AND3_X1   g193(.A1(new_n304_), .A2(new_n394_), .A3(new_n306_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n389_), .A2(new_n390_), .A3(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n381_), .A2(new_n385_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n302_), .A2(KEYINPUT32), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n316_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT94), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n399_), .B1(new_n400_), .B2(new_n296_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n398_), .B1(new_n296_), .B2(KEYINPUT94), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n397_), .A2(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n360_), .B1(new_n396_), .B2(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n259_), .B1(new_n387_), .B2(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n259_), .A2(new_n397_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n360_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n319_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n407_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n406_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G229gat), .A2(G233gat), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT73), .ZN(new_n414_));
  XOR2_X1   g213(.A(G15gat), .B(G22gat), .Z(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G1gat), .B(G8gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT72), .B(G1gat), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n418_), .A2(G8gat), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT14), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n416_), .B(new_n417_), .C1(new_n419_), .C2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n417_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n420_), .B1(new_n418_), .B2(G8gat), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n422_), .B1(new_n423_), .B2(new_n415_), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n421_), .A2(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G43gat), .B(G50gat), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G29gat), .B(G36gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(KEYINPUT69), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n428_), .A2(KEYINPUT69), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n427_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n431_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n433_), .A2(new_n429_), .A3(new_n426_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n432_), .A2(new_n434_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n414_), .B1(new_n425_), .B2(new_n435_), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n432_), .A2(new_n434_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n421_), .A2(new_n424_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n437_), .A2(KEYINPUT73), .A3(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n413_), .B1(new_n436_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT15), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n435_), .B(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(KEYINPUT74), .B1(new_n442_), .B2(new_n425_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n435_), .A2(new_n441_), .ZN(new_n444_));
  AOI21_X1  g243(.A(KEYINPUT15), .B1(new_n432_), .B2(new_n434_), .ZN(new_n445_));
  OAI211_X1 g244(.A(KEYINPUT74), .B(new_n425_), .C1(new_n444_), .C2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n440_), .B1(new_n443_), .B2(new_n447_), .ZN(new_n448_));
  NOR3_X1   g247(.A1(new_n425_), .A2(new_n414_), .A3(new_n435_), .ZN(new_n449_));
  AOI21_X1  g248(.A(KEYINPUT73), .B1(new_n437_), .B2(new_n438_), .ZN(new_n450_));
  OAI22_X1  g249(.A1(new_n449_), .A2(new_n450_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(new_n413_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G113gat), .B(G141gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G169gat), .B(G197gat), .ZN(new_n454_));
  XOR2_X1   g253(.A(new_n453_), .B(new_n454_), .Z(new_n455_));
  NAND3_X1  g254(.A1(new_n448_), .A2(new_n452_), .A3(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n455_), .B1(new_n448_), .B2(new_n452_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT13), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G230gat), .A2(G233gat), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(G85gat), .ZN(new_n464_));
  INV_X1    g263(.A(G92gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G85gat), .A2(G92gat), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT6), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n469_), .B1(G99gat), .B2(G106gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G99gat), .A2(G106gat), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n471_), .A2(KEYINPUT6), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n470_), .A2(new_n472_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(G99gat), .A2(G106gat), .ZN(new_n474_));
  NOR2_X1   g273(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  OAI22_X1  g275(.A1(KEYINPUT65), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n468_), .B1(new_n473_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT8), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n477_), .B(new_n476_), .C1(new_n470_), .C2(new_n472_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n482_), .A2(KEYINPUT8), .A3(new_n468_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n471_), .B(KEYINPUT6), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT9), .ZN(new_n485_));
  AND2_X1   g284(.A1(G85gat), .A2(G92gat), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n466_), .B(new_n485_), .C1(new_n486_), .C2(KEYINPUT64), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT64), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n466_), .A2(new_n488_), .A3(KEYINPUT9), .A4(new_n467_), .ZN(new_n489_));
  OR2_X1    g288(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n490_));
  INV_X1    g289(.A(G106gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n490_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n484_), .A2(new_n487_), .A3(new_n489_), .A4(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G57gat), .B(G64gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G71gat), .B(G78gat), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n495_), .A2(new_n496_), .A3(KEYINPUT11), .ZN(new_n497_));
  XOR2_X1   g296(.A(G71gat), .B(G78gat), .Z(new_n498_));
  INV_X1    g297(.A(G64gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(G57gat), .ZN(new_n500_));
  INV_X1    g299(.A(G57gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(G64gat), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n500_), .A2(new_n502_), .A3(KEYINPUT11), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n498_), .A2(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n495_), .A2(KEYINPUT11), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n497_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n481_), .A2(new_n483_), .A3(new_n494_), .A4(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT66), .ZN(new_n508_));
  AOI21_X1  g307(.A(KEYINPUT8), .B1(new_n482_), .B2(new_n468_), .ZN(new_n509_));
  AND4_X1   g308(.A1(new_n484_), .A2(new_n487_), .A3(new_n489_), .A4(new_n493_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT66), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n511_), .A2(new_n512_), .A3(new_n483_), .A4(new_n506_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n508_), .A2(new_n513_), .ZN(new_n514_));
  AND3_X1   g313(.A1(new_n482_), .A2(KEYINPUT8), .A3(new_n468_), .ZN(new_n515_));
  NOR3_X1   g314(.A1(new_n515_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n516_), .A2(new_n506_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n463_), .B1(new_n514_), .B2(new_n517_), .ZN(new_n518_));
  AND2_X1   g317(.A1(new_n507_), .A2(new_n462_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n481_), .A2(new_n483_), .A3(new_n494_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT12), .ZN(new_n521_));
  INV_X1    g320(.A(new_n506_), .ZN(new_n522_));
  AND3_X1   g321(.A1(new_n520_), .A2(new_n521_), .A3(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n521_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n519_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n518_), .A2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G120gat), .B(G148gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT5), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G176gat), .B(G204gat), .ZN(new_n529_));
  XOR2_X1   g328(.A(new_n528_), .B(new_n529_), .Z(new_n530_));
  NAND2_X1  g329(.A1(new_n526_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n530_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n518_), .A2(new_n525_), .A3(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n531_), .A2(KEYINPUT67), .A3(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(KEYINPUT67), .B1(new_n531_), .B2(new_n533_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n461_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n536_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n538_), .A2(new_n534_), .A3(KEYINPUT13), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n537_), .A2(new_n539_), .ZN(new_n540_));
  XOR2_X1   g339(.A(new_n540_), .B(KEYINPUT68), .Z(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n520_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT35), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G232gat), .A2(G233gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT34), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  AOI22_X1  g346(.A1(new_n516_), .A2(new_n437_), .B1(new_n544_), .B2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n543_), .A2(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n547_), .A2(new_n544_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n548_), .B(new_n543_), .C1(new_n544_), .C2(new_n547_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G190gat), .B(G218gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G134gat), .B(G162gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n555_), .A2(KEYINPUT36), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n551_), .A2(new_n552_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  XOR2_X1   g357(.A(new_n555_), .B(KEYINPUT36), .Z(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n560_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n561_));
  OAI21_X1  g360(.A(KEYINPUT37), .B1(new_n558_), .B2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT70), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n561_), .A2(KEYINPUT71), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT37), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n561_), .A2(KEYINPUT71), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n565_), .A2(new_n566_), .A3(new_n557_), .A4(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n562_), .A2(new_n563_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n564_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(G127gat), .B(G155gat), .Z(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT16), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G183gat), .B(G211gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT17), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n574_), .B(KEYINPUT17), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G231gat), .A2(G233gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n506_), .B(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(new_n425_), .ZN(new_n580_));
  MUX2_X1   g379(.A(new_n576_), .B(new_n577_), .S(new_n580_), .Z(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n570_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n411_), .A2(new_n460_), .A3(new_n542_), .A4(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n397_), .ZN(new_n586_));
  NOR3_X1   g385(.A1(new_n585_), .A2(new_n586_), .A3(new_n418_), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n587_), .A2(KEYINPUT38), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n565_), .A2(new_n557_), .A3(new_n567_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT97), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n591_), .B1(new_n406_), .B2(new_n410_), .ZN(new_n592_));
  NOR3_X1   g391(.A1(new_n540_), .A2(new_n581_), .A3(new_n459_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  OAI21_X1  g393(.A(G1gat), .B1(new_n594_), .B2(new_n586_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n587_), .A2(KEYINPUT38), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n588_), .A2(new_n595_), .A3(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT98), .ZN(G1324gat));
  OAI21_X1  g397(.A(G8gat), .B1(new_n594_), .B2(new_n409_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(KEYINPUT99), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(KEYINPUT39), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n599_), .A2(KEYINPUT99), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT40), .ZN(new_n604_));
  OR2_X1    g403(.A1(new_n409_), .A2(G8gat), .ZN(new_n605_));
  OAI22_X1  g404(.A1(new_n600_), .A2(KEYINPUT39), .B1(new_n585_), .B2(new_n605_), .ZN(new_n606_));
  OR3_X1    g405(.A1(new_n603_), .A2(new_n604_), .A3(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n604_), .B1(new_n603_), .B2(new_n606_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(G1325gat));
  OAI21_X1  g408(.A(G15gat), .B1(new_n594_), .B2(new_n259_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT41), .ZN(new_n611_));
  NOR3_X1   g410(.A1(new_n585_), .A2(G15gat), .A3(new_n259_), .ZN(new_n612_));
  OR2_X1    g411(.A1(new_n611_), .A2(new_n612_), .ZN(G1326gat));
  OAI21_X1  g412(.A(G22gat), .B1(new_n594_), .B2(new_n408_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT42), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n408_), .A2(G22gat), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n615_), .B1(new_n585_), .B2(new_n616_), .ZN(G1327gat));
  NOR2_X1   g416(.A1(new_n540_), .A2(new_n459_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n589_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(new_n581_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT101), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n411_), .A2(new_n618_), .A3(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(KEYINPUT102), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT102), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n411_), .A2(new_n618_), .A3(new_n624_), .A4(new_n621_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(G29gat), .B1(new_n627_), .B2(new_n397_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n618_), .A2(new_n581_), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n629_), .B(KEYINPUT100), .Z(new_n630_));
  INV_X1    g429(.A(KEYINPUT43), .ZN(new_n631_));
  INV_X1    g430(.A(new_n570_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n631_), .B1(new_n411_), .B2(new_n632_), .ZN(new_n633_));
  AOI211_X1 g432(.A(KEYINPUT43), .B(new_n570_), .C1(new_n406_), .C2(new_n410_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n630_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT44), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  OAI211_X1 g436(.A(new_n630_), .B(KEYINPUT44), .C1(new_n633_), .C2(new_n634_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n397_), .A2(G29gat), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n628_), .B1(new_n639_), .B2(new_n640_), .ZN(G1328gat));
  NAND3_X1  g440(.A1(new_n637_), .A2(new_n319_), .A3(new_n638_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(G36gat), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT103), .ZN(new_n644_));
  OAI21_X1  g443(.A(KEYINPUT104), .B1(new_n644_), .B2(KEYINPUT46), .ZN(new_n645_));
  NOR2_X1   g444(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n409_), .A2(G36gat), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n623_), .A2(new_n625_), .A3(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(KEYINPUT45), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT45), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n623_), .A2(new_n650_), .A3(new_n625_), .A4(new_n647_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n646_), .B1(new_n649_), .B2(new_n651_), .ZN(new_n652_));
  AND3_X1   g451(.A1(new_n643_), .A2(new_n645_), .A3(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n645_), .B1(new_n643_), .B2(new_n652_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1329gat));
  INV_X1    g454(.A(new_n259_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n637_), .A2(G43gat), .A3(new_n656_), .A4(new_n638_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n626_), .A2(new_n259_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n657_), .B1(G43gat), .B2(new_n658_), .ZN(new_n659_));
  XOR2_X1   g458(.A(KEYINPUT105), .B(KEYINPUT47), .Z(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(G1330gat));
  OR3_X1    g460(.A1(new_n626_), .A2(G50gat), .A3(new_n408_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT106), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n663_), .B1(new_n639_), .B2(new_n360_), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n637_), .A2(new_n663_), .A3(new_n360_), .A4(new_n638_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(G50gat), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n662_), .B1(new_n664_), .B2(new_n666_), .ZN(G1331gat));
  NOR3_X1   g466(.A1(new_n457_), .A2(new_n581_), .A3(new_n458_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n592_), .A2(new_n541_), .A3(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(G57gat), .B1(new_n669_), .B2(new_n586_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n460_), .B1(new_n406_), .B2(new_n410_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n671_), .A2(new_n540_), .A3(new_n584_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n397_), .A2(new_n501_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n670_), .B1(new_n672_), .B2(new_n673_), .ZN(G1332gat));
  OAI21_X1  g473(.A(G64gat), .B1(new_n669_), .B2(new_n409_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT48), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n319_), .A2(new_n499_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n676_), .B1(new_n672_), .B2(new_n677_), .ZN(G1333gat));
  OAI21_X1  g477(.A(G71gat), .B1(new_n669_), .B2(new_n259_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT49), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n259_), .A2(G71gat), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n680_), .B1(new_n672_), .B2(new_n681_), .ZN(G1334gat));
  OAI21_X1  g481(.A(G78gat), .B1(new_n669_), .B2(new_n408_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT50), .ZN(new_n684_));
  OR2_X1    g483(.A1(new_n408_), .A2(G78gat), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n684_), .B1(new_n672_), .B2(new_n685_), .ZN(G1335gat));
  AND2_X1   g485(.A1(new_n541_), .A2(new_n621_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n671_), .A2(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n464_), .B1(new_n688_), .B2(new_n586_), .ZN(new_n689_));
  OR2_X1    g488(.A1(new_n689_), .A2(KEYINPUT107), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(KEYINPUT107), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n633_), .A2(new_n634_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n540_), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n693_), .A2(new_n582_), .A3(new_n460_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n692_), .A2(new_n695_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n586_), .A2(new_n464_), .ZN(new_n697_));
  AOI22_X1  g496(.A1(new_n690_), .A2(new_n691_), .B1(new_n696_), .B2(new_n697_), .ZN(G1336gat));
  INV_X1    g497(.A(new_n688_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n699_), .A2(new_n465_), .A3(new_n319_), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n692_), .A2(new_n409_), .A3(new_n695_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n700_), .B1(new_n701_), .B2(new_n465_), .ZN(G1337gat));
  AND3_X1   g501(.A1(new_n656_), .A2(new_n490_), .A3(new_n492_), .ZN(new_n703_));
  AOI21_X1  g502(.A(KEYINPUT109), .B1(new_n699_), .B2(new_n703_), .ZN(new_n704_));
  OAI211_X1 g503(.A(new_n656_), .B(new_n694_), .C1(new_n633_), .C2(new_n634_), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n705_), .A2(KEYINPUT108), .A3(G99gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(KEYINPUT108), .B1(new_n705_), .B2(G99gat), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n704_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g508(.A1(new_n699_), .A2(new_n491_), .A3(new_n360_), .ZN(new_n710_));
  OAI211_X1 g509(.A(new_n360_), .B(new_n694_), .C1(new_n633_), .C2(new_n634_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT52), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n711_), .A2(new_n712_), .A3(G106gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n711_), .B2(G106gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n710_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g515(.A(KEYINPUT59), .ZN(new_n717_));
  NOR4_X1   g516(.A1(new_n319_), .A2(new_n259_), .A3(new_n586_), .A4(new_n360_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT58), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n507_), .A2(new_n462_), .ZN(new_n720_));
  OAI21_X1  g519(.A(KEYINPUT12), .B1(new_n516_), .B2(new_n506_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n520_), .A2(new_n521_), .A3(new_n522_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n720_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(KEYINPUT112), .B1(new_n723_), .B2(KEYINPUT55), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n523_), .A2(new_n524_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n463_), .B1(new_n725_), .B2(new_n514_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT112), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT55), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n525_), .A2(new_n727_), .A3(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n724_), .A2(new_n726_), .A3(new_n729_), .ZN(new_n730_));
  OAI211_X1 g529(.A(KEYINPUT55), .B(new_n519_), .C1(new_n523_), .C2(new_n524_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT113), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n721_), .A2(new_n722_), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n734_), .A2(KEYINPUT113), .A3(KEYINPUT55), .A4(new_n519_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n733_), .A2(new_n735_), .ZN(new_n736_));
  OAI211_X1 g535(.A(KEYINPUT56), .B(new_n530_), .C1(new_n730_), .C2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT116), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n733_), .A2(new_n735_), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n740_), .A2(new_n729_), .A3(new_n726_), .A4(new_n724_), .ZN(new_n741_));
  AOI21_X1  g540(.A(KEYINPUT56), .B1(new_n741_), .B2(new_n530_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n739_), .A2(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n530_), .B1(new_n730_), .B2(new_n736_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT56), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n744_), .A2(KEYINPUT116), .A3(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n412_), .B1(new_n436_), .B2(new_n439_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n747_), .B1(new_n443_), .B2(new_n447_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n455_), .B1(new_n451_), .B2(new_n412_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT115), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n748_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  AOI211_X1 g550(.A(KEYINPUT115), .B(new_n455_), .C1(new_n451_), .C2(new_n412_), .ZN(new_n752_));
  OAI211_X1 g551(.A(new_n456_), .B(new_n533_), .C1(new_n751_), .C2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n746_), .A2(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n719_), .B1(new_n743_), .B2(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n753_), .B1(new_n742_), .B2(KEYINPUT116), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n757_), .B(KEYINPUT58), .C1(new_n742_), .C2(new_n739_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n756_), .A2(new_n758_), .A3(new_n632_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n533_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n459_), .A2(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n737_), .B1(new_n742_), .B2(KEYINPUT114), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n744_), .A2(KEYINPUT114), .A3(new_n745_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n761_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  OAI221_X1 g563(.A(new_n456_), .B1(new_n752_), .B2(new_n751_), .C1(new_n535_), .C2(new_n536_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n619_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n759_), .B1(new_n766_), .B2(KEYINPUT57), .ZN(new_n767_));
  OR2_X1    g566(.A1(new_n767_), .A2(KEYINPUT118), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT57), .ZN(new_n769_));
  AOI211_X1 g568(.A(new_n769_), .B(new_n619_), .C1(new_n764_), .C2(new_n765_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n770_), .B1(new_n767_), .B2(KEYINPUT118), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n582_), .B1(new_n768_), .B2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n668_), .ZN(new_n773_));
  OAI21_X1  g572(.A(KEYINPUT110), .B1(new_n540_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT110), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n537_), .A2(new_n539_), .A3(new_n775_), .A4(new_n668_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n774_), .A2(new_n570_), .A3(new_n776_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(KEYINPUT111), .A2(KEYINPUT54), .ZN(new_n778_));
  NAND2_X1  g577(.A1(KEYINPUT111), .A2(KEYINPUT54), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n777_), .B1(new_n778_), .B2(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n781_), .B1(new_n777_), .B2(new_n780_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n717_), .B(new_n718_), .C1(new_n772_), .C2(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n460_), .A2(KEYINPUT119), .A3(G113gat), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n785_), .B1(KEYINPUT119), .B2(G113gat), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n581_), .B1(new_n767_), .B2(new_n770_), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n787_), .A2(KEYINPUT117), .A3(new_n782_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT117), .B1(new_n787_), .B2(new_n782_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n718_), .ZN(new_n790_));
  NOR3_X1   g589(.A1(new_n788_), .A2(new_n789_), .A3(new_n790_), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n784_), .B(new_n786_), .C1(new_n791_), .C2(new_n717_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n789_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n787_), .A2(new_n782_), .A3(KEYINPUT117), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n793_), .A2(new_n460_), .A3(new_n794_), .A4(new_n718_), .ZN(new_n795_));
  INV_X1    g594(.A(G113gat), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n792_), .A2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT120), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n792_), .A2(KEYINPUT120), .A3(new_n797_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(G1340gat));
  OAI21_X1  g601(.A(new_n784_), .B1(new_n791_), .B2(new_n717_), .ZN(new_n803_));
  OAI21_X1  g602(.A(G120gat), .B1(new_n803_), .B2(new_n542_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n693_), .A2(KEYINPUT60), .ZN(new_n805_));
  MUX2_X1   g604(.A(new_n805_), .B(KEYINPUT60), .S(G120gat), .Z(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT121), .B1(new_n791_), .B2(new_n806_), .ZN(new_n807_));
  AND3_X1   g606(.A1(new_n791_), .A2(KEYINPUT121), .A3(new_n806_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n804_), .B1(new_n807_), .B2(new_n808_), .ZN(G1341gat));
  INV_X1    g608(.A(G127gat), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n791_), .A2(new_n810_), .A3(new_n582_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n582_), .B(new_n784_), .C1(new_n791_), .C2(new_n717_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n811_), .B1(new_n813_), .B2(new_n810_), .ZN(G1342gat));
  INV_X1    g613(.A(G134gat), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n791_), .A2(new_n815_), .A3(new_n591_), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n632_), .B(new_n784_), .C1(new_n791_), .C2(new_n717_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n816_), .B1(new_n818_), .B2(new_n815_), .ZN(G1343gat));
  NOR2_X1   g618(.A1(new_n788_), .A2(new_n789_), .ZN(new_n820_));
  NOR4_X1   g619(.A1(new_n656_), .A2(new_n319_), .A3(new_n586_), .A4(new_n408_), .ZN(new_n821_));
  AND2_X1   g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n460_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n823_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g623(.A1(new_n820_), .A2(new_n821_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n825_), .A2(new_n542_), .ZN(new_n826_));
  XOR2_X1   g625(.A(KEYINPUT122), .B(G148gat), .Z(new_n827_));
  XNOR2_X1  g626(.A(new_n826_), .B(new_n827_), .ZN(G1345gat));
  NAND2_X1  g627(.A1(new_n822_), .A2(new_n582_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(KEYINPUT61), .B(G155gat), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n829_), .B(new_n830_), .ZN(G1346gat));
  NAND3_X1  g630(.A1(new_n822_), .A2(new_n321_), .A3(new_n591_), .ZN(new_n832_));
  OAI21_X1  g631(.A(G162gat), .B1(new_n825_), .B2(new_n570_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(G1347gat));
  NAND2_X1  g633(.A1(new_n407_), .A2(new_n319_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n835_), .A2(new_n360_), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n460_), .B(new_n836_), .C1(new_n772_), .C2(new_n783_), .ZN(new_n837_));
  AOI21_X1  g636(.A(KEYINPUT123), .B1(new_n837_), .B2(G169gat), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT62), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n837_), .A2(KEYINPUT123), .A3(G169gat), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n837_), .ZN(new_n843_));
  AOI22_X1  g642(.A1(new_n838_), .A2(new_n839_), .B1(new_n240_), .B2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n842_), .A2(new_n844_), .ZN(G1348gat));
  OAI21_X1  g644(.A(new_n836_), .B1(new_n772_), .B2(new_n783_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(G176gat), .B1(new_n847_), .B2(new_n540_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n788_), .A2(new_n789_), .A3(new_n360_), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n542_), .A2(new_n835_), .A3(new_n241_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n848_), .B1(new_n849_), .B2(new_n850_), .ZN(G1349gat));
  NOR3_X1   g650(.A1(new_n846_), .A2(new_n231_), .A3(new_n581_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n849_), .A2(new_n319_), .A3(new_n407_), .A4(new_n582_), .ZN(new_n853_));
  INV_X1    g652(.A(G183gat), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n852_), .B1(new_n853_), .B2(new_n854_), .ZN(G1350gat));
  OAI21_X1  g654(.A(G190gat), .B1(new_n846_), .B2(new_n570_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n591_), .A2(new_n232_), .ZN(new_n857_));
  XOR2_X1   g656(.A(new_n857_), .B(KEYINPUT124), .Z(new_n858_));
  OAI21_X1  g657(.A(new_n856_), .B1(new_n846_), .B2(new_n858_), .ZN(G1351gat));
  NOR3_X1   g658(.A1(new_n409_), .A2(new_n656_), .A3(new_n386_), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n793_), .A2(new_n794_), .A3(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n861_), .A2(G197gat), .A3(new_n460_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT125), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(G197gat), .ZN(new_n865_));
  INV_X1    g664(.A(new_n861_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(new_n866_), .B2(new_n459_), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n861_), .A2(KEYINPUT125), .A3(G197gat), .A4(new_n460_), .ZN(new_n868_));
  AND3_X1   g667(.A1(new_n864_), .A2(new_n867_), .A3(new_n868_), .ZN(G1352gat));
  NAND2_X1  g668(.A1(new_n861_), .A2(new_n541_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g670(.A(KEYINPUT63), .B(G211gat), .C1(new_n861_), .C2(new_n582_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n866_), .A2(new_n581_), .ZN(new_n873_));
  XOR2_X1   g672(.A(KEYINPUT63), .B(G211gat), .Z(new_n874_));
  AOI21_X1  g673(.A(new_n872_), .B1(new_n873_), .B2(new_n874_), .ZN(G1354gat));
  XNOR2_X1  g674(.A(KEYINPUT127), .B(G218gat), .ZN(new_n876_));
  NOR3_X1   g675(.A1(new_n866_), .A2(new_n570_), .A3(new_n876_), .ZN(new_n877_));
  NAND4_X1  g676(.A1(new_n793_), .A2(new_n591_), .A3(new_n794_), .A4(new_n860_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT126), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n878_), .B(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n877_), .B1(new_n880_), .B2(new_n876_), .ZN(G1355gat));
endmodule


