//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 1 0 0 1 0 1 1 0 0 0 1 0 1 1 0 1 0 1 0 0 1 1 0 1 0 0 0 1 0 1 1 0 0 0 1 0 0 1 1 0 0 1 1 1 1 1 1 1 1 1 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n786_, new_n787_, new_n788_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n885_, new_n887_, new_n888_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n917_,
    new_n918_, new_n919_, new_n921_, new_n922_, new_n923_, new_n924_,
    new_n926_, new_n927_, new_n928_, new_n930_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_;
  XOR2_X1   g000(.A(KEYINPUT10), .B(G99gat), .Z(new_n202_));
  INV_X1    g001(.A(G106gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G85gat), .ZN(new_n205_));
  INV_X1    g004(.A(G92gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G85gat), .A2(G92gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n207_), .A2(KEYINPUT9), .A3(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(G99gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT6), .B1(new_n210_), .B2(new_n203_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT6), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(G99gat), .A3(G106gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  OR2_X1    g013(.A1(new_n208_), .A2(KEYINPUT9), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n204_), .A2(new_n209_), .A3(new_n214_), .A4(new_n215_), .ZN(new_n216_));
  OR3_X1    g015(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT64), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT64), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n220_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n214_), .A2(new_n217_), .A3(new_n219_), .A4(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT8), .ZN(new_n223_));
  AND3_X1   g022(.A1(new_n207_), .A2(KEYINPUT65), .A3(new_n208_), .ZN(new_n224_));
  AND3_X1   g023(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n223_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n216_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G29gat), .B(G36gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G43gat), .B(G50gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  XOR2_X1   g029(.A(KEYINPUT68), .B(KEYINPUT15), .Z(new_n231_));
  XNOR2_X1  g030(.A(new_n230_), .B(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n227_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT69), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G232gat), .A2(G233gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT34), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT35), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  OAI211_X1 g038(.A(new_n230_), .B(new_n216_), .C1(new_n225_), .C2(new_n226_), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n233_), .A2(new_n234_), .A3(new_n239_), .A4(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n237_), .A2(new_n238_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n233_), .A2(new_n240_), .A3(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n239_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n245_), .B1(new_n233_), .B2(KEYINPUT69), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n241_), .B1(new_n244_), .B2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G190gat), .B(G218gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G134gat), .B(G162gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  XOR2_X1   g050(.A(KEYINPUT70), .B(KEYINPUT36), .Z(new_n252_));
  NAND3_X1  g051(.A1(new_n247_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n253_));
  XOR2_X1   g052(.A(new_n250_), .B(KEYINPUT36), .Z(new_n254_));
  OAI211_X1 g053(.A(new_n241_), .B(new_n254_), .C1(new_n244_), .C2(new_n246_), .ZN(new_n255_));
  XOR2_X1   g054(.A(KEYINPUT73), .B(KEYINPUT37), .Z(new_n256_));
  NAND3_X1  g055(.A1(new_n253_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT74), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n253_), .A2(KEYINPUT74), .A3(new_n255_), .A4(new_n256_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n255_), .A2(KEYINPUT71), .ZN(new_n262_));
  INV_X1    g061(.A(new_n246_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(new_n243_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT71), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n264_), .A2(new_n265_), .A3(new_n241_), .A4(new_n254_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n253_), .A2(new_n262_), .A3(new_n266_), .ZN(new_n267_));
  AND3_X1   g066(.A1(new_n267_), .A2(KEYINPUT72), .A3(KEYINPUT37), .ZN(new_n268_));
  AOI21_X1  g067(.A(KEYINPUT72), .B1(new_n267_), .B2(KEYINPUT37), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n261_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G57gat), .B(G64gat), .ZN(new_n272_));
  OR2_X1    g071(.A1(new_n272_), .A2(KEYINPUT11), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(KEYINPUT11), .ZN(new_n274_));
  XOR2_X1   g073(.A(G71gat), .B(G78gat), .Z(new_n275_));
  NAND3_X1  g074(.A1(new_n273_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n274_), .A2(new_n275_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n227_), .A2(new_n279_), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n216_), .B(new_n278_), .C1(new_n225_), .C2(new_n226_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT12), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n279_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n282_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n216_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n222_), .A2(new_n224_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT8), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n286_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n283_), .B1(new_n290_), .B2(new_n278_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT66), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G230gat), .A2(G233gat), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n280_), .A2(KEYINPUT66), .A3(new_n283_), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n285_), .A2(new_n293_), .A3(new_n294_), .A4(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n294_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n282_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(G120gat), .B(G148gat), .Z(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G176gat), .B(G204gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n299_), .B(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT13), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n299_), .B(new_n304_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT13), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n307_), .A2(new_n310_), .ZN(new_n311_));
  XOR2_X1   g110(.A(G127gat), .B(G155gat), .Z(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G183gat), .B(G211gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT17), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n317_), .A2(KEYINPUT77), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  OR2_X1    g118(.A1(new_n316_), .A2(KEYINPUT17), .ZN(new_n320_));
  XOR2_X1   g119(.A(G1gat), .B(G8gat), .Z(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G1gat), .A2(G8gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT14), .ZN(new_n324_));
  INV_X1    g123(.A(G15gat), .ZN(new_n325_));
  INV_X1    g124(.A(G22gat), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(G15gat), .A2(G22gat), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n324_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n329_), .A2(KEYINPUT75), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT76), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n329_), .A2(KEYINPUT75), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n331_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n332_), .B1(new_n331_), .B2(new_n333_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n322_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n336_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n338_), .A2(new_n321_), .A3(new_n334_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n340_), .A2(G231gat), .A3(G233gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G231gat), .A2(G233gat), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n337_), .A2(new_n339_), .A3(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n341_), .A2(new_n278_), .A3(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n278_), .B1(new_n341_), .B2(new_n343_), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n319_), .B(new_n320_), .C1(new_n345_), .C2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n341_), .A2(new_n343_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(new_n279_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n349_), .A2(new_n316_), .A3(new_n318_), .A4(new_n344_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n347_), .A2(new_n350_), .ZN(new_n351_));
  NOR3_X1   g150(.A1(new_n271_), .A2(new_n311_), .A3(new_n351_), .ZN(new_n352_));
  OR2_X1    g151(.A1(new_n352_), .A2(KEYINPUT79), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G127gat), .B(G134gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G113gat), .B(G120gat), .ZN(new_n355_));
  AND2_X1   g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n354_), .A2(new_n355_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(G155gat), .A2(G162gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G155gat), .A2(G162gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT85), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT85), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n363_), .A2(G155gat), .A3(G162gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n360_), .B1(new_n365_), .B2(KEYINPUT1), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT1), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n362_), .A2(new_n364_), .A3(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT86), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT86), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n362_), .A2(new_n364_), .A3(new_n370_), .A4(new_n367_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n366_), .A2(new_n369_), .A3(new_n371_), .ZN(new_n372_));
  XOR2_X1   g171(.A(G141gat), .B(G148gat), .Z(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT3), .ZN(new_n375_));
  INV_X1    g174(.A(G141gat), .ZN(new_n376_));
  INV_X1    g175(.A(G148gat), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n375_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G141gat), .A2(G148gat), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT2), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n382_));
  OAI21_X1  g181(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n378_), .A2(new_n381_), .A3(new_n382_), .A4(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n360_), .ZN(new_n385_));
  AND3_X1   g184(.A1(new_n384_), .A2(new_n365_), .A3(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n359_), .B1(new_n374_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n386_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(new_n359_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G225gat), .A2(G233gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(KEYINPUT96), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n389_), .A2(new_n391_), .A3(new_n394_), .ZN(new_n395_));
  AOI211_X1 g194(.A(new_n386_), .B(new_n358_), .C1(new_n372_), .C2(new_n373_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT4), .ZN(new_n397_));
  NOR3_X1   g196(.A1(new_n396_), .A2(new_n388_), .A3(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n374_), .A2(new_n387_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n399_), .A2(new_n397_), .A3(new_n358_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(new_n393_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n395_), .B1(new_n398_), .B2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G1gat), .B(G29gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(G85gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(KEYINPUT0), .B(G57gat), .ZN(new_n405_));
  XOR2_X1   g204(.A(new_n404_), .B(new_n405_), .Z(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n402_), .A2(new_n407_), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n395_), .B(new_n406_), .C1(new_n398_), .C2(new_n401_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n408_), .A2(KEYINPUT97), .A3(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT97), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n402_), .A2(new_n411_), .A3(new_n407_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT21), .ZN(new_n413_));
  AND2_X1   g212(.A1(G197gat), .A2(G204gat), .ZN(new_n414_));
  NOR2_X1   g213(.A1(G197gat), .A2(G204gat), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n413_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(G197gat), .ZN(new_n417_));
  INV_X1    g216(.A(G204gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G197gat), .A2(G204gat), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n419_), .A2(KEYINPUT21), .A3(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(G218gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(G211gat), .ZN(new_n423_));
  INV_X1    g222(.A(G211gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(G218gat), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n416_), .A2(new_n421_), .A3(new_n423_), .A4(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT87), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n424_), .A2(G218gat), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n422_), .A2(G211gat), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n427_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n423_), .A2(new_n425_), .A3(KEYINPUT87), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n430_), .A2(KEYINPUT21), .A3(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT88), .B1(new_n414_), .B2(new_n415_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT88), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n419_), .A2(new_n434_), .A3(new_n420_), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n426_), .B1(new_n432_), .B2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G183gat), .A2(G190gat), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT23), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n441_));
  INV_X1    g240(.A(G183gat), .ZN(new_n442_));
  INV_X1    g241(.A(G190gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n440_), .A2(new_n441_), .A3(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G169gat), .A2(G176gat), .ZN(new_n446_));
  OR2_X1    g245(.A1(KEYINPUT82), .A2(G176gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(KEYINPUT82), .A2(G176gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(G169gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT22), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT22), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(G169gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n451_), .A2(new_n453_), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n445_), .B(new_n446_), .C1(new_n449_), .C2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n438_), .A2(KEYINPUT23), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n439_), .A2(G183gat), .A3(G190gat), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT24), .ZN(new_n458_));
  NOR2_X1   g257(.A1(G169gat), .A2(G176gat), .ZN(new_n459_));
  AOI22_X1  g258(.A1(new_n456_), .A2(new_n457_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n459_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n461_), .A2(KEYINPUT24), .A3(new_n446_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT25), .B1(new_n442_), .B2(KEYINPUT81), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT81), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT25), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n465_), .A2(new_n466_), .A3(G183gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n443_), .A2(KEYINPUT26), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT26), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(G190gat), .ZN(new_n470_));
  AND4_X1   g269(.A1(new_n464_), .A2(new_n467_), .A3(new_n468_), .A4(new_n470_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n455_), .B1(new_n463_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n437_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT94), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n437_), .A2(new_n472_), .A3(KEYINPUT94), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n469_), .A2(G190gat), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n443_), .A2(KEYINPUT26), .ZN(new_n479_));
  OAI21_X1  g278(.A(KEYINPUT91), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(KEYINPUT25), .B(G183gat), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT91), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n468_), .A2(new_n470_), .A3(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n480_), .A2(new_n481_), .A3(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n446_), .A2(KEYINPUT24), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT92), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n446_), .A2(KEYINPUT92), .A3(KEYINPUT24), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n487_), .A2(new_n461_), .A3(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n484_), .A2(new_n460_), .A3(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n433_), .A2(new_n435_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n491_), .A2(KEYINPUT21), .A3(new_n431_), .A4(new_n430_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n446_), .B(KEYINPUT93), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n493_), .B(new_n445_), .C1(new_n449_), .C2(new_n454_), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n490_), .A2(new_n426_), .A3(new_n492_), .A4(new_n494_), .ZN(new_n495_));
  AND2_X1   g294(.A1(new_n495_), .A2(KEYINPUT20), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT95), .ZN(new_n497_));
  XNOR2_X1  g296(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G226gat), .A2(G233gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n477_), .A2(new_n496_), .A3(new_n497_), .A4(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n437_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n503_), .B1(new_n490_), .B2(new_n494_), .ZN(new_n504_));
  OAI21_X1  g303(.A(KEYINPUT20), .B1(new_n437_), .B2(new_n472_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n500_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n502_), .A2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G8gat), .B(G36gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT18), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G64gat), .B(G92gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(KEYINPUT32), .ZN(new_n513_));
  AND3_X1   g312(.A1(new_n437_), .A2(new_n472_), .A3(KEYINPUT94), .ZN(new_n514_));
  AOI21_X1  g313(.A(KEYINPUT94), .B1(new_n437_), .B2(new_n472_), .ZN(new_n515_));
  OAI211_X1 g314(.A(KEYINPUT20), .B(new_n495_), .C1(new_n514_), .C2(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(KEYINPUT95), .B1(new_n516_), .B2(new_n500_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n507_), .A2(new_n513_), .A3(new_n517_), .ZN(new_n518_));
  OR3_X1    g317(.A1(new_n504_), .A2(new_n500_), .A3(new_n505_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n495_), .A2(KEYINPUT20), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n520_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n519_), .B1(new_n501_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n513_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n410_), .A2(new_n412_), .A3(new_n518_), .A4(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT33), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n389_), .A2(new_n391_), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n394_), .B(new_n400_), .C1(new_n527_), .C2(new_n397_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n396_), .A2(new_n388_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n406_), .B1(new_n529_), .B2(new_n393_), .ZN(new_n530_));
  AOI22_X1  g329(.A1(new_n409_), .A2(new_n526_), .B1(new_n528_), .B2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n502_), .A2(new_n506_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n497_), .B1(new_n521_), .B2(new_n501_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n511_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n398_), .A2(new_n401_), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n535_), .A2(KEYINPUT33), .A3(new_n395_), .A4(new_n406_), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n517_), .A2(new_n512_), .A3(new_n506_), .A4(new_n502_), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n531_), .A2(new_n534_), .A3(new_n536_), .A4(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n525_), .A2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G22gat), .B(G50gat), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT28), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT29), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n390_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n542_), .B1(new_n390_), .B2(new_n543_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n541_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n546_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n548_), .A2(new_n544_), .A3(new_n540_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT89), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n503_), .B1(new_n399_), .B2(KEYINPUT29), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G228gat), .A2(G233gat), .ZN(new_n554_));
  INV_X1    g353(.A(G78gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(G106gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n553_), .B(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n547_), .A2(new_n549_), .A3(KEYINPUT89), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n552_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n550_), .A2(new_n558_), .A3(new_n551_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n539_), .A2(new_n563_), .ZN(new_n564_));
  AND3_X1   g363(.A1(new_n550_), .A2(new_n558_), .A3(new_n551_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n558_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n565_), .B1(new_n560_), .B2(new_n566_), .ZN(new_n567_));
  XOR2_X1   g366(.A(KEYINPUT98), .B(KEYINPUT27), .Z(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n512_), .B1(new_n507_), .B2(new_n517_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n537_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n569_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n410_), .A2(new_n412_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT27), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n574_), .B1(new_n522_), .B2(new_n511_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(new_n537_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n567_), .A2(new_n572_), .A3(new_n573_), .A4(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n564_), .A2(new_n577_), .ZN(new_n578_));
  XOR2_X1   g377(.A(G71gat), .B(G99gat), .Z(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(G43gat), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n472_), .A2(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n472_), .A2(new_n580_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G227gat), .A2(G233gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(new_n325_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT30), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  OR3_X1    g385(.A1(new_n581_), .A2(new_n582_), .A3(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT84), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n586_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n590_));
  XOR2_X1   g389(.A(new_n358_), .B(new_n590_), .Z(new_n591_));
  NAND4_X1  g390(.A1(new_n587_), .A2(new_n588_), .A3(new_n589_), .A4(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n587_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n591_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n588_), .B1(new_n587_), .B2(new_n589_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n592_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n597_), .B1(new_n410_), .B2(new_n412_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n598_), .A2(new_n572_), .A3(new_n563_), .A4(new_n576_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(KEYINPUT99), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n534_), .A2(new_n537_), .ZN(new_n601_));
  AOI22_X1  g400(.A1(new_n601_), .A2(new_n569_), .B1(new_n537_), .B2(new_n575_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT99), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n602_), .A2(new_n603_), .A3(new_n563_), .A4(new_n598_), .ZN(new_n604_));
  AOI22_X1  g403(.A1(new_n578_), .A2(new_n597_), .B1(new_n600_), .B2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G113gat), .B(G141gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G169gat), .B(G197gat), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n606_), .B(new_n607_), .Z(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n337_), .A2(new_n339_), .A3(new_n230_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(G229gat), .A2(G233gat), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT80), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n613_), .B1(new_n340_), .B2(new_n232_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n340_), .A2(new_n613_), .A3(new_n232_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n612_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n230_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n340_), .A2(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n611_), .B1(new_n619_), .B2(new_n610_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n609_), .B1(new_n617_), .B2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n620_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n616_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n623_), .A2(new_n614_), .ZN(new_n624_));
  OAI211_X1 g423(.A(new_n622_), .B(new_n608_), .C1(new_n624_), .C2(new_n612_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n621_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n605_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n352_), .A2(KEYINPUT79), .ZN(new_n629_));
  AND3_X1   g428(.A1(new_n353_), .A2(new_n628_), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(G1gat), .ZN(new_n631_));
  INV_X1    g430(.A(new_n573_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n630_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT38), .ZN(new_n634_));
  NOR3_X1   g433(.A1(new_n311_), .A2(new_n627_), .A3(new_n351_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT100), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n253_), .A2(new_n255_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n605_), .A2(new_n638_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n636_), .A2(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n631_), .B1(new_n640_), .B2(new_n632_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT101), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n634_), .A2(new_n642_), .ZN(G1324gat));
  INV_X1    g442(.A(G8gat), .ZN(new_n644_));
  INV_X1    g443(.A(new_n602_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n630_), .A2(new_n644_), .A3(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n640_), .A2(new_n645_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(KEYINPUT102), .A2(KEYINPUT39), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n644_), .B1(KEYINPUT102), .B2(KEYINPUT39), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n648_), .A2(new_n649_), .A3(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n649_), .B1(new_n648_), .B2(new_n650_), .ZN(new_n653_));
  OAI211_X1 g452(.A(new_n646_), .B(new_n647_), .C1(new_n652_), .C2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n648_), .A2(new_n650_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n649_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(new_n651_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n647_), .B1(new_n659_), .B2(new_n646_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n655_), .A2(new_n660_), .ZN(G1325gat));
  INV_X1    g460(.A(new_n597_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n630_), .A2(new_n325_), .A3(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n640_), .A2(new_n662_), .ZN(new_n664_));
  AND3_X1   g463(.A1(new_n664_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n665_));
  AOI21_X1  g464(.A(KEYINPUT41), .B1(new_n664_), .B2(G15gat), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n663_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT104), .ZN(G1326gat));
  XNOR2_X1  g467(.A(new_n563_), .B(KEYINPUT105), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n326_), .B1(new_n640_), .B2(new_n669_), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT42), .Z(new_n671_));
  NAND3_X1  g470(.A1(new_n630_), .A2(new_n326_), .A3(new_n669_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1327gat));
  INV_X1    g472(.A(KEYINPUT44), .ZN(new_n674_));
  INV_X1    g473(.A(new_n351_), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n311_), .A2(new_n627_), .A3(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  OAI21_X1  g476(.A(KEYINPUT43), .B1(new_n605_), .B2(new_n270_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT43), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n600_), .A2(new_n604_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n662_), .B1(new_n564_), .B2(new_n577_), .ZN(new_n681_));
  OAI211_X1 g480(.A(new_n679_), .B(new_n271_), .C1(new_n680_), .C2(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n677_), .B1(new_n678_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT106), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n674_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  AOI211_X1 g484(.A(KEYINPUT106), .B(new_n677_), .C1(new_n678_), .C2(new_n682_), .ZN(new_n686_));
  OAI21_X1  g485(.A(KEYINPUT107), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n577_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n567_), .B1(new_n525_), .B2(new_n538_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n597_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n600_), .A2(new_n604_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n679_), .B1(new_n692_), .B2(new_n271_), .ZN(new_n693_));
  AOI211_X1 g492(.A(KEYINPUT43), .B(new_n270_), .C1(new_n690_), .C2(new_n691_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n676_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(KEYINPUT106), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT107), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n678_), .A2(new_n682_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n698_), .A2(new_n684_), .A3(new_n676_), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n696_), .A2(new_n697_), .A3(new_n674_), .A4(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n687_), .A2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n683_), .A2(KEYINPUT44), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  OAI21_X1  g502(.A(G29gat), .B1(new_n703_), .B2(new_n573_), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n311_), .A2(new_n637_), .A3(new_n675_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n628_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(G29gat), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n632_), .A2(new_n708_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT108), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n704_), .B1(new_n707_), .B2(new_n710_), .ZN(G1328gat));
  INV_X1    g510(.A(G36gat), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n706_), .A2(new_n712_), .A3(new_n645_), .ZN(new_n713_));
  XOR2_X1   g512(.A(KEYINPUT109), .B(KEYINPUT45), .Z(new_n714_));
  XNOR2_X1  g513(.A(new_n713_), .B(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n702_), .A2(new_n645_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n716_), .B1(new_n687_), .B2(new_n700_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n715_), .B1(new_n717_), .B2(new_n712_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT46), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  OAI211_X1 g519(.A(KEYINPUT46), .B(new_n715_), .C1(new_n717_), .C2(new_n712_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1329gat));
  XNOR2_X1  g521(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n662_), .A2(G43gat), .ZN(new_n725_));
  INV_X1    g524(.A(new_n702_), .ZN(new_n726_));
  AOI211_X1 g525(.A(new_n725_), .B(new_n726_), .C1(new_n687_), .C2(new_n700_), .ZN(new_n727_));
  AOI21_X1  g526(.A(G43gat), .B1(new_n706_), .B2(new_n662_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n724_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n728_), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n730_), .B(new_n723_), .C1(new_n703_), .C2(new_n725_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(G1330gat));
  INV_X1    g531(.A(G50gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n706_), .A2(new_n733_), .A3(new_n669_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n726_), .A2(new_n563_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n701_), .A2(KEYINPUT111), .A3(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(G50gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(KEYINPUT111), .B1(new_n701_), .B2(new_n735_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n734_), .B1(new_n737_), .B2(new_n738_), .ZN(G1331gat));
  INV_X1    g538(.A(new_n311_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n740_), .A2(new_n626_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n692_), .A2(new_n741_), .A3(new_n675_), .A4(new_n270_), .ZN(new_n742_));
  XOR2_X1   g541(.A(new_n742_), .B(KEYINPUT112), .Z(new_n743_));
  INV_X1    g542(.A(G57gat), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n743_), .A2(new_n744_), .A3(new_n632_), .ZN(new_n745_));
  NOR3_X1   g544(.A1(new_n740_), .A2(new_n626_), .A3(new_n351_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n639_), .A2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  OAI21_X1  g547(.A(G57gat), .B1(new_n748_), .B2(new_n573_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n745_), .A2(new_n749_), .ZN(G1332gat));
  INV_X1    g549(.A(G64gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(new_n747_), .B2(new_n645_), .ZN(new_n752_));
  XOR2_X1   g551(.A(new_n752_), .B(KEYINPUT48), .Z(new_n753_));
  NAND3_X1  g552(.A1(new_n743_), .A2(new_n751_), .A3(new_n645_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(G1333gat));
  INV_X1    g554(.A(G71gat), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n743_), .A2(new_n756_), .A3(new_n662_), .ZN(new_n757_));
  OAI21_X1  g556(.A(G71gat), .B1(new_n748_), .B2(new_n597_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n758_), .A2(KEYINPUT49), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n758_), .A2(KEYINPUT49), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n757_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT113), .ZN(G1334gat));
  AOI21_X1  g561(.A(new_n555_), .B1(new_n747_), .B2(new_n669_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT114), .ZN(new_n764_));
  OR2_X1    g563(.A1(new_n764_), .A2(KEYINPUT50), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(KEYINPUT50), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n743_), .A2(new_n555_), .A3(new_n669_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n765_), .A2(new_n766_), .A3(new_n767_), .ZN(G1335gat));
  NAND2_X1  g567(.A1(new_n741_), .A2(new_n351_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n693_), .A2(new_n694_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n770_), .B2(KEYINPUT115), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n771_), .B1(KEYINPUT115), .B2(new_n770_), .ZN(new_n772_));
  OAI21_X1  g571(.A(G85gat), .B1(new_n772_), .B2(new_n573_), .ZN(new_n773_));
  AND4_X1   g572(.A1(new_n638_), .A2(new_n692_), .A3(new_n741_), .A4(new_n351_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n774_), .A2(new_n205_), .A3(new_n632_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(G1336gat));
  NAND2_X1  g575(.A1(new_n645_), .A2(G92gat), .ZN(new_n777_));
  OR2_X1    g576(.A1(new_n772_), .A2(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(G92gat), .B1(new_n774_), .B2(new_n645_), .ZN(new_n779_));
  XOR2_X1   g578(.A(new_n779_), .B(KEYINPUT116), .Z(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT117), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n778_), .A2(new_n780_), .A3(KEYINPUT117), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(G1337gat));
  OAI21_X1  g584(.A(G99gat), .B1(new_n772_), .B2(new_n597_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n774_), .A2(new_n202_), .A3(new_n662_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g588(.A1(new_n774_), .A2(new_n203_), .A3(new_n567_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT118), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n769_), .A2(new_n563_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n203_), .B1(new_n698_), .B2(new_n792_), .ZN(new_n793_));
  OR2_X1    g592(.A1(new_n793_), .A2(KEYINPUT52), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(KEYINPUT52), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n791_), .A2(new_n794_), .A3(new_n795_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT53), .ZN(G1339gat));
  AND4_X1   g596(.A1(new_n621_), .A2(new_n347_), .A3(new_n625_), .A4(new_n350_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n798_), .A2(new_n310_), .A3(new_n307_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT119), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n798_), .A2(new_n310_), .A3(new_n307_), .A4(KEYINPUT119), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n270_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT54), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n299_), .A2(new_n304_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n806_), .B1(new_n621_), .B2(new_n625_), .ZN(new_n807_));
  AOI22_X1  g606(.A1(new_n282_), .A2(new_n284_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n294_), .B1(new_n808_), .B2(new_n295_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n296_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n808_), .A2(KEYINPUT55), .A3(new_n294_), .A4(new_n295_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT56), .B1(new_n813_), .B2(new_n304_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT56), .ZN(new_n815_));
  AOI211_X1 g614(.A(new_n815_), .B(new_n305_), .C1(new_n811_), .C2(new_n812_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n807_), .B1(new_n814_), .B2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n619_), .A2(new_n610_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n608_), .B1(new_n818_), .B2(new_n611_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n610_), .A2(G229gat), .A3(G233gat), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n819_), .B1(new_n624_), .B2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n625_), .A2(new_n821_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n306_), .A2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n638_), .B1(new_n817_), .B2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(KEYINPUT57), .B1(new_n825_), .B2(KEYINPUT120), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT120), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT57), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n285_), .A2(new_n295_), .A3(new_n293_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n810_), .B1(new_n829_), .B2(new_n297_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n296_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n812_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n304_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n815_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n813_), .A2(KEYINPUT56), .A3(new_n304_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n823_), .B1(new_n837_), .B2(new_n807_), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n827_), .B(new_n828_), .C1(new_n838_), .C2(new_n638_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n822_), .A2(new_n806_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(new_n814_), .B2(new_n816_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT58), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n270_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n843_), .B1(new_n842_), .B2(new_n841_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n826_), .A2(new_n839_), .A3(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n351_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n805_), .A2(new_n846_), .ZN(new_n847_));
  NOR4_X1   g646(.A1(new_n645_), .A2(new_n573_), .A3(new_n567_), .A4(new_n597_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(G113gat), .B1(new_n850_), .B2(new_n626_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT121), .ZN(new_n852_));
  AND3_X1   g651(.A1(new_n845_), .A2(new_n852_), .A3(new_n351_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n852_), .B1(new_n845_), .B2(new_n351_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n805_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT59), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n848_), .A2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n855_), .A2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n849_), .A2(KEYINPUT59), .ZN(new_n860_));
  AND2_X1   g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n626_), .A2(G113gat), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(KEYINPUT122), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n851_), .B1(new_n861_), .B2(new_n863_), .ZN(G1340gat));
  INV_X1    g663(.A(G120gat), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n865_), .B1(new_n740_), .B2(KEYINPUT60), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n850_), .B(new_n866_), .C1(KEYINPUT60), .C2(new_n865_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n859_), .A2(new_n860_), .A3(new_n311_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n867_), .B1(new_n869_), .B2(new_n865_), .ZN(G1341gat));
  NAND3_X1  g669(.A1(new_n859_), .A2(new_n860_), .A3(new_n675_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(G127gat), .ZN(new_n872_));
  OR3_X1    g671(.A1(new_n849_), .A2(G127gat), .A3(new_n351_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(G1342gat));
  XNOR2_X1  g673(.A(KEYINPUT124), .B(G134gat), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n859_), .A2(new_n860_), .A3(new_n271_), .A4(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(G134gat), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n877_), .B1(new_n849_), .B2(new_n637_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT123), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  OAI211_X1 g679(.A(KEYINPUT123), .B(new_n877_), .C1(new_n849_), .C2(new_n637_), .ZN(new_n881_));
  AND3_X1   g680(.A1(new_n876_), .A2(new_n880_), .A3(new_n881_), .ZN(G1343gat));
  NOR3_X1   g681(.A1(new_n563_), .A2(new_n573_), .A3(new_n662_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n847_), .A2(new_n602_), .A3(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(new_n627_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(new_n376_), .ZN(G1344gat));
  NOR2_X1   g685(.A1(new_n884_), .A2(new_n740_), .ZN(new_n887_));
  XOR2_X1   g686(.A(KEYINPUT125), .B(G148gat), .Z(new_n888_));
  XNOR2_X1  g687(.A(new_n887_), .B(new_n888_), .ZN(G1345gat));
  NOR2_X1   g688(.A1(new_n884_), .A2(new_n351_), .ZN(new_n890_));
  XOR2_X1   g689(.A(KEYINPUT61), .B(G155gat), .Z(new_n891_));
  XNOR2_X1  g690(.A(new_n890_), .B(new_n891_), .ZN(G1346gat));
  OAI21_X1  g691(.A(G162gat), .B1(new_n884_), .B2(new_n270_), .ZN(new_n893_));
  OR2_X1    g692(.A1(new_n637_), .A2(G162gat), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n884_), .B2(new_n894_), .ZN(G1347gat));
  NAND2_X1  g694(.A1(new_n645_), .A2(new_n598_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n896_), .A2(new_n669_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n855_), .A2(new_n626_), .A3(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(G169gat), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT62), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  OR2_X1    g700(.A1(new_n898_), .A2(new_n454_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n898_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n901_), .A2(new_n902_), .A3(new_n903_), .ZN(G1348gat));
  INV_X1    g703(.A(new_n805_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n854_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n845_), .A2(new_n852_), .A3(new_n351_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n905_), .B1(new_n906_), .B2(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n897_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(new_n311_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n449_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n567_), .B1(new_n805_), .B2(new_n846_), .ZN(new_n913_));
  INV_X1    g712(.A(G176gat), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n740_), .A2(new_n914_), .A3(new_n896_), .ZN(new_n915_));
  AOI22_X1  g714(.A1(new_n911_), .A2(new_n912_), .B1(new_n913_), .B2(new_n915_), .ZN(G1349gat));
  NOR2_X1   g715(.A1(new_n896_), .A2(new_n351_), .ZN(new_n917_));
  AOI21_X1  g716(.A(G183gat), .B1(new_n913_), .B2(new_n917_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n351_), .A2(new_n481_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n918_), .B1(new_n910_), .B2(new_n919_), .ZN(G1350gat));
  NAND3_X1  g719(.A1(new_n638_), .A2(new_n480_), .A3(new_n483_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(KEYINPUT126), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n910_), .A2(new_n922_), .ZN(new_n923_));
  NOR3_X1   g722(.A1(new_n908_), .A2(new_n270_), .A3(new_n909_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n923_), .B1(new_n443_), .B2(new_n924_), .ZN(G1351gat));
  NOR3_X1   g724(.A1(new_n632_), .A2(new_n563_), .A3(new_n662_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n847_), .A2(new_n645_), .A3(new_n926_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n927_), .A2(new_n627_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(new_n417_), .ZN(G1352gat));
  NOR2_X1   g728(.A1(new_n927_), .A2(new_n740_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(new_n418_), .ZN(G1353gat));
  NOR2_X1   g730(.A1(new_n927_), .A2(new_n351_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n933_));
  INV_X1    g732(.A(new_n933_), .ZN(new_n934_));
  OAI21_X1  g733(.A(KEYINPUT127), .B1(new_n932_), .B2(new_n934_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT127), .ZN(new_n936_));
  OAI211_X1 g735(.A(new_n936_), .B(new_n933_), .C1(new_n927_), .C2(new_n351_), .ZN(new_n937_));
  XOR2_X1   g736(.A(KEYINPUT63), .B(G211gat), .Z(new_n938_));
  AOI22_X1  g737(.A1(new_n935_), .A2(new_n937_), .B1(new_n932_), .B2(new_n938_), .ZN(G1354gat));
  OAI21_X1  g738(.A(G218gat), .B1(new_n927_), .B2(new_n270_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n638_), .A2(new_n422_), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n940_), .B1(new_n927_), .B2(new_n941_), .ZN(G1355gat));
endmodule


