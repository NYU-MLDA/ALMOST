//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 1 1 1 0 1 0 0 1 1 1 0 0 0 0 1 0 1 1 1 0 1 1 0 1 1 1 0 0 0 1 0 1 0 1 0 0 1 0 0 0 0 1 1 1 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n780_, new_n781_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n918_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n928_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n960_,
    new_n961_, new_n962_, new_n963_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n971_, new_n972_, new_n973_, new_n974_,
    new_n976_, new_n977_, new_n978_, new_n980_, new_n981_, new_n982_,
    new_n983_, new_n984_, new_n985_;
  XNOR2_X1  g000(.A(G120gat), .B(G148gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT5), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G176gat), .B(G204gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  NAND2_X1  g004(.A1(G230gat), .A2(G233gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT64), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT6), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G85gat), .A2(G92gat), .ZN(new_n210_));
  OR2_X1    g009(.A1(new_n210_), .A2(KEYINPUT9), .ZN(new_n211_));
  OR2_X1    g010(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n212_));
  INV_X1    g011(.A(G106gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n212_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(G85gat), .ZN(new_n216_));
  INV_X1    g015(.A(G92gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(KEYINPUT9), .A3(new_n210_), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n209_), .A2(new_n211_), .A3(new_n215_), .A4(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  AND2_X1   g020(.A1(new_n218_), .A2(new_n210_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT6), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n208_), .B(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT7), .ZN(new_n225_));
  INV_X1    g024(.A(G99gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(new_n226_), .A3(new_n213_), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n222_), .B1(new_n224_), .B2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT8), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n223_), .B1(G99gat), .B2(G106gat), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n208_), .A2(KEYINPUT6), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n228_), .B(new_n227_), .C1(new_n232_), .C2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT8), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n234_), .A2(new_n235_), .A3(new_n222_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n221_), .B1(new_n231_), .B2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G57gat), .B(G64gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G71gat), .B(G78gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n238_), .A2(new_n239_), .A3(KEYINPUT11), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n238_), .A2(KEYINPUT11), .ZN(new_n241_));
  INV_X1    g040(.A(new_n239_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n238_), .A2(KEYINPUT11), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n240_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n237_), .A2(KEYINPUT65), .A3(new_n245_), .ZN(new_n246_));
  AND3_X1   g045(.A1(new_n234_), .A2(new_n235_), .A3(new_n222_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n235_), .B1(new_n234_), .B2(new_n222_), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n245_), .B(new_n220_), .C1(new_n247_), .C2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT65), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT66), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n246_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n220_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n245_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  AND2_X1   g055(.A1(new_n253_), .A2(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n252_), .B1(new_n246_), .B2(new_n251_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n207_), .B1(new_n257_), .B2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(KEYINPUT67), .A2(KEYINPUT12), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n261_), .B1(new_n237_), .B2(new_n245_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n207_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n263_), .B1(new_n237_), .B2(new_n245_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT67), .B(KEYINPUT12), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n254_), .A2(new_n255_), .A3(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n262_), .A2(new_n264_), .A3(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n262_), .A2(new_n264_), .A3(new_n266_), .A4(KEYINPUT68), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n205_), .B1(new_n260_), .B2(new_n271_), .ZN(new_n272_));
  AND2_X1   g071(.A1(new_n269_), .A2(new_n270_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n253_), .A2(new_n256_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n263_), .B1(new_n274_), .B2(new_n258_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n205_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n273_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n272_), .A2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT13), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G231gat), .A2(G233gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n245_), .B(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G1gat), .B(G8gat), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT77), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(G15gat), .ZN(new_n285_));
  INV_X1    g084(.A(G22gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G15gat), .A2(G22gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G1gat), .A2(G8gat), .ZN(new_n289_));
  AOI22_X1  g088(.A1(new_n287_), .A2(new_n288_), .B1(KEYINPUT14), .B2(new_n289_), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n284_), .A2(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n284_), .A2(new_n290_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n281_), .B(new_n293_), .ZN(new_n294_));
  XOR2_X1   g093(.A(G127gat), .B(G155gat), .Z(new_n295_));
  XNOR2_X1  g094(.A(G183gat), .B(G211gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  XOR2_X1   g096(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT17), .ZN(new_n300_));
  OR2_X1    g099(.A1(new_n294_), .A2(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n294_), .A2(KEYINPUT17), .A3(new_n299_), .ZN(new_n302_));
  AND2_X1   g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G190gat), .B(G218gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT70), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G134gat), .B(G162gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n305_), .A2(new_n306_), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT36), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT73), .ZN(new_n311_));
  OR2_X1    g110(.A1(new_n305_), .A2(new_n306_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT36), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n312_), .A2(new_n313_), .A3(new_n307_), .ZN(new_n314_));
  AND3_X1   g113(.A1(new_n310_), .A2(new_n311_), .A3(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n311_), .B1(new_n310_), .B2(new_n314_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G29gat), .B(G36gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G43gat), .B(G50gat), .ZN(new_n319_));
  OR2_X1    g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n319_), .ZN(new_n321_));
  AND2_X1   g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  OAI211_X1 g121(.A(new_n322_), .B(new_n220_), .C1(new_n247_), .C2(new_n248_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n320_), .A2(KEYINPUT15), .A3(new_n321_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(KEYINPUT15), .B1(new_n320_), .B2(new_n321_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n323_), .B1(new_n327_), .B2(new_n237_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT71), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n330_));
  AND2_X1   g129(.A1(G232gat), .A2(G233gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  AND2_X1   g131(.A1(new_n332_), .A2(KEYINPUT35), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n332_), .A2(KEYINPUT35), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n328_), .A2(new_n329_), .A3(new_n335_), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n323_), .B(new_n333_), .C1(new_n327_), .C2(new_n237_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n329_), .B1(new_n328_), .B2(new_n335_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n317_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(KEYINPUT74), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n328_), .A2(new_n335_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT71), .ZN(new_n343_));
  INV_X1    g142(.A(new_n314_), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n343_), .A2(new_n337_), .A3(new_n336_), .A4(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT72), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT74), .ZN(new_n348_));
  OAI211_X1 g147(.A(new_n348_), .B(new_n317_), .C1(new_n338_), .C2(new_n339_), .ZN(new_n349_));
  AND2_X1   g148(.A1(new_n336_), .A2(new_n337_), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n350_), .A2(KEYINPUT72), .A3(new_n343_), .A4(new_n344_), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n341_), .A2(new_n347_), .A3(new_n349_), .A4(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(KEYINPUT37), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT76), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n343_), .A2(new_n337_), .A3(new_n336_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT75), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT75), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n350_), .A2(new_n357_), .A3(new_n343_), .ZN(new_n358_));
  AND2_X1   g157(.A1(new_n310_), .A2(new_n314_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n356_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT37), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n360_), .A2(new_n361_), .A3(new_n345_), .ZN(new_n362_));
  AND3_X1   g161(.A1(new_n353_), .A2(new_n354_), .A3(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n354_), .B1(new_n353_), .B2(new_n362_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n279_), .B(new_n303_), .C1(new_n363_), .C2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT97), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT85), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G141gat), .A2(G148gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT81), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT81), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n370_), .A2(G141gat), .A3(G148gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n369_), .A2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(KEYINPUT84), .B(KEYINPUT2), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  AND3_X1   g173(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT3), .ZN(new_n377_));
  NOR3_X1   g176(.A1(new_n377_), .A2(G141gat), .A3(G148gat), .ZN(new_n378_));
  INV_X1    g177(.A(G141gat), .ZN(new_n379_));
  INV_X1    g178(.A(G148gat), .ZN(new_n380_));
  AOI21_X1  g179(.A(KEYINPUT3), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n376_), .B1(new_n378_), .B2(new_n381_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n367_), .B1(new_n374_), .B2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT2), .ZN(new_n384_));
  AND2_X1   g183(.A1(new_n384_), .A2(KEYINPUT84), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n384_), .A2(KEYINPUT84), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n369_), .B(new_n371_), .C1(new_n385_), .C2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n379_), .A2(new_n380_), .A3(KEYINPUT3), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n377_), .B1(G141gat), .B2(G148gat), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n375_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n387_), .A2(KEYINPUT85), .A3(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(G155gat), .ZN(new_n392_));
  INV_X1    g191(.A(G162gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G155gat), .A2(G162gat), .ZN(new_n395_));
  AND3_X1   g194(.A1(new_n394_), .A2(KEYINPUT86), .A3(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(KEYINPUT86), .B1(new_n394_), .B2(new_n395_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n383_), .A2(new_n391_), .A3(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n379_), .A2(new_n380_), .A3(KEYINPUT82), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT82), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n401_), .B1(G141gat), .B2(G148gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT1), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n394_), .A2(new_n404_), .A3(new_n395_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n369_), .A2(new_n371_), .A3(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(KEYINPUT83), .B1(new_n406_), .B2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n408_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT83), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n410_), .A2(new_n411_), .A3(new_n403_), .A4(new_n405_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n409_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n399_), .A2(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n414_), .A2(KEYINPUT29), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G22gat), .B(G50gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT28), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n415_), .B(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G78gat), .B(G106gat), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  OR2_X1    g219(.A1(G197gat), .A2(G204gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G197gat), .A2(G204gat), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n421_), .A2(KEYINPUT21), .A3(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT21), .ZN(new_n424_));
  AND2_X1   g223(.A1(G197gat), .A2(G204gat), .ZN(new_n425_));
  NOR2_X1   g224(.A1(G197gat), .A2(G204gat), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n424_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G211gat), .B(G218gat), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n423_), .A2(new_n427_), .A3(KEYINPUT87), .A4(new_n428_), .ZN(new_n429_));
  AND3_X1   g228(.A1(new_n423_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT87), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n431_), .B1(new_n423_), .B2(new_n428_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n429_), .B1(new_n430_), .B2(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n433_), .B1(new_n414_), .B2(KEYINPUT29), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G228gat), .A2(G233gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n435_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT29), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n438_), .B1(new_n399_), .B2(new_n413_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n437_), .B1(new_n439_), .B2(new_n433_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n420_), .B1(new_n436_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT88), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n418_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n440_), .ZN(new_n444_));
  NOR3_X1   g243(.A1(new_n439_), .A2(new_n437_), .A3(new_n433_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n419_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n436_), .A2(new_n440_), .A3(new_n420_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n443_), .A2(new_n448_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n446_), .A2(new_n418_), .A3(new_n442_), .A4(new_n447_), .ZN(new_n450_));
  AND2_X1   g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G1gat), .B(G29gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n452_), .B(G85gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(KEYINPUT0), .B(G57gat), .ZN(new_n454_));
  XOR2_X1   g253(.A(new_n453_), .B(new_n454_), .Z(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  XOR2_X1   g255(.A(G127gat), .B(G134gat), .Z(new_n457_));
  XOR2_X1   g256(.A(G113gat), .B(G120gat), .Z(new_n458_));
  XNOR2_X1  g257(.A(new_n457_), .B(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n391_), .A2(new_n398_), .ZN(new_n461_));
  AOI21_X1  g260(.A(KEYINPUT85), .B1(new_n387_), .B2(new_n390_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  AND2_X1   g262(.A1(new_n409_), .A2(new_n412_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n460_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n399_), .A2(new_n459_), .A3(new_n413_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n465_), .A2(KEYINPUT4), .A3(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G225gat), .A2(G233gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(KEYINPUT90), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n469_), .B(KEYINPUT91), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n459_), .B1(new_n399_), .B2(new_n413_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT4), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n471_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n465_), .A2(new_n466_), .A3(new_n469_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT92), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT92), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n465_), .A2(new_n477_), .A3(new_n466_), .A4(new_n469_), .ZN(new_n478_));
  AOI221_X4 g277(.A(new_n456_), .B1(new_n467_), .B2(new_n474_), .C1(new_n476_), .C2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n476_), .A2(new_n478_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n467_), .A2(new_n474_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n455_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n479_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G226gat), .A2(G233gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(KEYINPUT19), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT24), .ZN(new_n486_));
  INV_X1    g285(.A(G169gat), .ZN(new_n487_));
  INV_X1    g286(.A(G176gat), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n486_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G169gat), .A2(G176gat), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  OAI21_X1  g290(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n489_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G183gat), .A2(G190gat), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT23), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n493_), .A2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(KEYINPUT26), .B(G190gat), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT80), .ZN(new_n501_));
  INV_X1    g300(.A(G183gat), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n501_), .B1(new_n502_), .B2(KEYINPUT25), .ZN(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT25), .B(G183gat), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n500_), .B(new_n503_), .C1(new_n504_), .C2(new_n501_), .ZN(new_n505_));
  INV_X1    g304(.A(G190gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n502_), .A2(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n496_), .A2(new_n497_), .A3(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT22), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n509_), .A2(new_n488_), .A3(G169gat), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n487_), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  AOI22_X1  g311(.A1(new_n499_), .A2(new_n505_), .B1(new_n508_), .B2(new_n512_), .ZN(new_n513_));
  OAI21_X1  g312(.A(KEYINPUT20), .B1(new_n433_), .B2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n504_), .A2(new_n500_), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n496_), .A2(new_n497_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n487_), .A2(new_n488_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n517_), .A2(KEYINPUT24), .A3(new_n490_), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n515_), .A2(new_n516_), .A3(new_n518_), .A4(new_n489_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n508_), .A2(new_n512_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n423_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n522_), .B(new_n431_), .C1(new_n423_), .C2(new_n428_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n521_), .B1(new_n523_), .B2(new_n429_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n485_), .B1(new_n514_), .B2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(KEYINPUT95), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT95), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n527_), .B(new_n485_), .C1(new_n514_), .C2(new_n524_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT20), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n529_), .B1(new_n433_), .B2(new_n513_), .ZN(new_n530_));
  AND3_X1   g329(.A1(new_n508_), .A2(new_n512_), .A3(KEYINPUT89), .ZN(new_n531_));
  AOI21_X1  g330(.A(KEYINPUT89), .B1(new_n508_), .B2(new_n512_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n519_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n533_), .A2(new_n523_), .A3(new_n429_), .ZN(new_n534_));
  AND2_X1   g333(.A1(new_n530_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n485_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n526_), .A2(new_n528_), .A3(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G8gat), .B(G36gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT18), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G64gat), .B(G92gat), .ZN(new_n541_));
  XOR2_X1   g340(.A(new_n540_), .B(new_n541_), .Z(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n538_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT27), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT89), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n520_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n508_), .A2(new_n512_), .A3(KEYINPUT89), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n433_), .A2(new_n519_), .A3(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  OAI211_X1 g350(.A(KEYINPUT20), .B(new_n536_), .C1(new_n433_), .C2(new_n513_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n536_), .B1(new_n530_), .B2(new_n534_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n545_), .B1(new_n555_), .B2(new_n542_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n544_), .A2(new_n556_), .ZN(new_n557_));
  OR2_X1    g356(.A1(new_n433_), .A2(new_n513_), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n558_), .A2(new_n550_), .A3(KEYINPUT20), .A4(new_n536_), .ZN(new_n559_));
  OAI211_X1 g358(.A(new_n559_), .B(new_n542_), .C1(new_n535_), .C2(new_n536_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n543_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(new_n545_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n557_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n451_), .A2(new_n483_), .A3(new_n565_), .ZN(new_n566_));
  AND3_X1   g365(.A1(new_n399_), .A2(new_n459_), .A3(new_n413_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n567_), .A2(new_n472_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n477_), .B1(new_n568_), .B2(new_n469_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n478_), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n481_), .B(new_n455_), .C1(new_n569_), .C2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT33), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n455_), .A2(KEYINPUT33), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n574_), .B1(new_n467_), .B2(new_n474_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n562_), .B1(new_n480_), .B2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n472_), .A2(new_n473_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n467_), .A2(new_n469_), .A3(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT94), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n465_), .A2(new_n466_), .A3(new_n470_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(new_n456_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(KEYINPUT93), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n467_), .A2(KEYINPUT94), .A3(new_n469_), .A4(new_n577_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT93), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n581_), .A2(new_n585_), .A3(new_n456_), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n580_), .A2(new_n583_), .A3(new_n584_), .A4(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n573_), .A2(new_n576_), .A3(new_n587_), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n542_), .A2(KEYINPUT32), .ZN(new_n589_));
  NOR3_X1   g388(.A1(new_n589_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n590_), .B1(new_n538_), .B2(new_n589_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n591_), .B1(new_n479_), .B2(new_n482_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n588_), .A2(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n566_), .B1(new_n593_), .B2(new_n451_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G71gat), .B(G99gat), .ZN(new_n595_));
  INV_X1    g394(.A(G43gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n513_), .B(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(new_n459_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(G227gat), .A2(G233gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(new_n285_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT30), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT31), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n599_), .B(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(KEYINPUT96), .B1(new_n594_), .B2(new_n605_), .ZN(new_n606_));
  AOI22_X1  g405(.A1(new_n588_), .A2(new_n592_), .B1(new_n450_), .B2(new_n449_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n480_), .A2(new_n481_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(new_n456_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n609_), .A2(new_n557_), .A3(new_n571_), .A4(new_n563_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n449_), .A2(new_n450_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  OAI211_X1 g411(.A(KEYINPUT96), .B(new_n605_), .C1(new_n607_), .C2(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n451_), .A2(new_n564_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n614_), .A2(new_n604_), .A3(new_n483_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n613_), .A2(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n606_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT79), .ZN(new_n618_));
  INV_X1    g417(.A(new_n326_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(new_n324_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n618_), .B1(new_n293_), .B2(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n284_), .B(new_n290_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n327_), .A2(new_n622_), .A3(KEYINPUT79), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(G229gat), .A2(G233gat), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n320_), .A2(new_n321_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n626_), .B1(new_n293_), .B2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n293_), .A2(new_n627_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n622_), .A2(new_n322_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  AOI22_X1  g430(.A1(new_n624_), .A2(new_n628_), .B1(new_n631_), .B2(new_n626_), .ZN(new_n632_));
  XOR2_X1   g431(.A(G113gat), .B(G141gat), .Z(new_n633_));
  XNOR2_X1  g432(.A(G169gat), .B(G197gat), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n632_), .B(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n366_), .B1(new_n617_), .B2(new_n637_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n605_), .B1(new_n607_), .B2(new_n612_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT96), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n641_), .A2(new_n615_), .A3(new_n613_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n642_), .A2(KEYINPUT97), .A3(new_n636_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n365_), .B1(new_n638_), .B2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(G1gat), .ZN(new_n645_));
  INV_X1    g444(.A(new_n483_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n644_), .A2(new_n645_), .A3(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT38), .ZN(new_n648_));
  OR2_X1    g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n360_), .A2(new_n345_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n617_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n279_), .A2(new_n636_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n303_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n652_), .A2(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(G1gat), .B1(new_n656_), .B2(new_n483_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n647_), .A2(new_n648_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n649_), .A2(new_n657_), .A3(new_n658_), .ZN(G1324gat));
  INV_X1    g458(.A(KEYINPUT40), .ZN(new_n660_));
  OAI21_X1  g459(.A(G8gat), .B1(new_n656_), .B2(new_n565_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT98), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  OAI211_X1 g462(.A(KEYINPUT98), .B(G8gat), .C1(new_n656_), .C2(new_n565_), .ZN(new_n664_));
  AND3_X1   g463(.A1(new_n663_), .A2(KEYINPUT39), .A3(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT39), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n661_), .A2(new_n662_), .A3(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(G8gat), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n644_), .A2(new_n668_), .A3(new_n564_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n660_), .B1(new_n665_), .B2(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n663_), .A2(KEYINPUT39), .A3(new_n664_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n672_), .A2(KEYINPUT40), .A3(new_n667_), .A4(new_n669_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n671_), .A2(new_n673_), .ZN(G1325gat));
  OAI21_X1  g473(.A(G15gat), .B1(new_n656_), .B2(new_n605_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(KEYINPUT99), .B(KEYINPUT41), .ZN(new_n676_));
  OR2_X1    g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n644_), .A2(new_n285_), .A3(new_n604_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n675_), .A2(new_n676_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n677_), .A2(new_n678_), .A3(new_n679_), .ZN(G1326gat));
  NAND3_X1  g479(.A1(new_n652_), .A2(new_n451_), .A3(new_n655_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(G22gat), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(KEYINPUT100), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT100), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n681_), .A2(new_n684_), .A3(G22gat), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n683_), .A2(KEYINPUT42), .A3(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n644_), .A2(new_n286_), .A3(new_n451_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(KEYINPUT42), .B1(new_n683_), .B2(new_n685_), .ZN(new_n689_));
  OR2_X1    g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1327gat));
  NOR2_X1   g489(.A1(new_n653_), .A2(new_n303_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT43), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n363_), .A2(new_n364_), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n692_), .B(new_n693_), .C1(new_n606_), .C2(new_n616_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n692_), .B1(new_n642_), .B2(new_n693_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n691_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  OAI211_X1 g498(.A(KEYINPUT44), .B(new_n691_), .C1(new_n695_), .C2(new_n696_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  OAI21_X1  g500(.A(G29gat), .B1(new_n701_), .B2(new_n483_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n638_), .A2(new_n643_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n279_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n650_), .A2(new_n303_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n704_), .A2(new_n706_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n483_), .A2(G29gat), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT101), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n703_), .A2(new_n707_), .A3(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n702_), .A2(new_n710_), .ZN(G1328gat));
  XNOR2_X1  g510(.A(KEYINPUT102), .B(KEYINPUT46), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n565_), .A2(G36gat), .ZN(new_n714_));
  INV_X1    g513(.A(new_n643_), .ZN(new_n715_));
  AOI21_X1  g514(.A(KEYINPUT97), .B1(new_n642_), .B2(new_n636_), .ZN(new_n716_));
  OAI211_X1 g515(.A(new_n707_), .B(new_n714_), .C1(new_n715_), .C2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(KEYINPUT45), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT45), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n703_), .A2(new_n719_), .A3(new_n707_), .A4(new_n714_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n699_), .A2(new_n564_), .A3(new_n700_), .ZN(new_n721_));
  AOI221_X4 g520(.A(new_n713_), .B1(new_n718_), .B2(new_n720_), .C1(new_n721_), .C2(G36gat), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(G36gat), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n718_), .A2(new_n720_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n712_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n722_), .A2(new_n725_), .ZN(G1329gat));
  NAND2_X1  g525(.A1(new_n604_), .A2(G43gat), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n703_), .A2(new_n604_), .A3(new_n707_), .ZN(new_n728_));
  OAI22_X1  g527(.A1(new_n701_), .A2(new_n727_), .B1(new_n728_), .B2(G43gat), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g529(.A1(new_n451_), .A2(G50gat), .ZN(new_n731_));
  AND3_X1   g530(.A1(new_n703_), .A2(new_n451_), .A3(new_n707_), .ZN(new_n732_));
  OAI22_X1  g531(.A1(new_n701_), .A2(new_n731_), .B1(new_n732_), .B2(G50gat), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT103), .ZN(G1331gat));
  OAI21_X1  g533(.A(KEYINPUT104), .B1(new_n617_), .B2(new_n636_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT104), .ZN(new_n736_));
  OAI211_X1 g535(.A(new_n736_), .B(new_n637_), .C1(new_n606_), .C2(new_n616_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n353_), .A2(new_n362_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(KEYINPUT76), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n353_), .A2(new_n354_), .A3(new_n362_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n654_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  AND3_X1   g541(.A1(new_n738_), .A2(new_n704_), .A3(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT105), .ZN(new_n744_));
  OR2_X1    g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n744_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n483_), .A2(G57gat), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n745_), .A2(new_n746_), .A3(new_n747_), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n652_), .A2(new_n637_), .A3(new_n704_), .A4(new_n303_), .ZN(new_n749_));
  OAI21_X1  g548(.A(G57gat), .B1(new_n749_), .B2(new_n483_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n750_), .ZN(G1332gat));
  NOR2_X1   g550(.A1(new_n565_), .A2(G64gat), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n745_), .A2(new_n746_), .A3(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(G64gat), .B1(new_n749_), .B2(new_n565_), .ZN(new_n754_));
  XOR2_X1   g553(.A(KEYINPUT106), .B(KEYINPUT48), .Z(new_n755_));
  XNOR2_X1  g554(.A(new_n754_), .B(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n753_), .A2(new_n756_), .ZN(G1333gat));
  NOR2_X1   g556(.A1(new_n605_), .A2(G71gat), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n745_), .A2(new_n746_), .A3(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(G71gat), .B1(new_n749_), .B2(new_n605_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT49), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(G1334gat));
  NOR2_X1   g561(.A1(new_n611_), .A2(G78gat), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n745_), .A2(new_n746_), .A3(new_n763_), .ZN(new_n764_));
  OAI21_X1  g563(.A(G78gat), .B1(new_n749_), .B2(new_n611_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT50), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(G1335gat));
  NOR2_X1   g566(.A1(new_n279_), .A2(new_n706_), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n738_), .A2(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n769_), .A2(new_n216_), .A3(new_n646_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n636_), .A2(new_n303_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n704_), .A2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT107), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n772_), .B(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n696_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n776_), .B2(new_n694_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n777_), .A2(new_n646_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n770_), .B1(new_n778_), .B2(new_n216_), .ZN(G1336gat));
  NAND3_X1  g578(.A1(new_n769_), .A2(new_n217_), .A3(new_n564_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n777_), .A2(new_n564_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n780_), .B1(new_n781_), .B2(new_n217_), .ZN(G1337gat));
  AND3_X1   g581(.A1(new_n604_), .A2(new_n212_), .A3(new_n214_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n769_), .A2(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n226_), .B1(new_n777_), .B2(new_n604_), .ZN(new_n785_));
  OR3_X1    g584(.A1(new_n784_), .A2(new_n785_), .A3(KEYINPUT51), .ZN(new_n786_));
  OAI21_X1  g585(.A(KEYINPUT51), .B1(new_n784_), .B2(new_n785_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(G1338gat));
  OAI211_X1 g587(.A(new_n451_), .B(new_n774_), .C1(new_n695_), .C2(new_n696_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT109), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n789_), .A2(new_n790_), .A3(G106gat), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(KEYINPUT52), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n790_), .B1(new_n789_), .B2(G106gat), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n789_), .A2(G106gat), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n795_), .A2(KEYINPUT109), .A3(new_n796_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n611_), .A2(G106gat), .ZN(new_n798_));
  INV_X1    g597(.A(new_n737_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n736_), .B1(new_n642_), .B2(new_n637_), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n768_), .B(new_n798_), .C1(new_n799_), .C2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT108), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n738_), .A2(KEYINPUT108), .A3(new_n768_), .A4(new_n798_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n797_), .A2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(KEYINPUT53), .B1(new_n794_), .B2(new_n806_), .ZN(new_n807_));
  AOI22_X1  g606(.A1(new_n793_), .A2(new_n796_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n808_), .B(new_n809_), .C1(new_n793_), .C2(new_n792_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n807_), .A2(new_n810_), .ZN(G1339gat));
  NAND3_X1  g610(.A1(new_n614_), .A2(new_n604_), .A3(new_n646_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT58), .ZN(new_n813_));
  AND3_X1   g612(.A1(new_n273_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n632_), .A2(new_n635_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n624_), .A2(new_n629_), .A3(new_n626_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n635_), .B1(new_n631_), .B2(new_n625_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n815_), .A2(new_n818_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n814_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n269_), .A2(new_n821_), .A3(new_n270_), .ZN(new_n822_));
  AND3_X1   g621(.A1(new_n262_), .A2(new_n264_), .A3(new_n266_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n262_), .A2(new_n251_), .A3(new_n246_), .A4(new_n266_), .ZN(new_n824_));
  AOI22_X1  g623(.A1(new_n823_), .A2(KEYINPUT55), .B1(new_n824_), .B2(new_n263_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n276_), .B1(new_n822_), .B2(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(KEYINPUT112), .B1(new_n826_), .B2(KEYINPUT56), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT56), .ZN(new_n828_));
  AOI211_X1 g627(.A(new_n828_), .B(new_n276_), .C1(new_n822_), .C2(new_n825_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n820_), .B1(new_n827_), .B2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n822_), .A2(new_n825_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n205_), .ZN(new_n832_));
  NOR3_X1   g631(.A1(new_n832_), .A2(KEYINPUT112), .A3(new_n828_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n813_), .B1(new_n830_), .B2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n832_), .A2(new_n828_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n826_), .A2(KEYINPUT56), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n835_), .A2(KEYINPUT112), .A3(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n827_), .A2(new_n829_), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n837_), .A2(new_n838_), .A3(KEYINPUT58), .A4(new_n820_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n834_), .A2(new_n740_), .A3(new_n839_), .A4(new_n741_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n650_), .A2(KEYINPUT57), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT110), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n832_), .A2(new_n843_), .A3(new_n828_), .ZN(new_n844_));
  OAI21_X1  g643(.A(KEYINPUT110), .B1(new_n826_), .B2(KEYINPUT56), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n844_), .A2(new_n836_), .A3(new_n845_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n637_), .A2(new_n814_), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n819_), .ZN(new_n849_));
  AOI21_X1  g648(.A(KEYINPUT111), .B1(new_n278_), .B2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT111), .ZN(new_n851_));
  AOI211_X1 g650(.A(new_n851_), .B(new_n819_), .C1(new_n272_), .C2(new_n277_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n850_), .A2(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n842_), .B1(new_n848_), .B2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n276_), .B1(new_n273_), .B2(new_n275_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n849_), .B1(new_n814_), .B2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n851_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n278_), .A2(KEYINPUT111), .A3(new_n849_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n846_), .A2(new_n847_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n651_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n840_), .B(new_n854_), .C1(KEYINPUT57), .C2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n654_), .ZN(new_n863_));
  OAI21_X1  g662(.A(KEYINPUT54), .B1(new_n365_), .B2(new_n636_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n742_), .A2(new_n865_), .A3(new_n637_), .A4(new_n279_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n864_), .A2(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n812_), .B1(new_n863_), .B2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT113), .ZN(new_n869_));
  AOI21_X1  g668(.A(KEYINPUT59), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  AOI22_X1  g669(.A1(new_n862_), .A2(new_n654_), .B1(new_n864_), .B2(new_n866_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT59), .ZN(new_n872_));
  NOR4_X1   g671(.A1(new_n871_), .A2(KEYINPUT113), .A3(new_n872_), .A4(new_n812_), .ZN(new_n873_));
  OAI21_X1  g672(.A(KEYINPUT114), .B1(new_n870_), .B2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n812_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n841_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n650_), .B1(new_n848_), .B2(new_n853_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n876_), .B1(new_n877_), .B2(new_n878_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n303_), .B1(new_n879_), .B2(new_n840_), .ZN(new_n880_));
  AND2_X1   g679(.A1(new_n864_), .A2(new_n866_), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n869_), .B(new_n875_), .C1(new_n880_), .C2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(new_n872_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT114), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n868_), .A2(new_n869_), .A3(KEYINPUT59), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n883_), .A2(new_n884_), .A3(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT115), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n636_), .A2(new_n887_), .A3(G113gat), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n888_), .B1(new_n887_), .B2(G113gat), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n874_), .A2(new_n886_), .A3(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(G113gat), .ZN(new_n891_));
  INV_X1    g690(.A(new_n868_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n892_), .B2(new_n637_), .ZN(new_n893_));
  AND2_X1   g692(.A1(new_n890_), .A2(new_n893_), .ZN(G1340gat));
  INV_X1    g693(.A(G120gat), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n895_), .B1(new_n279_), .B2(KEYINPUT60), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n868_), .B(new_n896_), .C1(KEYINPUT60), .C2(new_n895_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n279_), .B1(new_n883_), .B2(new_n885_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n898_), .B2(new_n895_), .ZN(G1341gat));
  INV_X1    g698(.A(G127gat), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n654_), .A2(new_n900_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n874_), .A2(new_n886_), .A3(new_n901_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n900_), .B1(new_n892_), .B2(new_n654_), .ZN(new_n903_));
  AND2_X1   g702(.A1(new_n902_), .A2(new_n903_), .ZN(G1342gat));
  INV_X1    g703(.A(new_n693_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(KEYINPUT116), .B(G134gat), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n874_), .A2(new_n886_), .A3(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(G134gat), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n909_), .B1(new_n892_), .B2(new_n650_), .ZN(new_n910_));
  AND2_X1   g709(.A1(new_n908_), .A2(new_n910_), .ZN(G1343gat));
  INV_X1    g710(.A(new_n871_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n451_), .A2(new_n605_), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n913_), .A2(new_n483_), .A3(new_n564_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n912_), .A2(new_n914_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n915_), .A2(new_n637_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(new_n379_), .ZN(G1344gat));
  NOR2_X1   g716(.A1(new_n915_), .A2(new_n279_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(new_n380_), .ZN(G1345gat));
  AND2_X1   g718(.A1(new_n912_), .A2(new_n914_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT117), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n920_), .A2(new_n921_), .A3(new_n303_), .ZN(new_n922_));
  OAI21_X1  g721(.A(KEYINPUT117), .B1(new_n915_), .B2(new_n654_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(KEYINPUT61), .B(G155gat), .ZN(new_n924_));
  AND3_X1   g723(.A1(new_n922_), .A2(new_n923_), .A3(new_n924_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n924_), .B1(new_n922_), .B2(new_n923_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n925_), .A2(new_n926_), .ZN(G1346gat));
  NAND3_X1  g726(.A1(new_n920_), .A2(new_n393_), .A3(new_n651_), .ZN(new_n928_));
  OAI21_X1  g727(.A(G162gat), .B1(new_n915_), .B2(new_n905_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(G1347gat));
  NOR2_X1   g729(.A1(new_n871_), .A2(new_n451_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n646_), .A2(new_n565_), .ZN(new_n932_));
  INV_X1    g731(.A(new_n932_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n933_), .A2(new_n605_), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n931_), .A2(new_n636_), .A3(new_n934_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT62), .ZN(new_n936_));
  AND3_X1   g735(.A1(new_n935_), .A2(new_n936_), .A3(G169gat), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n936_), .B1(new_n935_), .B2(G169gat), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n931_), .A2(new_n934_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(KEYINPUT22), .B(G169gat), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n636_), .A2(new_n940_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(KEYINPUT118), .ZN(new_n942_));
  OAI22_X1  g741(.A1(new_n937_), .A2(new_n938_), .B1(new_n939_), .B2(new_n942_), .ZN(G1348gat));
  INV_X1    g742(.A(KEYINPUT119), .ZN(new_n944_));
  NAND3_X1  g743(.A1(new_n912_), .A2(new_n944_), .A3(new_n611_), .ZN(new_n945_));
  OAI21_X1  g744(.A(KEYINPUT119), .B1(new_n871_), .B2(new_n451_), .ZN(new_n946_));
  AND2_X1   g745(.A1(new_n945_), .A2(new_n946_), .ZN(new_n947_));
  INV_X1    g746(.A(new_n934_), .ZN(new_n948_));
  NOR3_X1   g747(.A1(new_n948_), .A2(new_n488_), .A3(new_n279_), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n931_), .A2(new_n704_), .A3(new_n934_), .ZN(new_n950_));
  AOI22_X1  g749(.A1(new_n947_), .A2(new_n949_), .B1(new_n950_), .B2(new_n488_), .ZN(G1349gat));
  NOR3_X1   g750(.A1(new_n939_), .A2(new_n504_), .A3(new_n654_), .ZN(new_n952_));
  INV_X1    g751(.A(KEYINPUT120), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n948_), .A2(new_n654_), .ZN(new_n954_));
  NAND4_X1  g753(.A1(new_n945_), .A2(new_n946_), .A3(new_n953_), .A4(new_n954_), .ZN(new_n955_));
  AND2_X1   g754(.A1(new_n955_), .A2(new_n502_), .ZN(new_n956_));
  NAND3_X1  g755(.A1(new_n945_), .A2(new_n946_), .A3(new_n954_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n957_), .A2(KEYINPUT120), .ZN(new_n958_));
  AOI21_X1  g757(.A(new_n952_), .B1(new_n956_), .B2(new_n958_), .ZN(G1350gat));
  NAND2_X1  g758(.A1(new_n651_), .A2(new_n500_), .ZN(new_n960_));
  XOR2_X1   g759(.A(new_n960_), .B(KEYINPUT121), .Z(new_n961_));
  NOR4_X1   g760(.A1(new_n871_), .A2(new_n451_), .A3(new_n905_), .A4(new_n948_), .ZN(new_n962_));
  OAI22_X1  g761(.A1(new_n939_), .A2(new_n961_), .B1(new_n962_), .B2(new_n506_), .ZN(new_n963_));
  XNOR2_X1  g762(.A(new_n963_), .B(KEYINPUT122), .ZN(G1351gat));
  NOR3_X1   g763(.A1(new_n871_), .A2(new_n913_), .A3(new_n933_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n965_), .A2(new_n636_), .ZN(new_n966_));
  INV_X1    g765(.A(G197gat), .ZN(new_n967_));
  AOI21_X1  g766(.A(new_n966_), .B1(KEYINPUT123), .B2(new_n967_), .ZN(new_n968_));
  XOR2_X1   g767(.A(KEYINPUT123), .B(G197gat), .Z(new_n969_));
  AOI21_X1  g768(.A(new_n968_), .B1(new_n966_), .B2(new_n969_), .ZN(G1352gat));
  AOI21_X1  g769(.A(new_n279_), .B1(KEYINPUT124), .B2(G204gat), .ZN(new_n971_));
  NAND2_X1  g770(.A1(new_n965_), .A2(new_n971_), .ZN(new_n972_));
  NOR2_X1   g771(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n973_));
  XNOR2_X1  g772(.A(new_n973_), .B(KEYINPUT125), .ZN(new_n974_));
  XNOR2_X1  g773(.A(new_n972_), .B(new_n974_), .ZN(G1353gat));
  NAND2_X1  g774(.A1(new_n965_), .A2(new_n303_), .ZN(new_n976_));
  OAI21_X1  g775(.A(new_n976_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n977_));
  XOR2_X1   g776(.A(KEYINPUT63), .B(G211gat), .Z(new_n978_));
  OAI21_X1  g777(.A(new_n977_), .B1(new_n976_), .B2(new_n978_), .ZN(G1354gat));
  XOR2_X1   g778(.A(KEYINPUT126), .B(G218gat), .Z(new_n980_));
  INV_X1    g779(.A(new_n980_), .ZN(new_n981_));
  AND3_X1   g780(.A1(new_n965_), .A2(new_n693_), .A3(new_n981_), .ZN(new_n982_));
  AOI21_X1  g781(.A(new_n981_), .B1(new_n965_), .B2(new_n651_), .ZN(new_n983_));
  OR3_X1    g782(.A1(new_n982_), .A2(new_n983_), .A3(KEYINPUT127), .ZN(new_n984_));
  OAI21_X1  g783(.A(KEYINPUT127), .B1(new_n982_), .B2(new_n983_), .ZN(new_n985_));
  NAND2_X1  g784(.A1(new_n984_), .A2(new_n985_), .ZN(G1355gat));
endmodule


