//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 1 0 1 0 1 1 1 1 1 1 0 0 1 0 0 0 0 1 0 1 1 0 0 1 1 0 1 1 1 0 1 0 1 1 0 0 1 1 1 0 0 0 1 1 0 1 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n711_, new_n712_, new_n713_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n837_, new_n838_,
    new_n840_, new_n841_, new_n843_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n875_, new_n876_,
    new_n877_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_, new_n913_;
  INV_X1    g000(.A(KEYINPUT8), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT7), .ZN(new_n203_));
  INV_X1    g002(.A(G99gat), .ZN(new_n204_));
  INV_X1    g003(.A(G106gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT6), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n211_));
  NAND4_X1  g010(.A1(new_n206_), .A2(new_n209_), .A3(new_n210_), .A4(new_n211_), .ZN(new_n212_));
  XOR2_X1   g011(.A(G85gat), .B(G92gat), .Z(new_n213_));
  AOI21_X1  g012(.A(new_n202_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT66), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT65), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n212_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(new_n202_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n213_), .B1(new_n212_), .B2(new_n216_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n215_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  AOI21_X1  g019(.A(KEYINPUT8), .B1(new_n212_), .B2(new_n216_), .ZN(new_n221_));
  AND2_X1   g020(.A1(new_n209_), .A2(new_n210_), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n222_), .A2(KEYINPUT65), .A3(new_n211_), .A4(new_n206_), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n221_), .A2(new_n223_), .A3(KEYINPUT66), .A4(new_n213_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n214_), .B1(new_n220_), .B2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(G85gat), .ZN(new_n226_));
  INV_X1    g025(.A(G92gat), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT64), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT9), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT9), .ZN(new_n230_));
  OAI211_X1 g029(.A(KEYINPUT64), .B(new_n230_), .C1(new_n226_), .C2(new_n227_), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n229_), .B(new_n231_), .C1(G85gat), .C2(G92gat), .ZN(new_n232_));
  XOR2_X1   g031(.A(KEYINPUT10), .B(G99gat), .Z(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(new_n205_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n232_), .A2(new_n222_), .A3(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(G71gat), .ZN(new_n237_));
  INV_X1    g036(.A(G78gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G71gat), .A2(G78gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G57gat), .B(G64gat), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n239_), .B(new_n240_), .C1(new_n241_), .C2(KEYINPUT11), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT67), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT68), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n247_), .B1(KEYINPUT11), .B2(new_n241_), .ZN(new_n248_));
  AND2_X1   g047(.A1(G57gat), .A2(G64gat), .ZN(new_n249_));
  NOR2_X1   g048(.A1(G57gat), .A2(G64gat), .ZN(new_n250_));
  OAI21_X1  g049(.A(KEYINPUT11), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT67), .B(KEYINPUT68), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n242_), .B1(new_n248_), .B2(new_n253_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n249_), .A2(new_n250_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT11), .ZN(new_n256_));
  AOI22_X1  g055(.A1(new_n255_), .A2(new_n256_), .B1(G71gat), .B2(G78gat), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n247_), .A2(new_n241_), .A3(KEYINPUT11), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n251_), .A2(new_n252_), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n257_), .A2(new_n258_), .A3(new_n259_), .A4(new_n239_), .ZN(new_n260_));
  AND3_X1   g059(.A1(new_n254_), .A2(new_n260_), .A3(KEYINPUT69), .ZN(new_n261_));
  AOI21_X1  g060(.A(KEYINPUT69), .B1(new_n254_), .B2(new_n260_), .ZN(new_n262_));
  OAI22_X1  g061(.A1(new_n225_), .A2(new_n236_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT12), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(KEYINPUT73), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT73), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n263_), .A2(new_n267_), .A3(new_n264_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n266_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT72), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n220_), .A2(new_n224_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n214_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n235_), .A2(KEYINPUT70), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT70), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n232_), .A2(new_n274_), .A3(new_n222_), .A4(new_n234_), .ZN(new_n275_));
  AOI22_X1  g074(.A1(new_n271_), .A2(new_n272_), .B1(new_n273_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n254_), .A2(new_n260_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n254_), .A2(new_n260_), .A3(KEYINPUT71), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n279_), .A2(KEYINPUT12), .A3(new_n280_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n270_), .B1(new_n276_), .B2(new_n281_), .ZN(new_n282_));
  AND3_X1   g081(.A1(new_n254_), .A2(new_n260_), .A3(KEYINPUT71), .ZN(new_n283_));
  AOI21_X1  g082(.A(KEYINPUT71), .B1(new_n254_), .B2(new_n260_), .ZN(new_n284_));
  NOR3_X1   g083(.A1(new_n283_), .A2(new_n284_), .A3(new_n264_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n273_), .A2(new_n275_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n285_), .B(KEYINPUT72), .C1(new_n225_), .C2(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n236_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n261_), .A2(new_n262_), .ZN(new_n290_));
  AOI22_X1  g089(.A1(new_n282_), .A2(new_n288_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G230gat), .A2(G233gat), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n269_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n289_), .A2(new_n290_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(new_n263_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n292_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n293_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT74), .B(KEYINPUT5), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G176gat), .B(G204gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G120gat), .B(G148gat), .ZN(new_n302_));
  XOR2_X1   g101(.A(new_n301_), .B(new_n302_), .Z(new_n303_));
  NAND2_X1  g102(.A1(new_n298_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n303_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n293_), .A2(new_n297_), .A3(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT13), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n304_), .A2(KEYINPUT13), .A3(new_n306_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT83), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT26), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n312_), .B1(new_n313_), .B2(G190gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(KEYINPUT25), .B(G183gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT26), .B(G190gat), .ZN(new_n316_));
  OAI211_X1 g115(.A(new_n314_), .B(new_n315_), .C1(new_n316_), .C2(new_n312_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G169gat), .A2(G176gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT84), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  OAI21_X1  g119(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n317_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT85), .ZN(new_n323_));
  OR2_X1    g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NOR3_X1   g123(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n325_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G183gat), .A2(G190gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT23), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n324_), .A2(new_n326_), .A3(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT86), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n330_), .B1(new_n327_), .B2(KEYINPUT23), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n331_), .B1(new_n328_), .B2(new_n330_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT87), .ZN(new_n333_));
  NOR2_X1   g132(.A1(G183gat), .A2(G190gat), .ZN(new_n334_));
  OR3_X1    g133(.A1(new_n332_), .A2(new_n333_), .A3(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT22), .B(G169gat), .ZN(new_n336_));
  INV_X1    g135(.A(G176gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n333_), .B1(new_n332_), .B2(new_n334_), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n335_), .A2(new_n319_), .A3(new_n338_), .A4(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n329_), .A2(new_n340_), .ZN(new_n341_));
  XOR2_X1   g140(.A(KEYINPUT88), .B(KEYINPUT31), .Z(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT30), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n341_), .B(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G15gat), .B(G43gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G227gat), .A2(G233gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n344_), .B(new_n347_), .ZN(new_n348_));
  XOR2_X1   g147(.A(G113gat), .B(G120gat), .Z(new_n349_));
  XNOR2_X1  g148(.A(G127gat), .B(G134gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  XOR2_X1   g150(.A(G71gat), .B(G99gat), .Z(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n348_), .B(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  XOR2_X1   g154(.A(G211gat), .B(G218gat), .Z(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(G197gat), .ZN(new_n358_));
  AND2_X1   g157(.A1(new_n358_), .A2(G204gat), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n358_), .A2(G204gat), .ZN(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT21), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  OR3_X1    g160(.A1(new_n358_), .A2(KEYINPUT90), .A3(G204gat), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n359_), .A2(KEYINPUT90), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n362_), .B1(new_n363_), .B2(new_n360_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n357_), .B(new_n361_), .C1(new_n364_), .C2(KEYINPUT21), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n364_), .A2(KEYINPUT21), .A3(new_n356_), .ZN(new_n366_));
  AND2_X1   g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  OR4_X1    g166(.A1(KEYINPUT89), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT2), .ZN(new_n369_));
  INV_X1    g168(.A(G141gat), .ZN(new_n370_));
  INV_X1    g169(.A(G148gat), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n369_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n373_));
  OAI22_X1  g172(.A1(KEYINPUT89), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n368_), .A2(new_n372_), .A3(new_n373_), .A4(new_n374_), .ZN(new_n375_));
  AND2_X1   g174(.A1(G155gat), .A2(G162gat), .ZN(new_n376_));
  NOR2_X1   g175(.A1(G155gat), .A2(G162gat), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n375_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT1), .ZN(new_n380_));
  AOI22_X1  g179(.A1(new_n378_), .A2(new_n380_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n381_));
  AOI22_X1  g180(.A1(new_n376_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n379_), .A2(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n367_), .B1(KEYINPUT29), .B2(new_n384_), .ZN(new_n385_));
  AND2_X1   g184(.A1(G228gat), .A2(G233gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT92), .ZN(new_n388_));
  XOR2_X1   g187(.A(G78gat), .B(G106gat), .Z(new_n389_));
  NOR2_X1   g188(.A1(new_n389_), .A2(KEYINPUT91), .ZN(new_n390_));
  XOR2_X1   g189(.A(new_n388_), .B(new_n390_), .Z(new_n391_));
  AOI21_X1  g190(.A(KEYINPUT92), .B1(new_n387_), .B2(new_n389_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n384_), .A2(KEYINPUT29), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT28), .B(G22gat), .ZN(new_n394_));
  INV_X1    g193(.A(G50gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n393_), .B(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n392_), .A2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n387_), .B(new_n389_), .ZN(new_n400_));
  AOI22_X1  g199(.A1(new_n391_), .A2(new_n399_), .B1(new_n400_), .B2(new_n398_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G1gat), .B(G29gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(G85gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(KEYINPUT0), .B(G57gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n384_), .B(new_n351_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G225gat), .A2(G233gat), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n406_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(KEYINPUT101), .ZN(new_n410_));
  INV_X1    g209(.A(new_n407_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT4), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT4), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n384_), .A2(new_n413_), .A3(new_n351_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n412_), .A2(new_n408_), .A3(new_n414_), .ZN(new_n415_));
  OR2_X1    g214(.A1(new_n415_), .A2(KEYINPUT102), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(KEYINPUT102), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n410_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT33), .ZN(new_n419_));
  INV_X1    g218(.A(new_n408_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n412_), .A2(new_n420_), .A3(new_n414_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT99), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n411_), .A2(new_n408_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n412_), .A2(KEYINPUT99), .A3(new_n420_), .A4(new_n414_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n406_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n423_), .A2(new_n424_), .A3(new_n425_), .A4(new_n426_), .ZN(new_n427_));
  OAI22_X1  g226(.A1(new_n418_), .A2(KEYINPUT103), .B1(new_n419_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT100), .ZN(new_n429_));
  AND3_X1   g228(.A1(new_n427_), .A2(new_n429_), .A3(new_n419_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n429_), .B1(new_n427_), .B2(new_n419_), .ZN(new_n431_));
  NOR3_X1   g230(.A1(new_n428_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT98), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G226gat), .A2(G233gat), .ZN(new_n434_));
  XOR2_X1   g233(.A(new_n434_), .B(KEYINPUT19), .Z(new_n435_));
  NAND2_X1  g234(.A1(new_n338_), .A2(new_n319_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n334_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n436_), .B1(new_n328_), .B2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n321_), .ZN(new_n439_));
  AOI22_X1  g238(.A1(new_n316_), .A2(new_n315_), .B1(new_n439_), .B2(new_n318_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT94), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n332_), .A2(new_n325_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n438_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(new_n367_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(KEYINPUT20), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT95), .ZN(new_n447_));
  INV_X1    g246(.A(new_n367_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n447_), .B1(new_n341_), .B2(new_n448_), .ZN(new_n449_));
  AOI211_X1 g248(.A(KEYINPUT95), .B(new_n367_), .C1(new_n329_), .C2(new_n340_), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n435_), .B(new_n446_), .C1(new_n449_), .C2(new_n450_), .ZN(new_n451_));
  OR2_X1    g250(.A1(new_n443_), .A2(new_n367_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n329_), .A2(new_n340_), .A3(new_n367_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n452_), .A2(new_n453_), .A3(KEYINPUT20), .ZN(new_n454_));
  XOR2_X1   g253(.A(new_n435_), .B(KEYINPUT93), .Z(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n454_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n451_), .A2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G64gat), .B(G92gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G8gat), .B(G36gat), .ZN(new_n462_));
  XOR2_X1   g261(.A(new_n461_), .B(new_n462_), .Z(new_n463_));
  AOI21_X1  g262(.A(new_n433_), .B1(new_n458_), .B2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n458_), .A2(new_n433_), .A3(new_n463_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n463_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n451_), .A2(new_n457_), .A3(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT97), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n451_), .A2(KEYINPUT97), .A3(new_n457_), .A4(new_n467_), .ZN(new_n471_));
  AOI22_X1  g270(.A1(new_n465_), .A2(new_n466_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n418_), .A2(KEYINPUT103), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n432_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(KEYINPUT104), .B1(new_n454_), .B2(new_n456_), .ZN(new_n475_));
  OR3_X1    g274(.A1(new_n454_), .A2(KEYINPUT104), .A3(new_n456_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n449_), .A2(new_n450_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n477_), .A2(new_n445_), .ZN(new_n478_));
  OAI211_X1 g277(.A(new_n475_), .B(new_n476_), .C1(new_n478_), .C2(new_n435_), .ZN(new_n479_));
  AND2_X1   g278(.A1(new_n467_), .A2(KEYINPUT32), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n423_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(new_n406_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(new_n427_), .ZN(new_n484_));
  OAI211_X1 g283(.A(new_n481_), .B(new_n484_), .C1(new_n458_), .C2(new_n480_), .ZN(new_n485_));
  AOI211_X1 g284(.A(new_n355_), .B(new_n402_), .C1(new_n474_), .C2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n479_), .A2(new_n463_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n487_), .A2(KEYINPUT27), .A3(new_n468_), .ZN(new_n488_));
  OAI211_X1 g287(.A(new_n401_), .B(new_n488_), .C1(new_n472_), .C2(KEYINPUT27), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(KEYINPUT105), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n470_), .A2(new_n471_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n466_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n491_), .B1(new_n492_), .B2(new_n464_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT27), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT105), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n495_), .A2(new_n496_), .A3(new_n401_), .A4(new_n488_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n490_), .A2(new_n355_), .A3(new_n497_), .ZN(new_n498_));
  AND2_X1   g297(.A1(new_n495_), .A2(new_n488_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n499_), .A2(new_n354_), .A3(new_n402_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n498_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n484_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n486_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G43gat), .B(G50gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(G36gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(KEYINPUT76), .B(G29gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT15), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G15gat), .B(G22gat), .ZN(new_n510_));
  INV_X1    g309(.A(G1gat), .ZN(new_n511_));
  INV_X1    g310(.A(G8gat), .ZN(new_n512_));
  OAI21_X1  g311(.A(KEYINPUT14), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n510_), .A2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G1gat), .B(G8gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n509_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT81), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G229gat), .A2(G233gat), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n507_), .A2(new_n516_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n509_), .A2(KEYINPUT81), .A3(new_n516_), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n519_), .A2(new_n520_), .A3(new_n521_), .A4(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n507_), .B(new_n516_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n524_), .A2(G229gat), .A3(G233gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G113gat), .B(G141gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G169gat), .B(G197gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT82), .B1(new_n526_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT82), .ZN(new_n531_));
  INV_X1    g330(.A(new_n529_), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n523_), .A2(new_n531_), .A3(new_n525_), .A4(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n530_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n526_), .A2(new_n529_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(KEYINPUT106), .B1(new_n503_), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT106), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n484_), .B1(new_n498_), .B2(new_n500_), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n539_), .B(new_n536_), .C1(new_n540_), .C2(new_n486_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n311_), .B1(new_n538_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT35), .ZN(new_n543_));
  INV_X1    g342(.A(new_n507_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n289_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT77), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n543_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT75), .B(KEYINPUT34), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G232gat), .A2(G233gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n547_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n271_), .A2(new_n272_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(new_n286_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n509_), .A2(new_n553_), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n550_), .A2(KEYINPUT35), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n551_), .A2(new_n545_), .A3(new_n554_), .A4(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n554_), .A2(new_n545_), .A3(new_n555_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n557_), .A2(new_n550_), .A3(new_n547_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G190gat), .B(G218gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G134gat), .B(G162gat), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n559_), .B(new_n560_), .Z(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n562_), .A2(KEYINPUT36), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n556_), .A2(new_n558_), .A3(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT78), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n556_), .A2(new_n558_), .A3(KEYINPUT78), .A4(new_n563_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n556_), .A2(new_n558_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n561_), .B(KEYINPUT36), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n568_), .A2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(KEYINPUT79), .B(KEYINPUT37), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n568_), .A2(new_n571_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n573_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n574_), .A2(new_n577_), .ZN(new_n578_));
  AND2_X1   g377(.A1(G231gat), .A2(G233gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n516_), .B(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n290_), .B(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G183gat), .B(G211gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  XOR2_X1   g384(.A(G127gat), .B(G155gat), .Z(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT17), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n283_), .A2(new_n284_), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n589_), .B(new_n580_), .Z(new_n590_));
  INV_X1    g389(.A(KEYINPUT17), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n587_), .A2(new_n591_), .ZN(new_n592_));
  AOI22_X1  g391(.A1(new_n582_), .A2(new_n588_), .B1(new_n590_), .B2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n578_), .A2(new_n594_), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n542_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n596_), .A2(new_n511_), .A3(new_n484_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT38), .ZN(new_n598_));
  OR2_X1    g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n501_), .A2(new_n502_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n486_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n311_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT107), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n603_), .A2(new_n604_), .A3(new_n536_), .ZN(new_n605_));
  OAI21_X1  g404(.A(KEYINPUT107), .B1(new_n311_), .B2(new_n537_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n605_), .A2(new_n606_), .A3(new_n593_), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n602_), .A2(KEYINPUT108), .A3(new_n575_), .A4(new_n607_), .ZN(new_n608_));
  OAI211_X1 g407(.A(new_n607_), .B(new_n575_), .C1(new_n540_), .C2(new_n486_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT108), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n608_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(G1gat), .B1(new_n613_), .B2(new_n502_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n597_), .A2(new_n598_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n599_), .A2(new_n614_), .A3(new_n615_), .ZN(G1324gat));
  INV_X1    g415(.A(new_n499_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n596_), .A2(new_n512_), .A3(new_n617_), .ZN(new_n618_));
  OAI21_X1  g417(.A(G8gat), .B1(new_n609_), .B2(new_n499_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT39), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT40), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n618_), .A2(KEYINPUT40), .A3(new_n620_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(G1325gat));
  INV_X1    g424(.A(G15gat), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n626_), .B1(new_n612_), .B2(new_n355_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT41), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n596_), .A2(new_n626_), .A3(new_n355_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(G1326gat));
  INV_X1    g429(.A(G22gat), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n542_), .A2(new_n631_), .A3(new_n402_), .A4(new_n595_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT42), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n612_), .A2(new_n402_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n633_), .B1(new_n634_), .B2(G22gat), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n401_), .B1(new_n608_), .B2(new_n611_), .ZN(new_n636_));
  NOR3_X1   g435(.A1(new_n636_), .A2(KEYINPUT42), .A3(new_n631_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n632_), .B1(new_n635_), .B2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT109), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  OAI211_X1 g439(.A(KEYINPUT109), .B(new_n632_), .C1(new_n635_), .C2(new_n637_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(G1327gat));
  INV_X1    g441(.A(KEYINPUT44), .ZN(new_n643_));
  INV_X1    g442(.A(new_n578_), .ZN(new_n644_));
  OAI21_X1  g443(.A(KEYINPUT43), .B1(new_n503_), .B2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT43), .ZN(new_n646_));
  OAI211_X1 g445(.A(new_n646_), .B(new_n578_), .C1(new_n540_), .C2(new_n486_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n605_), .A2(new_n606_), .A3(new_n594_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n643_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n649_), .B1(new_n645_), .B2(new_n647_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(KEYINPUT44), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n650_), .A2(G29gat), .A3(new_n484_), .A4(new_n652_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n575_), .A2(new_n593_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n542_), .A2(new_n484_), .A3(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(G29gat), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n653_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(KEYINPUT110), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT110), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n653_), .A2(new_n660_), .A3(new_n657_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n659_), .A2(new_n661_), .ZN(G1328gat));
  NAND2_X1  g461(.A1(new_n652_), .A2(new_n617_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n651_), .A2(KEYINPUT44), .ZN(new_n664_));
  OAI21_X1  g463(.A(G36gat), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n538_), .A2(new_n541_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n499_), .A2(G36gat), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n666_), .A2(new_n603_), .A3(new_n654_), .A4(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT45), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n542_), .A2(KEYINPUT45), .A3(new_n654_), .A4(new_n667_), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n665_), .A2(KEYINPUT46), .A3(new_n670_), .A4(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT46), .ZN(new_n673_));
  INV_X1    g472(.A(G36gat), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n499_), .B1(new_n651_), .B2(KEYINPUT44), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n674_), .B1(new_n650_), .B2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n670_), .A2(new_n671_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n673_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n672_), .A2(new_n678_), .ZN(G1329gat));
  NAND3_X1  g478(.A1(new_n542_), .A2(new_n355_), .A3(new_n654_), .ZN(new_n680_));
  INV_X1    g479(.A(G43gat), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n652_), .A2(G43gat), .A3(new_n355_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n682_), .B1(new_n683_), .B2(new_n664_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(KEYINPUT47), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT47), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n686_), .B(new_n682_), .C1(new_n683_), .C2(new_n664_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n685_), .A2(new_n687_), .ZN(G1330gat));
  AOI211_X1 g487(.A(new_n395_), .B(new_n401_), .C1(new_n651_), .C2(KEYINPUT44), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n542_), .A2(new_n402_), .A3(new_n654_), .ZN(new_n690_));
  AOI22_X1  g489(.A1(new_n689_), .A2(new_n650_), .B1(new_n395_), .B2(new_n690_), .ZN(G1331gat));
  NAND2_X1  g490(.A1(new_n311_), .A2(new_n537_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n692_), .A2(new_n594_), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n575_), .B(new_n693_), .C1(new_n540_), .C2(new_n486_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT112), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n694_), .B(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n696_), .A2(G57gat), .A3(new_n484_), .ZN(new_n697_));
  XOR2_X1   g496(.A(new_n697_), .B(KEYINPUT113), .Z(new_n698_));
  NAND2_X1  g497(.A1(new_n595_), .A2(new_n311_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT111), .Z(new_n700_));
  NOR2_X1   g499(.A1(new_n503_), .A2(new_n536_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(G57gat), .B1(new_n703_), .B2(new_n484_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n698_), .A2(new_n704_), .ZN(G1332gat));
  INV_X1    g504(.A(G64gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n706_), .B1(new_n696_), .B2(new_n617_), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT48), .Z(new_n708_));
  NAND3_X1  g507(.A1(new_n703_), .A2(new_n706_), .A3(new_n617_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1333gat));
  AOI21_X1  g509(.A(new_n237_), .B1(new_n696_), .B2(new_n355_), .ZN(new_n711_));
  XOR2_X1   g510(.A(new_n711_), .B(KEYINPUT49), .Z(new_n712_));
  NAND3_X1  g511(.A1(new_n703_), .A2(new_n237_), .A3(new_n355_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1334gat));
  NAND3_X1  g513(.A1(new_n703_), .A2(new_n238_), .A3(new_n402_), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n602_), .A2(new_n695_), .A3(new_n575_), .A4(new_n693_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n694_), .A2(KEYINPUT112), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n716_), .A2(new_n402_), .A3(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT50), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n718_), .A2(new_n719_), .A3(G78gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(new_n718_), .B2(G78gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n715_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT114), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  OAI211_X1 g523(.A(KEYINPUT114), .B(new_n715_), .C1(new_n720_), .C2(new_n721_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(G1335gat));
  AND2_X1   g525(.A1(new_n654_), .A2(new_n311_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n701_), .A2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(G85gat), .B1(new_n729_), .B2(new_n484_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n311_), .A2(new_n537_), .A3(new_n594_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n731_), .B1(new_n645_), .B2(new_n647_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n502_), .A2(new_n226_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n730_), .B1(new_n732_), .B2(new_n733_), .ZN(G1336gat));
  OAI21_X1  g533(.A(new_n227_), .B1(new_n728_), .B2(new_n499_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT115), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n617_), .A2(G92gat), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT116), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n736_), .B1(new_n732_), .B2(new_n738_), .ZN(G1337gat));
  NAND3_X1  g538(.A1(new_n729_), .A2(new_n233_), .A3(new_n355_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n732_), .A2(new_n355_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n740_), .B1(new_n741_), .B2(new_n204_), .ZN(new_n742_));
  AND2_X1   g541(.A1(KEYINPUT117), .A2(KEYINPUT51), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n742_), .B(new_n743_), .ZN(G1338gat));
  INV_X1    g543(.A(KEYINPUT52), .ZN(new_n745_));
  AOI211_X1 g544(.A(new_n401_), .B(new_n731_), .C1(new_n645_), .C2(new_n647_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n745_), .B1(new_n746_), .B2(new_n205_), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n701_), .A2(new_n205_), .A3(new_n402_), .A4(new_n727_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT118), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n732_), .A2(new_n402_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n750_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n747_), .A2(new_n749_), .A3(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT53), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT53), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n747_), .A2(new_n749_), .A3(new_n751_), .A4(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(G1339gat));
  NAND4_X1  g555(.A1(new_n574_), .A2(new_n577_), .A3(new_n537_), .A4(new_n593_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n757_), .A2(new_n311_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(KEYINPUT119), .B(KEYINPUT54), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n758_), .B(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n532_), .B1(new_n524_), .B2(new_n520_), .ZN(new_n762_));
  XOR2_X1   g561(.A(new_n762_), .B(KEYINPUT122), .Z(new_n763_));
  NAND3_X1  g562(.A1(new_n519_), .A2(new_n521_), .A3(new_n522_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n763_), .B1(new_n764_), .B2(new_n520_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n307_), .A2(new_n534_), .A3(new_n765_), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n263_), .A2(new_n267_), .A3(new_n264_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n267_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(KEYINPUT72), .B1(new_n553_), .B2(new_n285_), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n276_), .A2(new_n270_), .A3(new_n281_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n294_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n296_), .B1(new_n769_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT120), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT55), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n293_), .A2(new_n776_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n269_), .A2(new_n291_), .A3(KEYINPUT55), .A4(new_n292_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n282_), .A2(new_n288_), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n779_), .B(new_n294_), .C1(new_n767_), .C2(new_n768_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n780_), .A2(KEYINPUT120), .A3(new_n296_), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n775_), .A2(new_n777_), .A3(new_n778_), .A4(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(new_n303_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n783_), .A2(KEYINPUT121), .A3(KEYINPUT56), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(new_n536_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT121), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n786_), .B1(new_n782_), .B2(new_n303_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n306_), .B1(new_n787_), .B2(KEYINPUT56), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n766_), .B1(new_n785_), .B2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n789_), .A2(KEYINPUT57), .A3(new_n575_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT124), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n789_), .A2(new_n575_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT57), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n534_), .A2(new_n765_), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n777_), .A2(new_n778_), .ZN(new_n797_));
  AOI211_X1 g596(.A(new_n774_), .B(new_n292_), .C1(new_n269_), .C2(new_n291_), .ZN(new_n798_));
  AOI21_X1  g597(.A(KEYINPUT120), .B1(new_n780_), .B2(new_n296_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n305_), .B1(new_n797_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT56), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n796_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n306_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(new_n783_), .B2(KEYINPUT56), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT58), .ZN(new_n807_));
  AOI22_X1  g606(.A1(new_n806_), .A2(new_n807_), .B1(new_n574_), .B2(new_n577_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n803_), .A2(new_n805_), .A3(KEYINPUT58), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT123), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT123), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n803_), .A2(new_n805_), .A3(new_n811_), .A4(KEYINPUT58), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n808_), .A2(new_n810_), .A3(new_n812_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n789_), .A2(KEYINPUT124), .A3(KEYINPUT57), .A4(new_n575_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n792_), .A2(new_n795_), .A3(new_n813_), .A4(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n761_), .B1(new_n815_), .B2(new_n594_), .ZN(new_n816_));
  NOR3_X1   g615(.A1(new_n816_), .A2(new_n502_), .A3(new_n498_), .ZN(new_n817_));
  AOI21_X1  g616(.A(G113gat), .B1(new_n817_), .B2(new_n536_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT59), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n815_), .A2(new_n594_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n761_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n484_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n819_), .B1(new_n823_), .B2(new_n498_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n817_), .A2(KEYINPUT59), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n537_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n818_), .B1(new_n826_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g626(.A(KEYINPUT60), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n828_), .B1(new_n603_), .B2(G120gat), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n817_), .B(new_n829_), .C1(new_n828_), .C2(G120gat), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n603_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n831_));
  INV_X1    g630(.A(G120gat), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n830_), .B1(new_n831_), .B2(new_n832_), .ZN(G1341gat));
  AOI21_X1  g632(.A(G127gat), .B1(new_n817_), .B2(new_n593_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n594_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n834_), .B1(new_n835_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g635(.A(G134gat), .B1(new_n817_), .B2(new_n572_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n644_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n837_), .B1(new_n838_), .B2(G134gat), .ZN(G1343gat));
  NOR2_X1   g638(.A1(new_n823_), .A2(new_n500_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n536_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g641(.A1(new_n840_), .A2(new_n311_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n843_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g643(.A1(new_n840_), .A2(new_n593_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(KEYINPUT61), .B(G155gat), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n845_), .B(new_n846_), .ZN(G1346gat));
  AOI21_X1  g646(.A(G162gat), .B1(new_n840_), .B2(new_n572_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n578_), .A2(G162gat), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n848_), .B1(new_n840_), .B2(new_n849_), .ZN(G1347gat));
  NOR3_X1   g649(.A1(new_n402_), .A2(new_n484_), .A3(new_n354_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  NOR4_X1   g651(.A1(new_n816_), .A2(new_n499_), .A3(new_n537_), .A4(new_n852_), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n853_), .A2(new_n336_), .ZN(new_n854_));
  INV_X1    g653(.A(G169gat), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n853_), .A2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(KEYINPUT62), .B1(new_n854_), .B2(new_n856_), .ZN(new_n857_));
  OR2_X1    g656(.A1(new_n856_), .A2(KEYINPUT62), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(G1348gat));
  NAND2_X1  g658(.A1(new_n822_), .A2(new_n617_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n860_), .A2(new_n852_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(KEYINPUT125), .B(G176gat), .ZN(new_n862_));
  AND3_X1   g661(.A1(new_n861_), .A2(new_n311_), .A3(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n311_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(KEYINPUT125), .A2(G176gat), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n863_), .B1(new_n864_), .B2(new_n865_), .ZN(G1349gat));
  AOI21_X1  g665(.A(new_n499_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n867_), .A2(new_n593_), .A3(new_n851_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(G183gat), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT126), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n867_), .A2(new_n315_), .A3(new_n593_), .A4(new_n851_), .ZN(new_n871_));
  AND3_X1   g670(.A1(new_n869_), .A2(new_n870_), .A3(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n870_), .B1(new_n869_), .B2(new_n871_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n872_), .A2(new_n873_), .ZN(G1350gat));
  NAND3_X1  g673(.A1(new_n861_), .A2(new_n572_), .A3(new_n316_), .ZN(new_n875_));
  INV_X1    g674(.A(G190gat), .ZN(new_n876_));
  NOR3_X1   g675(.A1(new_n860_), .A2(new_n644_), .A3(new_n852_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n875_), .B1(new_n876_), .B2(new_n877_), .ZN(G1351gat));
  INV_X1    g677(.A(KEYINPUT127), .ZN(new_n879_));
  NOR3_X1   g678(.A1(new_n401_), .A2(new_n355_), .A3(new_n484_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n879_), .B1(new_n867_), .B2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n880_), .ZN(new_n882_));
  NOR4_X1   g681(.A1(new_n816_), .A2(KEYINPUT127), .A3(new_n499_), .A4(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n536_), .B1(new_n881_), .B2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(G197gat), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n802_), .B1(new_n801_), .B2(new_n786_), .ZN(new_n886_));
  NAND4_X1  g685(.A1(new_n886_), .A2(new_n536_), .A3(new_n306_), .A4(new_n784_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n572_), .B1(new_n887_), .B2(new_n766_), .ZN(new_n888_));
  AOI21_X1  g687(.A(KEYINPUT124), .B1(new_n888_), .B2(KEYINPUT57), .ZN(new_n889_));
  INV_X1    g688(.A(new_n814_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  AND2_X1   g690(.A1(new_n810_), .A2(new_n812_), .ZN(new_n892_));
  AOI22_X1  g691(.A1(new_n892_), .A2(new_n808_), .B1(new_n794_), .B2(new_n793_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n593_), .B1(new_n891_), .B2(new_n893_), .ZN(new_n894_));
  OAI211_X1 g693(.A(new_n617_), .B(new_n880_), .C1(new_n894_), .C2(new_n761_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(KEYINPUT127), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n867_), .A2(new_n879_), .A3(new_n880_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n898_), .A2(new_n358_), .A3(new_n536_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n885_), .A2(new_n899_), .ZN(G1352gat));
  AOI21_X1  g699(.A(G204gat), .B1(new_n898_), .B2(new_n311_), .ZN(new_n901_));
  OAI211_X1 g700(.A(G204gat), .B(new_n311_), .C1(new_n881_), .C2(new_n883_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n901_), .A2(new_n903_), .ZN(G1353gat));
  XOR2_X1   g703(.A(KEYINPUT63), .B(G211gat), .Z(new_n905_));
  OAI211_X1 g704(.A(new_n593_), .B(new_n905_), .C1(new_n881_), .C2(new_n883_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n594_), .B1(new_n896_), .B2(new_n897_), .ZN(new_n907_));
  OR2_X1    g706(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n906_), .B1(new_n907_), .B2(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n909_), .ZN(G1354gat));
  OAI211_X1 g709(.A(G218gat), .B(new_n578_), .C1(new_n881_), .C2(new_n883_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n575_), .B1(new_n896_), .B2(new_n897_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n911_), .B1(new_n912_), .B2(G218gat), .ZN(new_n913_));
  INV_X1    g712(.A(new_n913_), .ZN(G1355gat));
endmodule


