//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 0 0 1 1 0 1 0 0 0 1 1 1 1 1 0 0 1 0 0 1 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 0 0 1 0 1 1 0 0 1 0 0 1 0 1 1 0 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n691_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n838_, new_n839_, new_n841_, new_n842_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n849_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n881_, new_n882_,
    new_n883_, new_n885_, new_n886_, new_n887_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_;
  INV_X1    g000(.A(KEYINPUT37), .ZN(new_n202_));
  XOR2_X1   g001(.A(KEYINPUT10), .B(G99gat), .Z(new_n203_));
  INV_X1    g002(.A(G106gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G85gat), .ZN(new_n206_));
  INV_X1    g005(.A(G92gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G85gat), .A2(G92gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n208_), .A2(KEYINPUT9), .A3(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G99gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT6), .B1(new_n211_), .B2(new_n204_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT6), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n213_), .A2(G99gat), .A3(G106gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n209_), .A2(KEYINPUT9), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n205_), .A2(new_n210_), .A3(new_n215_), .A4(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT8), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT64), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT7), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n219_), .B(new_n220_), .C1(G99gat), .C2(G106gat), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n211_), .B(new_n204_), .C1(KEYINPUT64), .C2(KEYINPUT7), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT66), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT66), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n221_), .A2(new_n222_), .A3(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n224_), .A2(new_n226_), .A3(new_n215_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n208_), .A2(new_n209_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT65), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT65), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n208_), .A2(new_n230_), .A3(new_n209_), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n218_), .B1(new_n227_), .B2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n223_), .A2(new_n215_), .ZN(new_n234_));
  AND4_X1   g033(.A1(new_n218_), .A2(new_n234_), .A3(new_n229_), .A4(new_n231_), .ZN(new_n235_));
  OAI211_X1 g034(.A(KEYINPUT67), .B(new_n217_), .C1(new_n233_), .C2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n232_), .A2(new_n218_), .A3(new_n234_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n229_), .A2(new_n231_), .ZN(new_n239_));
  AOI22_X1  g038(.A1(new_n223_), .A2(KEYINPUT66), .B1(new_n212_), .B2(new_n214_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n239_), .B1(new_n240_), .B2(new_n226_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n238_), .B1(new_n241_), .B2(new_n218_), .ZN(new_n242_));
  AOI21_X1  g041(.A(KEYINPUT67), .B1(new_n242_), .B2(new_n217_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n237_), .A2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G29gat), .B(G36gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G43gat), .B(G50gat), .ZN(new_n246_));
  XOR2_X1   g045(.A(new_n245_), .B(new_n246_), .Z(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT71), .B(KEYINPUT72), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n244_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT15), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n247_), .A2(new_n248_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n247_), .A2(new_n248_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n251_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n245_), .B(new_n246_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(new_n248_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT15), .ZN(new_n257_));
  AND2_X1   g056(.A1(new_n254_), .A2(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n217_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n258_), .A2(KEYINPUT73), .A3(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT73), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n254_), .A2(new_n257_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n259_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n261_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n250_), .A2(new_n260_), .A3(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G232gat), .A2(G233gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT34), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT35), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  OR2_X1    g069(.A1(new_n270_), .A2(KEYINPUT75), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(KEYINPUT75), .ZN(new_n272_));
  OAI211_X1 g071(.A(new_n271_), .B(new_n272_), .C1(KEYINPUT35), .C2(new_n267_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n273_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n274_));
  AOI22_X1  g073(.A1(new_n265_), .A2(new_n270_), .B1(new_n250_), .B2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G190gat), .B(G218gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT74), .ZN(new_n277_));
  XOR2_X1   g076(.A(G134gat), .B(G162gat), .Z(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT36), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n275_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n279_), .A2(KEYINPUT36), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n275_), .A2(KEYINPUT76), .A3(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(KEYINPUT76), .B1(new_n275_), .B2(new_n283_), .ZN(new_n286_));
  OAI211_X1 g085(.A(new_n202_), .B(new_n282_), .C1(new_n285_), .C2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT76), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n265_), .A2(new_n270_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n274_), .A2(new_n250_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n283_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n288_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n280_), .B(KEYINPUT77), .ZN(new_n294_));
  AOI22_X1  g093(.A1(new_n293_), .A2(new_n284_), .B1(new_n291_), .B2(new_n294_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n287_), .B1(new_n295_), .B2(new_n202_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G57gat), .B(G64gat), .ZN(new_n297_));
  OR2_X1    g096(.A1(new_n297_), .A2(KEYINPUT11), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(KEYINPUT11), .ZN(new_n299_));
  XOR2_X1   g098(.A(G71gat), .B(G78gat), .Z(new_n300_));
  NAND3_X1  g099(.A1(new_n298_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n301_));
  OR2_X1    g100(.A1(new_n299_), .A2(new_n300_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G231gat), .A2(G233gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(KEYINPUT79), .ZN(new_n306_));
  INV_X1    g105(.A(G1gat), .ZN(new_n307_));
  INV_X1    g106(.A(G8gat), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT14), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT78), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT78), .ZN(new_n311_));
  OAI211_X1 g110(.A(new_n311_), .B(KEYINPUT14), .C1(new_n307_), .C2(new_n308_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G15gat), .B(G22gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n310_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G1gat), .B(G8gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n306_), .B(new_n317_), .ZN(new_n318_));
  XOR2_X1   g117(.A(G127gat), .B(G155gat), .Z(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT16), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G183gat), .B(G211gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT17), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  AND2_X1   g123(.A1(new_n322_), .A2(new_n323_), .ZN(new_n325_));
  OR3_X1    g124(.A1(new_n318_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n318_), .A2(new_n324_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n296_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n303_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n331_), .B1(new_n237_), .B2(new_n243_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT68), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT67), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n259_), .A2(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n335_), .A2(new_n303_), .A3(new_n236_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n332_), .A2(new_n333_), .A3(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G230gat), .A2(G233gat), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  OAI211_X1 g138(.A(new_n337_), .B(new_n339_), .C1(new_n333_), .C2(new_n332_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n259_), .A2(KEYINPUT12), .A3(new_n331_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n342_), .B1(new_n244_), .B2(new_n303_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT12), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n332_), .A2(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n343_), .A2(new_n345_), .A3(new_n338_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n340_), .A2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G120gat), .B(G148gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT5), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G176gat), .B(G204gat), .ZN(new_n350_));
  XOR2_X1   g149(.A(new_n349_), .B(new_n350_), .Z(new_n351_));
  OR2_X1    g150(.A1(new_n347_), .A2(new_n351_), .ZN(new_n352_));
  XOR2_X1   g151(.A(new_n351_), .B(KEYINPUT69), .Z(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n347_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT13), .ZN(new_n356_));
  OAI211_X1 g155(.A(new_n352_), .B(new_n355_), .C1(KEYINPUT70), .C2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n355_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n347_), .A2(new_n351_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT70), .B(KEYINPUT13), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n357_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n330_), .A2(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT80), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G8gat), .B(G36gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT18), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G64gat), .B(G92gat), .ZN(new_n368_));
  XOR2_X1   g167(.A(new_n367_), .B(new_n368_), .Z(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(G197gat), .ZN(new_n371_));
  OAI21_X1  g170(.A(KEYINPUT94), .B1(new_n371_), .B2(G204gat), .ZN(new_n372_));
  INV_X1    g171(.A(G204gat), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n372_), .B1(G197gat), .B2(new_n373_), .ZN(new_n374_));
  NOR3_X1   g173(.A1(new_n371_), .A2(KEYINPUT94), .A3(G204gat), .ZN(new_n375_));
  OAI21_X1  g174(.A(KEYINPUT21), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G211gat), .B(G218gat), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT95), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n378_), .B1(new_n371_), .B2(G204gat), .ZN(new_n379_));
  NOR3_X1   g178(.A1(new_n373_), .A2(KEYINPUT95), .A3(G197gat), .ZN(new_n380_));
  OAI22_X1  g179(.A1(new_n379_), .A2(new_n380_), .B1(new_n371_), .B2(G204gat), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n376_), .B(new_n377_), .C1(new_n381_), .C2(KEYINPUT21), .ZN(new_n382_));
  INV_X1    g181(.A(new_n377_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n381_), .A2(KEYINPUT21), .A3(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n382_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G183gat), .A2(G190gat), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT87), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT23), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n387_), .A2(KEYINPUT23), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n391_), .A2(KEYINPUT88), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n389_), .A2(KEYINPUT88), .A3(KEYINPUT23), .ZN(new_n394_));
  NOR2_X1   g193(.A1(G169gat), .A2(G176gat), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT85), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT24), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n393_), .A2(new_n394_), .A3(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(KEYINPUT96), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT96), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n393_), .A2(new_n402_), .A3(new_n394_), .A4(new_n399_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(G169gat), .ZN(new_n405_));
  INV_X1    g204(.A(G176gat), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT24), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  OR2_X1    g206(.A1(new_n397_), .A2(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(KEYINPUT25), .B(G183gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(KEYINPUT26), .B(G190gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n408_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n404_), .A2(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n389_), .A2(KEYINPUT23), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n387_), .A2(KEYINPUT23), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT86), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  OR2_X1    g217(.A1(new_n415_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT97), .ZN(new_n420_));
  OR2_X1    g219(.A1(G183gat), .A2(G190gat), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n419_), .A2(new_n420_), .A3(new_n421_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(G169gat), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n421_), .B1(new_n415_), .B2(new_n418_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(KEYINPUT97), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n422_), .A2(new_n424_), .A3(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n386_), .B1(new_n414_), .B2(new_n427_), .ZN(new_n428_));
  AND3_X1   g227(.A1(new_n408_), .A2(new_n411_), .A3(new_n399_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(new_n419_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n393_), .A2(new_n421_), .A3(new_n394_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(new_n424_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n430_), .A2(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT20), .B1(new_n433_), .B2(new_n385_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G226gat), .A2(G233gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(KEYINPUT19), .ZN(new_n436_));
  NOR3_X1   g235(.A1(new_n428_), .A2(new_n434_), .A3(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n436_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n414_), .A2(new_n386_), .A3(new_n427_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT20), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n440_), .B1(new_n433_), .B2(new_n385_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n438_), .B1(new_n439_), .B2(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n370_), .B1(new_n437_), .B2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(KEYINPUT27), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT98), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n445_), .B(new_n436_), .C1(new_n428_), .C2(new_n434_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n439_), .A2(new_n441_), .A3(new_n438_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  AND3_X1   g247(.A1(new_n422_), .A2(new_n424_), .A3(new_n426_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n412_), .B1(new_n401_), .B2(new_n403_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n385_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  AOI22_X1  g250(.A1(new_n429_), .A2(new_n419_), .B1(new_n424_), .B2(new_n431_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n440_), .B1(new_n452_), .B2(new_n386_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n438_), .B1(new_n451_), .B2(new_n453_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n454_), .A2(new_n445_), .ZN(new_n455_));
  NOR3_X1   g254(.A1(new_n448_), .A2(new_n455_), .A3(new_n370_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT106), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n444_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  OR2_X1    g257(.A1(new_n454_), .A2(new_n445_), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n459_), .A2(new_n369_), .A3(new_n447_), .A4(new_n446_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT106), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n370_), .B1(new_n448_), .B2(new_n455_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  XOR2_X1   g262(.A(KEYINPUT107), .B(KEYINPUT27), .Z(new_n464_));
  AOI22_X1  g263(.A1(new_n458_), .A2(new_n461_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G227gat), .A2(G233gat), .ZN(new_n466_));
  XOR2_X1   g265(.A(new_n466_), .B(G15gat), .Z(new_n467_));
  XNOR2_X1  g266(.A(new_n433_), .B(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(KEYINPUT31), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G71gat), .B(G99gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n470_), .B(G43gat), .ZN(new_n471_));
  XOR2_X1   g270(.A(KEYINPUT89), .B(KEYINPUT30), .Z(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  XOR2_X1   g272(.A(G127gat), .B(G134gat), .Z(new_n474_));
  XOR2_X1   g273(.A(G113gat), .B(G120gat), .Z(new_n475_));
  XOR2_X1   g274(.A(new_n474_), .B(new_n475_), .Z(new_n476_));
  XNOR2_X1  g275(.A(new_n473_), .B(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n469_), .B(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT3), .ZN(new_n479_));
  INV_X1    g278(.A(G141gat), .ZN(new_n480_));
  INV_X1    g279(.A(G148gat), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n479_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G141gat), .A2(G148gat), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT2), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n482_), .A2(new_n485_), .A3(new_n486_), .A4(new_n487_), .ZN(new_n488_));
  XOR2_X1   g287(.A(G155gat), .B(G162gat), .Z(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT91), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(G155gat), .A2(G162gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G155gat), .A2(G162gat), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n493_), .B1(KEYINPUT1), .B2(new_n494_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n495_), .B1(KEYINPUT1), .B2(new_n494_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n480_), .A2(new_n481_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n496_), .A2(new_n483_), .A3(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n492_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(new_n476_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT99), .ZN(new_n501_));
  INV_X1    g300(.A(new_n476_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n492_), .A2(new_n502_), .A3(new_n498_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n500_), .A2(new_n501_), .A3(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n499_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n505_), .A2(KEYINPUT99), .A3(new_n502_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G225gat), .A2(G233gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  XOR2_X1   g308(.A(new_n508_), .B(KEYINPUT100), .Z(new_n510_));
  INV_X1    g309(.A(KEYINPUT4), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n499_), .A2(new_n511_), .A3(new_n476_), .ZN(new_n512_));
  AND2_X1   g311(.A1(new_n512_), .A2(KEYINPUT101), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n512_), .A2(KEYINPUT101), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n510_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n511_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n509_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G1gat), .B(G29gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(KEYINPUT102), .B(KEYINPUT0), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G57gat), .B(G85gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n517_), .A2(new_n523_), .ZN(new_n524_));
  OAI211_X1 g323(.A(new_n522_), .B(new_n509_), .C1(new_n515_), .C2(new_n516_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT29), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n385_), .B1(new_n505_), .B2(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(KEYINPUT92), .B(KEYINPUT28), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n505_), .A2(new_n528_), .ZN(new_n532_));
  XOR2_X1   g331(.A(G22gat), .B(G50gat), .Z(new_n533_));
  OR2_X1    g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  AND2_X1   g333(.A1(KEYINPUT93), .A2(G228gat), .ZN(new_n535_));
  NOR2_X1   g334(.A1(KEYINPUT93), .A2(G228gat), .ZN(new_n536_));
  OAI21_X1  g335(.A(G233gat), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(G78gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(G106gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n532_), .A2(new_n533_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n534_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n540_), .B1(new_n534_), .B2(new_n541_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n531_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n544_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n531_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n546_), .A2(new_n547_), .A3(new_n542_), .ZN(new_n548_));
  AND2_X1   g347(.A1(new_n545_), .A2(new_n548_), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n465_), .A2(new_n478_), .A3(new_n527_), .A4(new_n549_), .ZN(new_n550_));
  OAI211_X1 g349(.A(KEYINPUT32), .B(new_n369_), .C1(new_n437_), .C2(new_n442_), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n551_), .A2(KEYINPUT105), .ZN(new_n552_));
  INV_X1    g351(.A(new_n448_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n369_), .A2(KEYINPUT32), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n553_), .A2(new_n459_), .A3(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n551_), .A2(KEYINPUT105), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n552_), .A2(new_n526_), .A3(new_n555_), .A4(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n522_), .B1(new_n507_), .B2(new_n510_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n508_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n558_), .B1(new_n516_), .B2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(KEYINPUT104), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT104), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n558_), .B(new_n562_), .C1(new_n516_), .C2(new_n559_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n525_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(KEYINPUT33), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n564_), .A2(new_n566_), .A3(new_n460_), .A4(new_n462_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT103), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT33), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n525_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n568_), .B1(new_n525_), .B2(new_n569_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n557_), .B1(new_n567_), .B2(new_n573_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n549_), .A2(new_n526_), .ZN(new_n575_));
  AOI22_X1  g374(.A1(new_n574_), .A2(new_n549_), .B1(new_n465_), .B2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n478_), .B(KEYINPUT90), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n550_), .B1(new_n576_), .B2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  XOR2_X1   g379(.A(G113gat), .B(G141gat), .Z(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT82), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G169gat), .B(G197gat), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n582_), .B(new_n583_), .Z(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT81), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n249_), .A2(new_n586_), .A3(new_n317_), .ZN(new_n587_));
  OAI21_X1  g386(.A(KEYINPUT81), .B1(new_n256_), .B2(new_n316_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n256_), .A2(new_n316_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G229gat), .A2(G233gat), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n254_), .A2(new_n257_), .A3(new_n316_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n589_), .A2(new_n592_), .A3(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n585_), .B1(new_n594_), .B2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n594_), .A2(new_n596_), .A3(new_n585_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(KEYINPUT83), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT83), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n594_), .A2(new_n596_), .A3(new_n600_), .A4(new_n585_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n597_), .B1(new_n599_), .B2(new_n601_), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n602_), .B(KEYINPUT84), .Z(new_n603_));
  NOR2_X1   g402(.A1(new_n580_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n365_), .A2(new_n604_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n526_), .A2(KEYINPUT108), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n526_), .A2(KEYINPUT108), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(new_n307_), .ZN(new_n609_));
  OR3_X1    g408(.A1(new_n605_), .A2(KEYINPUT109), .A3(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(KEYINPUT109), .B1(new_n605_), .B2(new_n609_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n610_), .A2(KEYINPUT38), .A3(new_n611_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n282_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n602_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n362_), .A2(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n615_), .A2(new_n328_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n579_), .A2(new_n613_), .A3(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT110), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n617_), .A2(new_n618_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n526_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(G1gat), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n612_), .A2(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(KEYINPUT38), .B1(new_n610_), .B2(new_n611_), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n623_), .A2(new_n624_), .ZN(G1324gat));
  NOR2_X1   g424(.A1(new_n465_), .A2(G8gat), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n365_), .A2(new_n604_), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT111), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n617_), .A2(new_n465_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n630_), .A2(KEYINPUT39), .A3(G8gat), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(G8gat), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT39), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n629_), .A2(new_n631_), .A3(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT40), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n629_), .A2(KEYINPUT40), .A3(new_n631_), .A4(new_n634_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(G1325gat));
  OR3_X1    g438(.A1(new_n605_), .A2(G15gat), .A3(new_n577_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n578_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n641_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n642_));
  AOI21_X1  g441(.A(KEYINPUT41), .B1(new_n641_), .B2(G15gat), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n640_), .B1(new_n642_), .B2(new_n643_), .ZN(G1326gat));
  OR3_X1    g443(.A1(new_n605_), .A2(G22gat), .A3(new_n549_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n549_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n646_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT42), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n647_), .A2(new_n648_), .A3(G22gat), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n648_), .B1(new_n647_), .B2(G22gat), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n645_), .B1(new_n649_), .B2(new_n650_), .ZN(G1327gat));
  NOR2_X1   g450(.A1(new_n615_), .A2(new_n329_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT43), .ZN(new_n653_));
  INV_X1    g452(.A(new_n296_), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n579_), .A2(new_n653_), .A3(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n653_), .B1(new_n579_), .B2(new_n654_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n652_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT44), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  OAI211_X1 g458(.A(KEYINPUT44), .B(new_n652_), .C1(new_n655_), .C2(new_n656_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n608_), .ZN(new_n662_));
  INV_X1    g461(.A(G29gat), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n613_), .A2(new_n329_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n362_), .A2(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n604_), .A2(new_n526_), .A3(new_n666_), .ZN(new_n667_));
  AOI22_X1  g466(.A1(new_n661_), .A2(new_n664_), .B1(new_n663_), .B2(new_n667_), .ZN(G1328gat));
  INV_X1    g467(.A(new_n465_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n659_), .A2(new_n669_), .A3(new_n660_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(G36gat), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n465_), .A2(KEYINPUT112), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n465_), .A2(KEYINPUT112), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n674_), .A2(G36gat), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n604_), .A2(new_n666_), .A3(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT45), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n671_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT46), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n671_), .A2(KEYINPUT46), .A3(new_n677_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(G1329gat));
  NAND4_X1  g481(.A1(new_n659_), .A2(G43gat), .A3(new_n478_), .A4(new_n660_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n603_), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n579_), .A2(new_n578_), .A3(new_n684_), .A4(new_n666_), .ZN(new_n685_));
  XOR2_X1   g484(.A(KEYINPUT113), .B(G43gat), .Z(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n687_), .B(KEYINPUT114), .Z(new_n688_));
  NAND2_X1  g487(.A1(new_n683_), .A2(new_n688_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g489(.A(G50gat), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n549_), .A2(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n604_), .A2(new_n646_), .A3(new_n666_), .ZN(new_n693_));
  AOI22_X1  g492(.A1(new_n661_), .A2(new_n692_), .B1(new_n691_), .B2(new_n693_), .ZN(G1331gat));
  OAI21_X1  g493(.A(KEYINPUT115), .B1(new_n580_), .B2(new_n614_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT115), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n579_), .A2(new_n696_), .A3(new_n602_), .ZN(new_n697_));
  AOI211_X1 g496(.A(new_n362_), .B(new_n330_), .C1(new_n695_), .C2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(G57gat), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n698_), .A2(new_n699_), .A3(new_n608_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n613_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n580_), .A2(new_n701_), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n684_), .A2(new_n362_), .A3(new_n328_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n702_), .A2(new_n526_), .A3(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(G57gat), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n700_), .A2(new_n705_), .ZN(G1332gat));
  INV_X1    g505(.A(G64gat), .ZN(new_n707_));
  INV_X1    g506(.A(new_n674_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n698_), .A2(new_n707_), .A3(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n702_), .A2(new_n708_), .A3(new_n703_), .ZN(new_n710_));
  XOR2_X1   g509(.A(KEYINPUT116), .B(KEYINPUT48), .Z(new_n711_));
  AND3_X1   g510(.A1(new_n710_), .A2(G64gat), .A3(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n711_), .B1(new_n710_), .B2(G64gat), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n709_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT117), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  OAI211_X1 g515(.A(new_n709_), .B(KEYINPUT117), .C1(new_n713_), .C2(new_n712_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(G1333gat));
  NAND3_X1  g517(.A1(new_n702_), .A2(new_n578_), .A3(new_n703_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(G71gat), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(KEYINPUT118), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT118), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n719_), .A2(new_n722_), .A3(G71gat), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n721_), .A2(KEYINPUT49), .A3(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(G71gat), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n698_), .A2(new_n725_), .A3(new_n578_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(KEYINPUT49), .B1(new_n721_), .B2(new_n723_), .ZN(new_n728_));
  OR2_X1    g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1334gat));
  NAND3_X1  g528(.A1(new_n702_), .A2(new_n646_), .A3(new_n703_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(G78gat), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(KEYINPUT119), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT119), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n730_), .A2(new_n733_), .A3(G78gat), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n732_), .A2(KEYINPUT50), .A3(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n698_), .A2(new_n538_), .A3(new_n646_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(KEYINPUT50), .B1(new_n732_), .B2(new_n734_), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n737_), .A2(new_n738_), .ZN(G1335gat));
  NAND2_X1  g538(.A1(new_n363_), .A2(new_n665_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(new_n695_), .B2(new_n697_), .ZN(new_n741_));
  AOI21_X1  g540(.A(G85gat), .B1(new_n741_), .B2(new_n608_), .ZN(new_n742_));
  NOR3_X1   g541(.A1(new_n362_), .A2(new_n329_), .A3(new_n614_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n743_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT120), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n527_), .A2(new_n206_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n742_), .B1(new_n745_), .B2(new_n746_), .ZN(G1336gat));
  AOI21_X1  g546(.A(G92gat), .B1(new_n741_), .B2(new_n669_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n674_), .A2(new_n207_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n745_), .B2(new_n749_), .ZN(G1337gat));
  AND2_X1   g549(.A1(new_n478_), .A2(new_n203_), .ZN(new_n751_));
  AOI22_X1  g550(.A1(new_n741_), .A2(new_n751_), .B1(KEYINPUT121), .B2(KEYINPUT51), .ZN(new_n752_));
  OAI21_X1  g551(.A(G99gat), .B1(new_n744_), .B2(new_n577_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(KEYINPUT121), .A2(KEYINPUT51), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT122), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n754_), .B(new_n756_), .ZN(G1338gat));
  NAND3_X1  g556(.A1(new_n741_), .A2(new_n204_), .A3(new_n646_), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n646_), .B(new_n743_), .C1(new_n655_), .C2(new_n656_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT52), .ZN(new_n760_));
  AND3_X1   g559(.A1(new_n759_), .A2(new_n760_), .A3(G106gat), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n760_), .B1(new_n759_), .B2(G106gat), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n758_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g563(.A1(new_n296_), .A2(new_n362_), .A3(new_n603_), .A4(new_n329_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT54), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n765_), .B(new_n766_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n602_), .A2(new_n359_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n338_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT55), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n346_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n343_), .A2(new_n345_), .A3(KEYINPUT55), .A4(new_n338_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(KEYINPUT56), .B1(new_n773_), .B2(new_n354_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT56), .ZN(new_n775_));
  AOI211_X1 g574(.A(new_n775_), .B(new_n353_), .C1(new_n771_), .C2(new_n772_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n768_), .B1(new_n774_), .B2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n599_), .A2(new_n601_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n591_), .A2(new_n592_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n589_), .A2(new_n593_), .A3(new_n595_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n779_), .A2(new_n780_), .A3(new_n584_), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n778_), .B(new_n781_), .C1(new_n358_), .C2(new_n359_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n701_), .B1(new_n777_), .B2(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(KEYINPUT57), .B1(new_n783_), .B2(KEYINPUT123), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT123), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT57), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n778_), .A2(new_n781_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n787_), .B1(new_n355_), .B2(new_n352_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n303_), .B1(new_n335_), .B2(new_n236_), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n336_), .B(new_n341_), .C1(new_n789_), .C2(KEYINPUT12), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n770_), .B1(new_n790_), .B2(new_n339_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n790_), .A2(new_n339_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n772_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n354_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n775_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n773_), .A2(KEYINPUT56), .A3(new_n354_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n788_), .B1(new_n798_), .B2(new_n768_), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n785_), .B(new_n786_), .C1(new_n799_), .C2(new_n701_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n787_), .A2(new_n359_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n801_), .B1(new_n774_), .B2(new_n776_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT58), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n798_), .A2(KEYINPUT58), .A3(new_n801_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n654_), .A2(new_n804_), .A3(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n784_), .A2(new_n800_), .A3(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n767_), .B1(new_n328_), .B2(new_n807_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n465_), .A2(new_n608_), .A3(new_n478_), .A4(new_n549_), .ZN(new_n809_));
  OAI21_X1  g608(.A(KEYINPUT59), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  XNOR2_X1  g609(.A(KEYINPUT125), .B(G113gat), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n603_), .A2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n807_), .A2(new_n328_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT124), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n807_), .A2(KEYINPUT124), .A3(new_n328_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n767_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  OR2_X1    g616(.A1(new_n809_), .A2(KEYINPUT59), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n810_), .B(new_n812_), .C1(new_n817_), .C2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(G113gat), .ZN(new_n820_));
  INV_X1    g619(.A(new_n767_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n813_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n809_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n820_), .B1(new_n824_), .B2(new_n602_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n819_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(KEYINPUT126), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT126), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n819_), .A2(new_n828_), .A3(new_n825_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n827_), .A2(new_n829_), .ZN(G1340gat));
  NOR2_X1   g629(.A1(new_n362_), .A2(KEYINPUT60), .ZN(new_n831_));
  MUX2_X1   g630(.A(new_n831_), .B(KEYINPUT60), .S(G120gat), .Z(new_n832_));
  NAND3_X1  g631(.A1(new_n822_), .A2(new_n823_), .A3(new_n832_), .ZN(new_n833_));
  XOR2_X1   g632(.A(new_n833_), .B(KEYINPUT127), .Z(new_n834_));
  OAI21_X1  g633(.A(new_n810_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n835_));
  OAI21_X1  g634(.A(G120gat), .B1(new_n835_), .B2(new_n362_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n836_), .ZN(G1341gat));
  OAI21_X1  g636(.A(G127gat), .B1(new_n835_), .B2(new_n328_), .ZN(new_n838_));
  OR2_X1    g637(.A1(new_n328_), .A2(G127gat), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n838_), .B1(new_n824_), .B2(new_n839_), .ZN(G1342gat));
  OAI21_X1  g639(.A(G134gat), .B1(new_n835_), .B2(new_n296_), .ZN(new_n841_));
  OR2_X1    g640(.A1(new_n613_), .A2(G134gat), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(new_n824_), .B2(new_n842_), .ZN(G1343gat));
  NOR2_X1   g642(.A1(new_n808_), .A2(new_n578_), .ZN(new_n844_));
  NOR3_X1   g643(.A1(new_n708_), .A2(new_n549_), .A3(new_n662_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n846_), .A2(new_n602_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n847_), .B(new_n480_), .ZN(G1344gat));
  NOR2_X1   g647(.A1(new_n846_), .A2(new_n362_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(new_n481_), .ZN(G1345gat));
  NOR2_X1   g649(.A1(new_n846_), .A2(new_n328_), .ZN(new_n851_));
  XOR2_X1   g650(.A(KEYINPUT61), .B(G155gat), .Z(new_n852_));
  XNOR2_X1  g651(.A(new_n851_), .B(new_n852_), .ZN(G1346gat));
  OAI21_X1  g652(.A(G162gat), .B1(new_n846_), .B2(new_n296_), .ZN(new_n854_));
  OR2_X1    g653(.A1(new_n613_), .A2(G162gat), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n846_), .B2(new_n855_), .ZN(G1347gat));
  AND3_X1   g655(.A1(new_n807_), .A2(KEYINPUT124), .A3(new_n328_), .ZN(new_n857_));
  AOI21_X1  g656(.A(KEYINPUT124), .B1(new_n807_), .B2(new_n328_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n821_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT22), .ZN(new_n860_));
  NOR3_X1   g659(.A1(new_n674_), .A2(new_n577_), .A3(new_n608_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n549_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n859_), .A2(new_n860_), .A3(new_n614_), .A4(new_n863_), .ZN(new_n864_));
  AND3_X1   g663(.A1(new_n864_), .A2(KEYINPUT62), .A3(new_n405_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(KEYINPUT62), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n817_), .A2(new_n602_), .A3(new_n862_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT62), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n405_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n865_), .B1(new_n866_), .B2(new_n869_), .ZN(G1348gat));
  NOR2_X1   g669(.A1(new_n817_), .A2(new_n862_), .ZN(new_n871_));
  AOI21_X1  g670(.A(G176gat), .B1(new_n871_), .B2(new_n363_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n808_), .A2(new_n646_), .ZN(new_n873_));
  AND3_X1   g672(.A1(new_n861_), .A2(G176gat), .A3(new_n363_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n872_), .B1(new_n873_), .B2(new_n874_), .ZN(G1349gat));
  NAND2_X1  g674(.A1(new_n861_), .A2(new_n329_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(G183gat), .B1(new_n873_), .B2(new_n877_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n328_), .A2(new_n409_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n878_), .B1(new_n871_), .B2(new_n879_), .ZN(G1350gat));
  NAND3_X1  g679(.A1(new_n871_), .A2(new_n410_), .A3(new_n701_), .ZN(new_n881_));
  INV_X1    g680(.A(G190gat), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n817_), .A2(new_n296_), .A3(new_n862_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n881_), .B1(new_n882_), .B2(new_n883_), .ZN(G1351gat));
  NOR3_X1   g683(.A1(new_n674_), .A2(new_n526_), .A3(new_n549_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n844_), .A2(new_n885_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n886_), .A2(new_n602_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(new_n371_), .ZN(G1352gat));
  NOR2_X1   g687(.A1(new_n886_), .A2(new_n362_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(new_n373_), .ZN(G1353gat));
  NAND3_X1  g689(.A1(new_n844_), .A2(new_n329_), .A3(new_n885_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n892_));
  AND2_X1   g691(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n893_));
  NOR3_X1   g692(.A1(new_n891_), .A2(new_n892_), .A3(new_n893_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n894_), .B1(new_n891_), .B2(new_n892_), .ZN(G1354gat));
  OAI21_X1  g694(.A(G218gat), .B1(new_n886_), .B2(new_n296_), .ZN(new_n896_));
  OR2_X1    g695(.A1(new_n613_), .A2(G218gat), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n886_), .B2(new_n897_), .ZN(G1355gat));
endmodule


