//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 0 1 0 1 1 1 1 1 1 0 0 0 1 0 1 0 1 0 1 0 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 1 0 0 0 1 0 0 1 0 1 0 1 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n836_,
    new_n837_, new_n838_, new_n840_, new_n841_, new_n842_, new_n844_,
    new_n845_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n853_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_, new_n884_, new_n885_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT69), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G29gat), .B(G36gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(KEYINPUT70), .B(KEYINPUT15), .Z(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  XOR2_X1   g006(.A(KEYINPUT10), .B(G99gat), .Z(new_n208_));
  INV_X1    g007(.A(G106gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  XOR2_X1   g009(.A(G85gat), .B(G92gat), .Z(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT9), .ZN(new_n212_));
  INV_X1    g011(.A(G85gat), .ZN(new_n213_));
  INV_X1    g012(.A(G92gat), .ZN(new_n214_));
  OR3_X1    g013(.A1(new_n213_), .A2(new_n214_), .A3(KEYINPUT9), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G99gat), .A2(G106gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT6), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n210_), .A2(new_n212_), .A3(new_n215_), .A4(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n219_));
  OR3_X1    g018(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n217_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(KEYINPUT64), .A2(KEYINPUT8), .ZN(new_n222_));
  AND3_X1   g021(.A1(new_n221_), .A2(new_n211_), .A3(new_n222_), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n222_), .B1(new_n221_), .B2(new_n211_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n218_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G232gat), .A2(G233gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT34), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  XOR2_X1   g027(.A(KEYINPUT68), .B(KEYINPUT35), .Z(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  AOI22_X1  g029(.A1(new_n207_), .A2(new_n225_), .B1(new_n228_), .B2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n225_), .A2(KEYINPUT65), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT65), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n233_), .B(new_n218_), .C1(new_n223_), .C2(new_n224_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n232_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(new_n205_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n231_), .A2(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n228_), .A2(new_n230_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n237_), .B(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G134gat), .B(G162gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT71), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G190gat), .B(G218gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n244_), .A2(KEYINPUT36), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n240_), .A2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n237_), .B(new_n238_), .ZN(new_n247_));
  XOR2_X1   g046(.A(new_n244_), .B(KEYINPUT36), .Z(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n246_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT37), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT37), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n246_), .A2(new_n249_), .A3(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G127gat), .B(G155gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(G211gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT16), .B(G183gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT17), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G15gat), .B(G22gat), .ZN(new_n261_));
  INV_X1    g060(.A(G1gat), .ZN(new_n262_));
  INV_X1    g061(.A(G8gat), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT14), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n261_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G1gat), .B(G8gat), .ZN(new_n266_));
  XOR2_X1   g065(.A(new_n265_), .B(new_n266_), .Z(new_n267_));
  NAND2_X1  g066(.A1(G231gat), .A2(G233gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  XOR2_X1   g068(.A(G57gat), .B(G64gat), .Z(new_n270_));
  INV_X1    g069(.A(KEYINPUT11), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT66), .ZN(new_n273_));
  XOR2_X1   g072(.A(G71gat), .B(G78gat), .Z(new_n274_));
  NAND3_X1  g073(.A1(new_n272_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n273_), .B1(new_n272_), .B2(new_n274_), .ZN(new_n277_));
  OAI22_X1  g076(.A1(new_n276_), .A2(new_n277_), .B1(new_n271_), .B2(new_n270_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n277_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n270_), .A2(new_n271_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n279_), .A2(new_n275_), .A3(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n278_), .A2(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n269_), .B(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT73), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n260_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n285_), .B1(new_n284_), .B2(new_n283_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n259_), .A2(KEYINPUT17), .ZN(new_n287_));
  XOR2_X1   g086(.A(new_n287_), .B(KEYINPUT72), .Z(new_n288_));
  OR2_X1    g087(.A1(new_n283_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n286_), .A2(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n255_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT74), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT96), .ZN(new_n293_));
  XOR2_X1   g092(.A(G64gat), .B(G92gat), .Z(new_n294_));
  XNOR2_X1  g093(.A(G8gat), .B(G36gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  AND3_X1   g097(.A1(KEYINPUT19), .A2(G226gat), .A3(G233gat), .ZN(new_n299_));
  AOI21_X1  g098(.A(KEYINPUT19), .B1(G226gat), .B2(G233gat), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  XOR2_X1   g100(.A(new_n301_), .B(KEYINPUT88), .Z(new_n302_));
  NAND2_X1  g101(.A1(G183gat), .A2(G190gat), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT23), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n306_));
  OAI211_X1 g105(.A(new_n305_), .B(new_n306_), .C1(G183gat), .C2(G190gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G169gat), .A2(G176gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(G169gat), .ZN(new_n310_));
  OR2_X1    g109(.A1(new_n310_), .A2(KEYINPUT22), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(KEYINPUT22), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n313_), .A2(G176gat), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n309_), .A2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT26), .B(G190gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT25), .B(G183gat), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT24), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n318_), .B1(G169gat), .B2(G176gat), .ZN(new_n319_));
  INV_X1    g118(.A(G176gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n310_), .A2(new_n320_), .ZN(new_n321_));
  AOI22_X1  g120(.A1(new_n316_), .A2(new_n317_), .B1(new_n319_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT89), .ZN(new_n323_));
  AND3_X1   g122(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n324_));
  AOI21_X1  g123(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n318_), .A2(new_n310_), .A3(new_n320_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n323_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  AND4_X1   g127(.A1(new_n323_), .A2(new_n327_), .A3(new_n305_), .A4(new_n306_), .ZN(new_n329_));
  OAI211_X1 g128(.A(KEYINPUT90), .B(new_n322_), .C1(new_n328_), .C2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n327_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT89), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n327_), .A2(new_n305_), .A3(new_n323_), .A4(new_n306_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(KEYINPUT90), .B1(new_n335_), .B2(new_n322_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n315_), .B1(new_n331_), .B2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G197gat), .B(G204gat), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT21), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G211gat), .B(G218gat), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(G204gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(G197gat), .ZN(new_n344_));
  INV_X1    g143(.A(G197gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(G204gat), .ZN(new_n346_));
  AND2_X1   g145(.A1(KEYINPUT83), .A2(KEYINPUT21), .ZN(new_n347_));
  NOR2_X1   g146(.A1(KEYINPUT83), .A2(KEYINPUT21), .ZN(new_n348_));
  OAI211_X1 g147(.A(new_n344_), .B(new_n346_), .C1(new_n347_), .C2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT84), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT83), .B(KEYINPUT21), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n338_), .A2(new_n352_), .A3(KEYINPUT84), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n344_), .A2(new_n346_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(KEYINPUT21), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n351_), .A2(new_n353_), .A3(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n342_), .B1(new_n356_), .B2(new_n341_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n337_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT20), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n356_), .A2(new_n341_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n342_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT78), .ZN(new_n363_));
  INV_X1    g162(.A(G183gat), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n363_), .B1(new_n364_), .B2(KEYINPUT25), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT25), .ZN(new_n366_));
  OR2_X1    g165(.A1(new_n366_), .A2(G183gat), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n366_), .A2(KEYINPUT78), .A3(G183gat), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n316_), .A2(new_n365_), .A3(new_n367_), .A4(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n319_), .A2(new_n321_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n369_), .A2(new_n326_), .A3(new_n327_), .A4(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n311_), .A2(KEYINPUT79), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT79), .B1(new_n310_), .B2(KEYINPUT22), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n373_), .A2(new_n320_), .A3(new_n312_), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n308_), .B(new_n307_), .C1(new_n372_), .C2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n371_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n359_), .B1(new_n362_), .B2(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n302_), .B1(new_n358_), .B2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n301_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT20), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n381_), .B1(new_n357_), .B2(new_n376_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n382_), .B1(new_n337_), .B2(new_n357_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n298_), .B1(new_n379_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n298_), .ZN(new_n386_));
  OAI21_X1  g185(.A(KEYINPUT20), .B1(new_n357_), .B2(new_n376_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n387_), .B1(new_n357_), .B2(new_n337_), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n386_), .B(new_n383_), .C1(new_n388_), .C2(new_n302_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n385_), .A2(KEYINPUT92), .A3(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT27), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n379_), .A2(new_n384_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT92), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n392_), .A2(new_n393_), .A3(new_n386_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n390_), .A2(new_n391_), .A3(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT95), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n389_), .A2(KEYINPUT27), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n388_), .A2(new_n302_), .ZN(new_n398_));
  OAI21_X1  g197(.A(KEYINPUT20), .B1(new_n362_), .B2(new_n377_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n322_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n315_), .A2(new_n400_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n401_), .A2(new_n357_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n301_), .B1(new_n399_), .B2(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n386_), .B1(new_n398_), .B2(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n396_), .B1(new_n397_), .B2(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n309_), .A2(new_n314_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT90), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n400_), .A2(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n406_), .B1(new_n408_), .B2(new_n330_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n378_), .B1(new_n362_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n302_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n403_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(new_n298_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n413_), .A2(KEYINPUT95), .A3(KEYINPUT27), .A4(new_n389_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n395_), .A2(new_n405_), .A3(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G225gat), .A2(G233gat), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT4), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT3), .ZN(new_n419_));
  INV_X1    g218(.A(G141gat), .ZN(new_n420_));
  INV_X1    g219(.A(G148gat), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n419_), .A2(new_n420_), .A3(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G141gat), .A2(G148gat), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT2), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n426_));
  NAND3_X1  g225(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n422_), .A2(new_n425_), .A3(new_n426_), .A4(new_n427_), .ZN(new_n428_));
  OR2_X1    g227(.A1(G155gat), .A2(G162gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G155gat), .A2(G162gat), .ZN(new_n430_));
  AND2_X1   g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n428_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n430_), .A2(KEYINPUT1), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT1), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n434_), .A2(G155gat), .A3(G162gat), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n433_), .A2(new_n435_), .A3(new_n429_), .ZN(new_n436_));
  XOR2_X1   g235(.A(G141gat), .B(G148gat), .Z(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n432_), .A2(new_n438_), .ZN(new_n439_));
  OR2_X1    g238(.A1(G127gat), .A2(G134gat), .ZN(new_n440_));
  INV_X1    g239(.A(G113gat), .ZN(new_n441_));
  INV_X1    g240(.A(G120gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G127gat), .A2(G134gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(G113gat), .A2(G120gat), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n440_), .A2(new_n443_), .A3(new_n444_), .A4(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(KEYINPUT80), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n440_), .A2(new_n444_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n443_), .A2(new_n445_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  AND2_X1   g249(.A1(new_n450_), .A2(new_n446_), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n439_), .B(new_n447_), .C1(new_n451_), .C2(KEYINPUT80), .ZN(new_n452_));
  AOI22_X1  g251(.A1(new_n428_), .A2(new_n431_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n450_), .A2(new_n446_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n418_), .B1(new_n452_), .B2(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(KEYINPUT80), .B1(new_n450_), .B2(new_n446_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n447_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(KEYINPUT4), .B1(new_n459_), .B2(new_n439_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n417_), .B1(new_n456_), .B2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n452_), .A2(new_n455_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n416_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n461_), .A2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G1gat), .B(G29gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(new_n213_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(KEYINPUT0), .B(G57gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n465_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n461_), .A2(new_n464_), .A3(new_n469_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT81), .B(KEYINPUT28), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n439_), .A2(KEYINPUT29), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G22gat), .B(G50gat), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n477_), .A2(new_n479_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n476_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n482_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n484_), .A2(new_n475_), .A3(new_n480_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n439_), .A2(KEYINPUT29), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n487_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n360_), .A2(KEYINPUT85), .A3(new_n361_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(KEYINPUT82), .A2(G233gat), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(KEYINPUT82), .A2(G233gat), .ZN(new_n492_));
  OAI21_X1  g291(.A(G228gat), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n488_), .A2(new_n489_), .A3(new_n494_), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n357_), .B(new_n487_), .C1(KEYINPUT85), .C2(new_n493_), .ZN(new_n496_));
  XOR2_X1   g295(.A(G78gat), .B(G106gat), .Z(new_n497_));
  NAND3_X1  g296(.A1(new_n495_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT86), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n495_), .A2(KEYINPUT86), .A3(new_n496_), .A4(new_n497_), .ZN(new_n501_));
  AND2_X1   g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT87), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n495_), .A2(new_n496_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n497_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n503_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  AOI211_X1 g305(.A(KEYINPUT87), .B(new_n497_), .C1(new_n495_), .C2(new_n496_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n486_), .B1(new_n502_), .B2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n504_), .A2(new_n505_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n486_), .A2(new_n510_), .A3(new_n498_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n474_), .B1(new_n509_), .B2(new_n512_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n293_), .B1(new_n415_), .B2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n510_), .A2(KEYINPUT87), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n504_), .A2(new_n503_), .A3(new_n505_), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n515_), .A2(new_n500_), .A3(new_n501_), .A4(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n486_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n473_), .B1(new_n519_), .B2(new_n511_), .ZN(new_n520_));
  AND2_X1   g319(.A1(new_n405_), .A2(new_n414_), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n520_), .A2(new_n521_), .A3(KEYINPUT96), .A4(new_n395_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n512_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT33), .ZN(new_n524_));
  NOR3_X1   g323(.A1(new_n453_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n455_), .ZN(new_n526_));
  OAI21_X1  g325(.A(KEYINPUT4), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n460_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(new_n416_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n469_), .B1(new_n463_), .B2(new_n417_), .ZN(new_n531_));
  AOI22_X1  g330(.A1(new_n472_), .A2(new_n524_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n462_), .A2(new_n417_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n533_), .B1(new_n529_), .B2(new_n417_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT93), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n534_), .A2(new_n535_), .A3(KEYINPUT33), .A4(new_n469_), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n461_), .A2(new_n464_), .A3(KEYINPUT33), .A4(new_n469_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT93), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n532_), .A2(new_n536_), .A3(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n539_), .B1(new_n394_), .B2(new_n390_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT32), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n298_), .A2(new_n541_), .ZN(new_n542_));
  XOR2_X1   g341(.A(new_n542_), .B(KEYINPUT94), .Z(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(new_n392_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n412_), .A2(new_n542_), .ZN(new_n545_));
  AND3_X1   g344(.A1(new_n544_), .A2(new_n473_), .A3(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n523_), .B1(new_n540_), .B2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n514_), .A2(new_n522_), .A3(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G227gat), .A2(G233gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n376_), .B(new_n549_), .ZN(new_n550_));
  XOR2_X1   g349(.A(G71gat), .B(G99gat), .Z(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(KEYINPUT30), .B(G15gat), .ZN(new_n554_));
  XOR2_X1   g353(.A(new_n459_), .B(new_n554_), .Z(new_n555_));
  XOR2_X1   g354(.A(KEYINPUT31), .B(G43gat), .Z(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n553_), .B(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n548_), .A2(new_n559_), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n523_), .A2(new_n395_), .A3(new_n405_), .A4(new_n414_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT97), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n521_), .A2(KEYINPUT97), .A3(new_n523_), .A4(new_n395_), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n563_), .A2(new_n564_), .A3(new_n474_), .A4(new_n558_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n560_), .A2(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n282_), .A2(KEYINPUT12), .A3(new_n225_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n282_), .B1(new_n232_), .B2(new_n234_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G230gat), .A2(G233gat), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n232_), .A2(new_n282_), .A3(new_n234_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT12), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n570_), .A2(new_n571_), .A3(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n282_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n235_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(new_n572_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n571_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n575_), .A2(new_n580_), .ZN(new_n581_));
  XOR2_X1   g380(.A(G176gat), .B(G204gat), .Z(new_n582_));
  XNOR2_X1  g381(.A(G120gat), .B(G148gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n585_));
  XOR2_X1   g384(.A(new_n584_), .B(new_n585_), .Z(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n581_), .A2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n575_), .A2(new_n580_), .A3(new_n586_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n590_), .A2(KEYINPUT13), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(KEYINPUT13), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n205_), .B(KEYINPUT75), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(new_n267_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n267_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n207_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(G229gat), .A2(G233gat), .ZN(new_n599_));
  AND3_X1   g398(.A1(new_n596_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n595_), .B(new_n267_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n599_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n601_), .A2(new_n604_), .ZN(new_n605_));
  XOR2_X1   g404(.A(G169gat), .B(G197gat), .Z(new_n606_));
  XNOR2_X1  g405(.A(G113gat), .B(G141gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n605_), .A2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n601_), .A2(new_n604_), .A3(new_n610_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n594_), .A2(new_n615_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n566_), .A2(new_n616_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n292_), .A2(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n618_), .A2(new_n262_), .A3(new_n473_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT38), .ZN(new_n620_));
  OR2_X1    g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT98), .ZN(new_n622_));
  OR2_X1    g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n250_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n624_), .A2(new_n290_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n617_), .A2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT99), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(G1gat), .B1(new_n628_), .B2(new_n474_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n619_), .A2(new_n620_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n621_), .A2(new_n622_), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n623_), .A2(new_n629_), .A3(new_n630_), .A4(new_n631_), .ZN(G1324gat));
  NAND3_X1  g431(.A1(new_n618_), .A2(new_n263_), .A3(new_n415_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n617_), .A2(new_n415_), .A3(new_n625_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT39), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n634_), .A2(new_n635_), .A3(G8gat), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n635_), .B1(new_n634_), .B2(G8gat), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n633_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  XOR2_X1   g437(.A(new_n638_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g438(.A(G15gat), .B1(new_n628_), .B2(new_n559_), .ZN(new_n640_));
  OR2_X1    g439(.A1(new_n640_), .A2(KEYINPUT41), .ZN(new_n641_));
  INV_X1    g440(.A(G15gat), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n618_), .A2(new_n642_), .A3(new_n558_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT100), .Z(new_n644_));
  NAND2_X1  g443(.A1(new_n640_), .A2(KEYINPUT41), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n641_), .A2(new_n644_), .A3(new_n645_), .ZN(G1326gat));
  XNOR2_X1  g445(.A(new_n523_), .B(KEYINPUT101), .ZN(new_n647_));
  INV_X1    g446(.A(G22gat), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT102), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n618_), .A2(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n648_), .B1(new_n627_), .B2(new_n647_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT42), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n652_), .A2(new_n653_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n651_), .B1(new_n654_), .B2(new_n655_), .ZN(G1327gat));
  INV_X1    g455(.A(KEYINPUT44), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n616_), .A2(new_n290_), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n563_), .A2(new_n558_), .A3(new_n564_), .ZN(new_n659_));
  AOI22_X1  g458(.A1(new_n659_), .A2(new_n474_), .B1(new_n548_), .B2(new_n559_), .ZN(new_n660_));
  OAI21_X1  g459(.A(KEYINPUT43), .B1(new_n660_), .B2(new_n254_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT43), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n566_), .A2(new_n662_), .A3(new_n255_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n658_), .B1(new_n661_), .B2(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n657_), .B1(new_n664_), .B2(KEYINPUT103), .ZN(new_n665_));
  INV_X1    g464(.A(new_n658_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n660_), .A2(KEYINPUT43), .A3(new_n254_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n662_), .B1(new_n566_), .B2(new_n255_), .ZN(new_n668_));
  OAI211_X1 g467(.A(KEYINPUT103), .B(new_n666_), .C1(new_n667_), .C2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  OAI21_X1  g469(.A(KEYINPUT104), .B1(new_n665_), .B2(new_n670_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n666_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT103), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT104), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n674_), .A2(new_n675_), .A3(new_n657_), .A4(new_n669_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n664_), .A2(KEYINPUT44), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n671_), .A2(new_n473_), .A3(new_n676_), .A4(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(G29gat), .ZN(new_n679_));
  INV_X1    g478(.A(new_n290_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n250_), .A2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n617_), .A2(new_n681_), .ZN(new_n682_));
  OR3_X1    g481(.A1(new_n682_), .A2(G29gat), .A3(new_n474_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n679_), .A2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(KEYINPUT105), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT105), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n679_), .A2(new_n686_), .A3(new_n683_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n685_), .A2(new_n687_), .ZN(G1328gat));
  INV_X1    g487(.A(new_n415_), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n682_), .A2(G36gat), .A3(new_n689_), .ZN(new_n690_));
  XOR2_X1   g489(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n691_));
  XNOR2_X1  g490(.A(new_n690_), .B(new_n691_), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n671_), .A2(new_n415_), .A3(new_n676_), .A4(new_n677_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n692_), .B1(new_n693_), .B2(G36gat), .ZN(new_n694_));
  XNOR2_X1  g493(.A(KEYINPUT107), .B(KEYINPUT46), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n695_), .ZN(new_n697_));
  AOI211_X1 g496(.A(new_n697_), .B(new_n692_), .C1(new_n693_), .C2(G36gat), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n696_), .A2(new_n698_), .ZN(G1329gat));
  NAND4_X1  g498(.A1(new_n671_), .A2(new_n558_), .A3(new_n676_), .A4(new_n677_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(G43gat), .ZN(new_n701_));
  OR3_X1    g500(.A1(new_n682_), .A2(G43gat), .A3(new_n559_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT47), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n701_), .A2(KEYINPUT47), .A3(new_n702_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(G1330gat));
  INV_X1    g506(.A(new_n523_), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n671_), .A2(new_n708_), .A3(new_n676_), .A4(new_n677_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(G50gat), .ZN(new_n710_));
  INV_X1    g509(.A(G50gat), .ZN(new_n711_));
  NAND4_X1  g510(.A1(new_n617_), .A2(new_n711_), .A3(new_n647_), .A4(new_n681_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(KEYINPUT108), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT108), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n710_), .A2(new_n715_), .A3(new_n712_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n716_), .ZN(G1331gat));
  NOR2_X1   g516(.A1(new_n593_), .A2(new_n614_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n660_), .A2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(new_n625_), .ZN(new_n721_));
  INV_X1    g520(.A(G57gat), .ZN(new_n722_));
  NOR3_X1   g521(.A1(new_n721_), .A2(new_n722_), .A3(new_n474_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n292_), .A2(new_n720_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(new_n473_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n723_), .B1(new_n726_), .B2(new_n722_), .ZN(G1332gat));
  OAI21_X1  g526(.A(G64gat), .B1(new_n721_), .B2(new_n689_), .ZN(new_n728_));
  XOR2_X1   g527(.A(KEYINPUT109), .B(KEYINPUT48), .Z(new_n729_));
  XNOR2_X1  g528(.A(new_n728_), .B(new_n729_), .ZN(new_n730_));
  OR2_X1    g529(.A1(new_n689_), .A2(G64gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n730_), .B1(new_n724_), .B2(new_n731_), .ZN(G1333gat));
  OAI21_X1  g531(.A(G71gat), .B1(new_n721_), .B2(new_n559_), .ZN(new_n733_));
  XOR2_X1   g532(.A(KEYINPUT110), .B(KEYINPUT49), .Z(new_n734_));
  XNOR2_X1  g533(.A(new_n733_), .B(new_n734_), .ZN(new_n735_));
  OR2_X1    g534(.A1(new_n559_), .A2(G71gat), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n735_), .B1(new_n724_), .B2(new_n736_), .ZN(G1334gat));
  NAND3_X1  g536(.A1(new_n720_), .A2(new_n625_), .A3(new_n647_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(G78gat), .ZN(new_n739_));
  XOR2_X1   g538(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n740_));
  XNOR2_X1  g539(.A(new_n739_), .B(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(G78gat), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n725_), .A2(new_n742_), .A3(new_n647_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(G1335gat));
  AND2_X1   g543(.A1(new_n720_), .A2(new_n681_), .ZN(new_n745_));
  AOI21_X1  g544(.A(G85gat), .B1(new_n745_), .B2(new_n473_), .ZN(new_n746_));
  AOI211_X1 g545(.A(new_n680_), .B(new_n719_), .C1(new_n661_), .C2(new_n663_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n474_), .A2(new_n213_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n746_), .B1(new_n747_), .B2(new_n748_), .ZN(G1336gat));
  AOI21_X1  g548(.A(G92gat), .B1(new_n745_), .B2(new_n415_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n689_), .A2(new_n214_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(new_n747_), .B2(new_n751_), .ZN(G1337gat));
  NAND3_X1  g551(.A1(new_n745_), .A2(new_n208_), .A3(new_n558_), .ZN(new_n753_));
  OR2_X1    g552(.A1(new_n753_), .A2(KEYINPUT112), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(KEYINPUT112), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n747_), .A2(new_n558_), .ZN(new_n756_));
  AOI22_X1  g555(.A1(new_n754_), .A2(new_n755_), .B1(G99gat), .B2(new_n756_), .ZN(new_n757_));
  XOR2_X1   g556(.A(new_n757_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g557(.A1(new_n745_), .A2(new_n209_), .A3(new_n708_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n747_), .A2(new_n708_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(G106gat), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n761_), .A2(KEYINPUT52), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n761_), .A2(KEYINPUT52), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n759_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(KEYINPUT53), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT53), .ZN(new_n766_));
  OAI211_X1 g565(.A(new_n766_), .B(new_n759_), .C1(new_n762_), .C2(new_n763_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n765_), .A2(new_n767_), .ZN(G1339gat));
  INV_X1    g567(.A(new_n659_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n614_), .A2(new_n589_), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n570_), .A2(KEYINPUT55), .A3(new_n571_), .A4(new_n574_), .ZN(new_n771_));
  OR2_X1    g570(.A1(new_n771_), .A2(KEYINPUT114), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(KEYINPUT114), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT55), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n575_), .A2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n570_), .A2(new_n574_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n579_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n772_), .A2(new_n773_), .A3(new_n775_), .A4(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(KEYINPUT56), .B1(new_n778_), .B2(new_n587_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(KEYINPUT115), .A2(KEYINPUT56), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n770_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n773_), .A2(new_n775_), .A3(new_n777_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n771_), .A2(KEYINPUT114), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n587_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT56), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n778_), .A2(KEYINPUT56), .A3(new_n587_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n786_), .A2(KEYINPUT115), .A3(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n781_), .A2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n602_), .A2(new_n599_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n596_), .A2(new_n598_), .A3(new_n603_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n790_), .A2(new_n611_), .A3(new_n791_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n613_), .A2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(new_n590_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n789_), .A2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n795_), .A2(KEYINPUT57), .A3(new_n250_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT57), .ZN(new_n797_));
  AOI22_X1  g596(.A1(new_n781_), .A2(new_n788_), .B1(new_n590_), .B2(new_n793_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n797_), .B1(new_n798_), .B2(new_n624_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n793_), .A2(new_n589_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n784_), .A2(new_n785_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n801_), .B1(new_n802_), .B2(new_n779_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT116), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n803_), .A2(new_n804_), .A3(KEYINPUT58), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT58), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n800_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n806_), .B1(new_n807_), .B2(KEYINPUT116), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n254_), .B1(new_n805_), .B2(new_n808_), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n796_), .B(new_n799_), .C1(new_n809_), .C2(KEYINPUT117), .ZN(new_n810_));
  AND2_X1   g609(.A1(new_n809_), .A2(KEYINPUT117), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n290_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n594_), .A2(new_n614_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n291_), .A2(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(KEYINPUT113), .B1(new_n814_), .B2(KEYINPUT54), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(KEYINPUT54), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT113), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n291_), .A2(new_n817_), .A3(new_n818_), .A4(new_n813_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n815_), .A2(new_n816_), .A3(new_n819_), .ZN(new_n820_));
  AOI211_X1 g619(.A(new_n474_), .B(new_n769_), .C1(new_n812_), .C2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(G113gat), .B1(new_n821_), .B2(new_n614_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n805_), .A2(new_n808_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n255_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n824_), .A2(new_n796_), .A3(new_n799_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n290_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n820_), .ZN(new_n827_));
  XOR2_X1   g626(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n828_));
  NOR3_X1   g627(.A1(new_n769_), .A2(new_n474_), .A3(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n827_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT59), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n830_), .B1(new_n821_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n615_), .A2(new_n441_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n822_), .B1(new_n833_), .B2(new_n834_), .ZN(G1340gat));
  OAI21_X1  g634(.A(G120gat), .B1(new_n832_), .B2(new_n593_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n442_), .B1(new_n593_), .B2(KEYINPUT60), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n821_), .B(new_n837_), .C1(KEYINPUT60), .C2(new_n442_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n838_), .ZN(G1341gat));
  AOI21_X1  g638(.A(G127gat), .B1(new_n821_), .B2(new_n680_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n680_), .A2(G127gat), .ZN(new_n841_));
  XOR2_X1   g640(.A(new_n841_), .B(KEYINPUT119), .Z(new_n842_));
  AOI21_X1  g641(.A(new_n840_), .B1(new_n833_), .B2(new_n842_), .ZN(G1342gat));
  AOI21_X1  g642(.A(G134gat), .B1(new_n821_), .B2(new_n624_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n255_), .A2(G134gat), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n844_), .B1(new_n833_), .B2(new_n845_), .ZN(G1343gat));
  NOR3_X1   g645(.A1(new_n415_), .A2(new_n558_), .A3(new_n523_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  AOI211_X1 g647(.A(new_n474_), .B(new_n848_), .C1(new_n812_), .C2(new_n820_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n614_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(KEYINPUT120), .B(G141gat), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n850_), .B(new_n851_), .ZN(G1344gat));
  NAND2_X1  g651(.A1(new_n849_), .A2(new_n594_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g653(.A(KEYINPUT61), .B(G155gat), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT121), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n857_), .B1(new_n849_), .B2(new_n680_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n812_), .A2(new_n820_), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n859_), .A2(new_n473_), .A3(new_n680_), .A4(new_n847_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n860_), .A2(KEYINPUT121), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n856_), .B1(new_n858_), .B2(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n849_), .A2(new_n857_), .A3(new_n680_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n860_), .A2(KEYINPUT121), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n863_), .A2(new_n864_), .A3(new_n855_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n862_), .A2(new_n865_), .ZN(G1346gat));
  AOI21_X1  g665(.A(G162gat), .B1(new_n849_), .B2(new_n624_), .ZN(new_n867_));
  AND2_X1   g666(.A1(new_n255_), .A2(G162gat), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n867_), .B1(new_n849_), .B2(new_n868_), .ZN(G1347gat));
  INV_X1    g668(.A(KEYINPUT62), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n558_), .A2(new_n474_), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n647_), .A2(new_n689_), .A3(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n873_), .B1(new_n826_), .B2(new_n820_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n614_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n870_), .B1(new_n875_), .B2(G169gat), .ZN(new_n876_));
  AOI211_X1 g675(.A(KEYINPUT62), .B(new_n310_), .C1(new_n874_), .C2(new_n614_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n874_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n615_), .A2(new_n313_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(KEYINPUT122), .ZN(new_n880_));
  OAI22_X1  g679(.A1(new_n876_), .A2(new_n877_), .B1(new_n878_), .B2(new_n880_), .ZN(G1348gat));
  AOI21_X1  g680(.A(G176gat), .B1(new_n874_), .B2(new_n594_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n871_), .A2(new_n708_), .ZN(new_n883_));
  AND3_X1   g682(.A1(new_n859_), .A2(new_n415_), .A3(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n593_), .A2(new_n320_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n882_), .B1(new_n884_), .B2(new_n885_), .ZN(G1349gat));
  NOR3_X1   g685(.A1(new_n878_), .A2(new_n317_), .A3(new_n290_), .ZN(new_n887_));
  NAND4_X1  g686(.A1(new_n859_), .A2(new_n415_), .A3(new_n680_), .A4(new_n883_), .ZN(new_n888_));
  OR2_X1    g687(.A1(new_n888_), .A2(KEYINPUT123), .ZN(new_n889_));
  AOI21_X1  g688(.A(G183gat), .B1(new_n888_), .B2(KEYINPUT123), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n887_), .B1(new_n889_), .B2(new_n890_), .ZN(G1350gat));
  NAND2_X1  g690(.A1(new_n874_), .A2(new_n255_), .ZN(new_n892_));
  AND2_X1   g691(.A1(new_n624_), .A2(new_n316_), .ZN(new_n893_));
  AOI22_X1  g692(.A1(new_n892_), .A2(G190gat), .B1(new_n874_), .B2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT124), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n894_), .B(new_n895_), .ZN(G1351gat));
  NOR2_X1   g695(.A1(new_n513_), .A2(new_n558_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  AOI211_X1 g697(.A(new_n689_), .B(new_n898_), .C1(new_n812_), .C2(new_n820_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n899_), .A2(G197gat), .A3(new_n614_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(KEYINPUT125), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n899_), .A2(new_n614_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(new_n345_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT125), .ZN(new_n904_));
  NAND4_X1  g703(.A1(new_n899_), .A2(new_n904_), .A3(G197gat), .A4(new_n614_), .ZN(new_n905_));
  AND3_X1   g704(.A1(new_n901_), .A2(new_n903_), .A3(new_n905_), .ZN(G1352gat));
  NAND2_X1  g705(.A1(new_n899_), .A2(new_n594_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g707(.A(KEYINPUT63), .ZN(new_n909_));
  INV_X1    g708(.A(G211gat), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT126), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n290_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n912_), .B1(new_n899_), .B2(new_n913_), .ZN(new_n914_));
  NAND4_X1  g713(.A1(new_n859_), .A2(new_n415_), .A3(new_n897_), .A4(new_n913_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n915_), .A2(KEYINPUT126), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n911_), .B1(new_n914_), .B2(new_n916_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n899_), .A2(new_n912_), .A3(new_n913_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n915_), .A2(KEYINPUT126), .ZN(new_n919_));
  NAND4_X1  g718(.A1(new_n918_), .A2(new_n919_), .A3(new_n909_), .A4(new_n910_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n917_), .A2(new_n920_), .ZN(G1354gat));
  AOI21_X1  g720(.A(G218gat), .B1(new_n899_), .B2(new_n624_), .ZN(new_n922_));
  AND2_X1   g721(.A1(new_n255_), .A2(G218gat), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n922_), .B1(new_n899_), .B2(new_n923_), .ZN(G1355gat));
endmodule


