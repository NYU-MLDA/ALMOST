//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 0 0 0 0 0 1 1 0 1 0 0 1 1 0 0 1 0 0 1 1 1 1 0 1 1 1 0 1 1 1 1 0 0 0 0 1 0 0 1 0 0 1 1 1 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n766_, new_n767_, new_n768_, new_n770_,
    new_n771_, new_n772_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n785_, new_n786_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n885_, new_n887_, new_n888_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n903_, new_n904_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_, new_n924_, new_n926_, new_n927_, new_n929_, new_n930_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n938_,
    new_n940_, new_n941_, new_n942_, new_n944_, new_n945_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT66), .ZN(new_n204_));
  XOR2_X1   g003(.A(G57gat), .B(G64gat), .Z(new_n205_));
  INV_X1    g004(.A(KEYINPUT11), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(G71gat), .ZN(new_n208_));
  INV_X1    g007(.A(G78gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G71gat), .A2(G78gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n207_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT65), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n205_), .A2(new_n206_), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  OR2_X1    g015(.A1(new_n212_), .A2(KEYINPUT65), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n212_), .A2(KEYINPUT65), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n217_), .A2(new_n218_), .A3(new_n214_), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n216_), .A2(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(G99gat), .A2(G106gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n221_), .B(KEYINPUT7), .ZN(new_n222_));
  OR2_X1    g021(.A1(new_n222_), .A2(KEYINPUT64), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(KEYINPUT64), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G99gat), .A2(G106gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(KEYINPUT6), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n223_), .A2(new_n224_), .A3(new_n226_), .ZN(new_n227_));
  XOR2_X1   g026(.A(G85gat), .B(G92gat), .Z(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(KEYINPUT8), .A3(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT8), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n222_), .A2(new_n226_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n228_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n230_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT9), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n234_), .A2(G85gat), .A3(G92gat), .ZN(new_n235_));
  AND2_X1   g034(.A1(new_n226_), .A2(new_n235_), .ZN(new_n236_));
  XOR2_X1   g035(.A(KEYINPUT10), .B(G99gat), .Z(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  OAI221_X1 g037(.A(new_n236_), .B1(new_n234_), .B2(new_n232_), .C1(G106gat), .C2(new_n238_), .ZN(new_n239_));
  AND3_X1   g038(.A1(new_n229_), .A2(new_n233_), .A3(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n204_), .B1(new_n220_), .B2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n216_), .A2(new_n219_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n229_), .A2(new_n233_), .A3(new_n239_), .ZN(new_n243_));
  NOR3_X1   g042(.A1(new_n242_), .A2(KEYINPUT66), .A3(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n241_), .A2(new_n244_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n220_), .A2(new_n240_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n203_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT12), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n248_), .B1(new_n220_), .B2(new_n240_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n220_), .A2(new_n240_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n242_), .A2(KEYINPUT12), .A3(new_n243_), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n249_), .A2(new_n202_), .A3(new_n250_), .A4(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G120gat), .B(G148gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT5), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(G176gat), .ZN(new_n255_));
  INV_X1    g054(.A(G204gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n255_), .B(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT67), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n247_), .A2(new_n252_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n258_), .B1(new_n247_), .B2(new_n252_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT13), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT13), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n264_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n265_));
  AND2_X1   g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT91), .ZN(new_n268_));
  AND2_X1   g067(.A1(G211gat), .A2(G218gat), .ZN(new_n269_));
  NOR2_X1   g068(.A1(G211gat), .A2(G218gat), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n268_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(G211gat), .ZN(new_n272_));
  INV_X1    g071(.A(G218gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G211gat), .A2(G218gat), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n274_), .A2(KEYINPUT91), .A3(new_n275_), .ZN(new_n276_));
  AND2_X1   g075(.A1(new_n271_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT92), .ZN(new_n278_));
  INV_X1    g077(.A(G197gat), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n279_), .A2(G204gat), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT88), .B(G197gat), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n281_), .B1(new_n282_), .B2(new_n256_), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n277_), .A2(new_n278_), .A3(KEYINPUT21), .A4(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n271_), .A2(new_n276_), .A3(KEYINPUT21), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n279_), .A2(KEYINPUT88), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT88), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(G197gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n280_), .B1(new_n289_), .B2(G204gat), .ZN(new_n290_));
  OAI21_X1  g089(.A(KEYINPUT92), .B1(new_n285_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n284_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G197gat), .A2(G204gat), .ZN(new_n293_));
  OAI211_X1 g092(.A(KEYINPUT21), .B(new_n293_), .C1(new_n282_), .C2(G204gat), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT89), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT90), .B(KEYINPUT21), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n290_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n289_), .A2(new_n256_), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n299_), .A2(KEYINPUT89), .A3(KEYINPUT21), .A4(new_n293_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n271_), .A2(new_n276_), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n296_), .A2(new_n298_), .A3(new_n300_), .A4(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n292_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(G183gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT25), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT25), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(G183gat), .ZN(new_n307_));
  AND2_X1   g106(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n308_));
  NOR2_X1   g107(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n305_), .B(new_n307_), .C1(new_n308_), .C2(new_n309_), .ZN(new_n310_));
  AND3_X1   g109(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n311_));
  AOI21_X1  g110(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(G169gat), .ZN(new_n314_));
  INV_X1    g113(.A(G176gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G169gat), .A2(G176gat), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n316_), .A2(KEYINPUT24), .A3(new_n317_), .ZN(new_n318_));
  OR3_X1    g117(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n310_), .A2(new_n313_), .A3(new_n318_), .A4(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G183gat), .A2(G190gat), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT23), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  OR2_X1    g122(.A1(G183gat), .A2(G190gat), .ZN(new_n324_));
  NAND3_X1  g123(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n323_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n314_), .A2(KEYINPUT22), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT22), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(G169gat), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n327_), .A2(new_n329_), .A3(new_n315_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n326_), .A2(new_n330_), .A3(new_n317_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n320_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n303_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G226gat), .A2(G233gat), .ZN(new_n334_));
  XOR2_X1   g133(.A(new_n334_), .B(KEYINPUT93), .Z(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT19), .ZN(new_n336_));
  AND3_X1   g135(.A1(new_n313_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT26), .B(G190gat), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT75), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n305_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT25), .B(G183gat), .ZN(new_n341_));
  OAI211_X1 g140(.A(new_n338_), .B(new_n340_), .C1(new_n341_), .C2(new_n339_), .ZN(new_n342_));
  AND2_X1   g141(.A1(new_n326_), .A2(new_n317_), .ZN(new_n343_));
  OAI21_X1  g142(.A(KEYINPUT76), .B1(new_n328_), .B2(G169gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT22), .B(G169gat), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n315_), .B(new_n344_), .C1(new_n345_), .C2(KEYINPUT76), .ZN(new_n346_));
  AOI22_X1  g145(.A1(new_n337_), .A2(new_n342_), .B1(new_n343_), .B2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n292_), .A2(new_n302_), .A3(new_n347_), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n333_), .A2(KEYINPUT20), .A3(new_n336_), .A4(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n332_), .ZN(new_n350_));
  AND3_X1   g149(.A1(new_n292_), .A2(new_n302_), .A3(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n347_), .B1(new_n292_), .B2(new_n302_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT20), .ZN(new_n353_));
  NOR3_X1   g152(.A1(new_n351_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n349_), .B1(new_n354_), .B2(new_n336_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G8gat), .B(G36gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(KEYINPUT18), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(G64gat), .ZN(new_n358_));
  INV_X1    g157(.A(G92gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n355_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n352_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n292_), .A2(new_n302_), .A3(new_n350_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n362_), .A2(KEYINPUT20), .A3(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n336_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n360_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n366_), .A2(new_n349_), .A3(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(KEYINPUT27), .B1(new_n361_), .B2(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n367_), .B1(new_n366_), .B2(new_n349_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n332_), .A2(KEYINPUT97), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT97), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n320_), .A2(new_n372_), .A3(new_n331_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n292_), .A2(new_n302_), .A3(new_n371_), .A4(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT98), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n374_), .A2(new_n375_), .A3(KEYINPUT20), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(new_n362_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n375_), .B1(new_n374_), .B2(KEYINPUT20), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n336_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n333_), .A2(KEYINPUT20), .A3(new_n365_), .A4(new_n348_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n370_), .B1(new_n381_), .B2(new_n367_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n369_), .B1(new_n382_), .B2(KEYINPUT27), .ZN(new_n383_));
  INV_X1    g182(.A(G120gat), .ZN(new_n384_));
  INV_X1    g183(.A(G127gat), .ZN(new_n385_));
  INV_X1    g184(.A(G134gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G127gat), .A2(G134gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT79), .ZN(new_n390_));
  INV_X1    g189(.A(G113gat), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT79), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n387_), .A2(new_n392_), .A3(new_n388_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n390_), .A2(new_n391_), .A3(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n391_), .B1(new_n390_), .B2(new_n393_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n384_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n390_), .A2(new_n393_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(G113gat), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n399_), .A2(G120gat), .A3(new_n394_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n397_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT85), .ZN(new_n402_));
  INV_X1    g201(.A(G141gat), .ZN(new_n403_));
  INV_X1    g202(.A(G148gat), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n402_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT3), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT85), .B1(G141gat), .B2(G148gat), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n405_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT86), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n405_), .A2(KEYINPUT86), .A3(new_n406_), .A4(new_n407_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G141gat), .A2(G148gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(KEYINPUT2), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT2), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n415_), .A2(G141gat), .A3(G148gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n403_), .A2(new_n404_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT3), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n412_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT87), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT83), .ZN(new_n424_));
  INV_X1    g223(.A(G155gat), .ZN(new_n425_));
  INV_X1    g224(.A(G162gat), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n424_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT83), .B1(G155gat), .B2(G162gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n420_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT87), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n430_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G155gat), .A2(G162gat), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n423_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(KEYINPUT1), .ZN(new_n436_));
  INV_X1    g235(.A(new_n428_), .ZN(new_n437_));
  NOR3_X1   g236(.A1(KEYINPUT83), .A2(G155gat), .A3(G162gat), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n436_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT84), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n429_), .A2(KEYINPUT84), .A3(new_n436_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n434_), .A2(KEYINPUT1), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n418_), .B(new_n413_), .C1(new_n443_), .C2(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n401_), .B1(new_n435_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT96), .ZN(new_n447_));
  OR2_X1    g246(.A1(KEYINPUT95), .A2(KEYINPUT4), .ZN(new_n448_));
  NAND2_X1  g247(.A1(KEYINPUT95), .A2(KEYINPUT4), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n446_), .A2(new_n447_), .A3(new_n448_), .A4(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n412_), .A2(new_n432_), .A3(new_n421_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(new_n429_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n434_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n445_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  AND2_X1   g253(.A1(new_n397_), .A2(new_n400_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n454_), .A2(new_n455_), .A3(new_n448_), .A4(new_n449_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT96), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n450_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G225gat), .A2(G233gat), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n454_), .A2(new_n455_), .ZN(new_n461_));
  OAI211_X1 g260(.A(new_n401_), .B(new_n445_), .C1(new_n452_), .C2(new_n453_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n461_), .A2(new_n462_), .A3(KEYINPUT4), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT94), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT94), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n461_), .A2(new_n462_), .A3(new_n465_), .A4(KEYINPUT4), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n458_), .A2(new_n460_), .A3(new_n464_), .A4(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G1gat), .B(G29gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(G85gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n469_), .B(KEYINPUT0), .ZN(new_n470_));
  INV_X1    g269(.A(G57gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n470_), .B(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n461_), .A2(new_n462_), .A3(new_n459_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n467_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n467_), .A2(new_n473_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n472_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n383_), .A2(new_n474_), .A3(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G78gat), .B(G106gat), .ZN(new_n479_));
  AOI22_X1  g278(.A1(new_n454_), .A2(KEYINPUT29), .B1(new_n302_), .B2(new_n292_), .ZN(new_n480_));
  INV_X1    g279(.A(G50gat), .ZN(new_n481_));
  AND2_X1   g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n480_), .A2(new_n481_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n479_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  OR2_X1    g283(.A1(new_n480_), .A2(new_n481_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n479_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n480_), .A2(new_n481_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n485_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n484_), .A2(new_n488_), .ZN(new_n489_));
  OR3_X1    g288(.A1(new_n454_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT28), .B1(new_n454_), .B2(KEYINPUT29), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G228gat), .A2(G233gat), .ZN(new_n492_));
  INV_X1    g291(.A(G22gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  AND3_X1   g294(.A1(new_n490_), .A2(new_n491_), .A3(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n495_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n489_), .B(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n478_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G227gat), .A2(G233gat), .ZN(new_n501_));
  XOR2_X1   g300(.A(new_n501_), .B(KEYINPUT30), .Z(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(KEYINPUT76), .B1(new_n327_), .B2(new_n329_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n344_), .A2(new_n315_), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n317_), .B(new_n326_), .C1(new_n504_), .C2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT77), .ZN(new_n507_));
  INV_X1    g306(.A(new_n342_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n313_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n506_), .B(new_n507_), .C1(new_n508_), .C2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n337_), .A2(new_n342_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n507_), .B1(new_n512_), .B2(new_n506_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n503_), .B1(new_n511_), .B2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(KEYINPUT78), .B(G43gat), .ZN(new_n515_));
  XOR2_X1   g314(.A(new_n515_), .B(G99gat), .Z(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n506_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT77), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n519_), .A2(new_n510_), .A3(new_n502_), .ZN(new_n520_));
  AND3_X1   g319(.A1(new_n514_), .A2(new_n517_), .A3(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n517_), .B1(new_n514_), .B2(new_n520_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G15gat), .B(G71gat), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NOR3_X1   g323(.A1(new_n521_), .A2(new_n522_), .A3(new_n524_), .ZN(new_n525_));
  NOR3_X1   g324(.A1(new_n511_), .A2(new_n513_), .A3(new_n503_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n502_), .B1(new_n519_), .B2(new_n510_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n516_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n514_), .A2(new_n517_), .A3(new_n520_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n523_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  OAI21_X1  g329(.A(KEYINPUT81), .B1(new_n525_), .B2(new_n530_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n524_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT81), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n528_), .A2(new_n523_), .A3(new_n529_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n532_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n535_));
  XOR2_X1   g334(.A(KEYINPUT80), .B(KEYINPUT31), .Z(new_n536_));
  XNOR2_X1  g335(.A(new_n401_), .B(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n531_), .A2(new_n535_), .A3(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n537_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n532_), .A2(new_n534_), .A3(new_n533_), .A4(new_n539_), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n538_), .A2(KEYINPUT82), .A3(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(KEYINPUT82), .B1(new_n538_), .B2(new_n540_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n500_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n360_), .A2(KEYINPUT32), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n546_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n547_), .B1(new_n355_), .B2(new_n546_), .ZN(new_n548_));
  AND3_X1   g347(.A1(new_n467_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n472_), .B1(new_n467_), .B2(new_n473_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n548_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(KEYINPUT99), .ZN(new_n552_));
  XOR2_X1   g351(.A(new_n489_), .B(new_n498_), .Z(new_n553_));
  INV_X1    g352(.A(KEYINPUT33), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n474_), .A2(new_n554_), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n361_), .A2(new_n368_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n458_), .A2(new_n459_), .A3(new_n464_), .A4(new_n466_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n461_), .A2(new_n462_), .A3(new_n460_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n557_), .A2(new_n476_), .A3(new_n558_), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n467_), .A2(KEYINPUT33), .A3(new_n472_), .A4(new_n473_), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n555_), .A2(new_n556_), .A3(new_n559_), .A4(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT99), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n562_), .B(new_n548_), .C1(new_n549_), .C2(new_n550_), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n552_), .A2(new_n553_), .A3(new_n561_), .A4(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n545_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n538_), .A2(new_n540_), .ZN(new_n566_));
  NOR3_X1   g365(.A1(new_n478_), .A2(new_n499_), .A3(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n565_), .A2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G29gat), .B(G36gat), .ZN(new_n570_));
  INV_X1    g369(.A(G43gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(new_n481_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT15), .ZN(new_n574_));
  XOR2_X1   g373(.A(KEYINPUT70), .B(G1gat), .Z(new_n575_));
  INV_X1    g374(.A(G8gat), .ZN(new_n576_));
  OAI21_X1  g375(.A(KEYINPUT14), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G15gat), .B(G22gat), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(G1gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(G8gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n579_), .B(G1gat), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(new_n576_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n574_), .A2(new_n582_), .A3(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n582_), .A2(new_n584_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(new_n573_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(G229gat), .A2(G233gat), .ZN(new_n588_));
  XOR2_X1   g387(.A(new_n588_), .B(KEYINPUT72), .Z(new_n589_));
  NAND3_X1  g388(.A1(new_n585_), .A2(new_n587_), .A3(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n573_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n586_), .B(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n590_), .B1(new_n592_), .B2(new_n588_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G113gat), .B(G141gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(new_n314_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(new_n279_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n593_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n596_), .ZN(new_n598_));
  OAI211_X1 g397(.A(new_n590_), .B(new_n598_), .C1(new_n592_), .C2(new_n588_), .ZN(new_n599_));
  AND3_X1   g398(.A1(new_n597_), .A2(KEYINPUT73), .A3(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(KEYINPUT73), .B1(new_n597_), .B2(new_n599_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n602_), .A2(KEYINPUT74), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n602_), .A2(KEYINPUT74), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n569_), .A2(KEYINPUT100), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT100), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n567_), .B1(new_n545_), .B2(new_n564_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n608_), .B1(new_n609_), .B2(new_n605_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n267_), .B1(new_n607_), .B2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(G231gat), .A2(G233gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n586_), .B(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(new_n220_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT71), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G127gat), .B(G155gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT16), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(G183gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(new_n272_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT17), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n616_), .B(new_n622_), .Z(new_n623_));
  INV_X1    g422(.A(new_n614_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n624_), .A2(new_n621_), .A3(new_n620_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n574_), .A2(new_n243_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n240_), .A2(new_n573_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(G232gat), .A2(G233gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT34), .ZN(new_n631_));
  OAI211_X1 g430(.A(new_n628_), .B(new_n629_), .C1(KEYINPUT35), .C2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(KEYINPUT35), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT68), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n632_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n632_), .A2(new_n634_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(G190gat), .B(G218gat), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(G134gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(new_n426_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n641_), .A2(KEYINPUT36), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n637_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n642_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n641_), .A2(KEYINPUT36), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n645_), .A2(KEYINPUT37), .A3(new_n648_), .ZN(new_n649_));
  AND3_X1   g448(.A1(new_n646_), .A2(KEYINPUT69), .A3(new_n647_), .ZN(new_n650_));
  AOI21_X1  g449(.A(KEYINPUT69), .B1(new_n646_), .B2(new_n647_), .ZN(new_n651_));
  NOR3_X1   g450(.A1(new_n650_), .A2(new_n651_), .A3(new_n644_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n649_), .B1(new_n652_), .B2(KEYINPUT37), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n627_), .A2(new_n653_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n611_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(new_n575_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n477_), .A2(new_n474_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT102), .ZN(new_n660_));
  OR3_X1    g459(.A1(new_n659_), .A2(new_n660_), .A3(KEYINPUT38), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n659_), .A2(KEYINPUT38), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n660_), .B1(new_n659_), .B2(KEYINPUT38), .ZN(new_n663_));
  OR2_X1    g462(.A1(new_n600_), .A2(new_n601_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n263_), .A2(new_n664_), .A3(new_n265_), .ZN(new_n665_));
  XOR2_X1   g464(.A(new_n665_), .B(KEYINPUT101), .Z(new_n666_));
  NOR2_X1   g465(.A1(new_n609_), .A2(new_n652_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n666_), .A2(new_n626_), .A3(new_n667_), .ZN(new_n668_));
  OAI21_X1  g467(.A(G1gat), .B1(new_n668_), .B2(new_n658_), .ZN(new_n669_));
  NAND4_X1  g468(.A1(new_n661_), .A2(new_n662_), .A3(new_n663_), .A4(new_n669_), .ZN(G1324gat));
  INV_X1    g469(.A(KEYINPUT103), .ZN(new_n671_));
  INV_X1    g470(.A(new_n383_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n611_), .A2(new_n576_), .A3(new_n654_), .A4(new_n672_), .ZN(new_n673_));
  NAND4_X1  g472(.A1(new_n666_), .A2(new_n626_), .A3(new_n672_), .A4(new_n667_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT39), .ZN(new_n675_));
  AND3_X1   g474(.A1(new_n674_), .A2(new_n675_), .A3(G8gat), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n674_), .B2(G8gat), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n673_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(KEYINPUT104), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT104), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n680_), .B(new_n673_), .C1(new_n676_), .C2(new_n677_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n671_), .B1(new_n679_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n679_), .A2(new_n671_), .A3(new_n681_), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n683_), .A2(KEYINPUT40), .A3(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(KEYINPUT40), .B1(new_n683_), .B2(new_n684_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n685_), .A2(new_n686_), .ZN(G1325gat));
  OAI21_X1  g486(.A(G15gat), .B1(new_n668_), .B2(new_n543_), .ZN(new_n688_));
  XOR2_X1   g487(.A(new_n688_), .B(KEYINPUT41), .Z(new_n689_));
  INV_X1    g488(.A(G15gat), .ZN(new_n690_));
  INV_X1    g489(.A(new_n542_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n538_), .A2(KEYINPUT82), .A3(new_n540_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n655_), .A2(new_n690_), .A3(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n689_), .A2(new_n694_), .ZN(G1326gat));
  XNOR2_X1  g494(.A(new_n553_), .B(KEYINPUT105), .ZN(new_n696_));
  OAI21_X1  g495(.A(G22gat), .B1(new_n668_), .B2(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT42), .ZN(new_n698_));
  INV_X1    g497(.A(new_n696_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n655_), .A2(new_n493_), .A3(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n698_), .A2(new_n700_), .ZN(G1327gat));
  INV_X1    g500(.A(KEYINPUT43), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n562_), .B1(new_n657_), .B2(new_n548_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n563_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n553_), .A2(new_n561_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n544_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n702_), .B(new_n653_), .C1(new_n707_), .C2(new_n567_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT106), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n653_), .ZN(new_n711_));
  OAI21_X1  g510(.A(KEYINPUT43), .B1(new_n711_), .B2(new_n609_), .ZN(new_n712_));
  NAND4_X1  g511(.A1(new_n569_), .A2(KEYINPUT106), .A3(new_n702_), .A4(new_n653_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n710_), .A2(new_n712_), .A3(new_n713_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n666_), .A2(new_n627_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(KEYINPUT44), .B1(new_n716_), .B2(KEYINPUT107), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT107), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n719_));
  AOI211_X1 g518(.A(new_n718_), .B(new_n719_), .C1(new_n714_), .C2(new_n715_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n657_), .B1(new_n717_), .B2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(G29gat), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n611_), .A2(new_n652_), .A3(new_n627_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT108), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n611_), .A2(KEYINPUT108), .A3(new_n652_), .A4(new_n627_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(G29gat), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n727_), .A2(new_n728_), .A3(new_n657_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n722_), .A2(new_n729_), .ZN(new_n730_));
  XOR2_X1   g529(.A(new_n730_), .B(KEYINPUT109), .Z(G1328gat));
  OAI21_X1  g530(.A(new_n672_), .B1(new_n717_), .B2(new_n720_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(KEYINPUT110), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT110), .ZN(new_n734_));
  OAI211_X1 g533(.A(new_n734_), .B(new_n672_), .C1(new_n717_), .C2(new_n720_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n733_), .A2(G36gat), .A3(new_n735_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(KEYINPUT111), .B(KEYINPUT46), .ZN(new_n737_));
  INV_X1    g536(.A(G36gat), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n725_), .A2(new_n738_), .A3(new_n672_), .A4(new_n726_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT45), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n736_), .A2(new_n737_), .A3(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n737_), .B1(new_n736_), .B2(new_n740_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n741_), .A2(new_n742_), .ZN(G1329gat));
  NOR2_X1   g542(.A1(new_n717_), .A2(new_n720_), .ZN(new_n744_));
  OAI21_X1  g543(.A(G43gat), .B1(new_n744_), .B2(new_n566_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n727_), .A2(new_n571_), .A3(new_n693_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n747_), .B(new_n749_), .ZN(G1330gat));
  OAI21_X1  g549(.A(G50gat), .B1(new_n744_), .B2(new_n553_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n727_), .A2(new_n481_), .A3(new_n699_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(G1331gat));
  NAND2_X1  g552(.A1(new_n654_), .A2(new_n267_), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT113), .Z(new_n755_));
  NOR3_X1   g554(.A1(new_n755_), .A2(new_n664_), .A3(new_n609_), .ZN(new_n756_));
  AOI21_X1  g555(.A(G57gat), .B1(new_n756_), .B2(new_n657_), .ZN(new_n757_));
  AND4_X1   g556(.A1(new_n626_), .A2(new_n667_), .A3(new_n267_), .A4(new_n605_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n658_), .A2(new_n471_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n757_), .B1(new_n758_), .B2(new_n759_), .ZN(G1332gat));
  INV_X1    g559(.A(G64gat), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n761_), .B1(new_n758_), .B2(new_n672_), .ZN(new_n762_));
  XOR2_X1   g561(.A(new_n762_), .B(KEYINPUT48), .Z(new_n763_));
  NAND3_X1  g562(.A1(new_n756_), .A2(new_n761_), .A3(new_n672_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(G1333gat));
  AOI21_X1  g564(.A(new_n208_), .B1(new_n758_), .B2(new_n693_), .ZN(new_n766_));
  XOR2_X1   g565(.A(new_n766_), .B(KEYINPUT49), .Z(new_n767_));
  NAND3_X1  g566(.A1(new_n756_), .A2(new_n208_), .A3(new_n693_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(G1334gat));
  AOI21_X1  g568(.A(new_n209_), .B1(new_n758_), .B2(new_n699_), .ZN(new_n770_));
  XOR2_X1   g569(.A(new_n770_), .B(KEYINPUT50), .Z(new_n771_));
  NAND3_X1  g570(.A1(new_n756_), .A2(new_n209_), .A3(new_n699_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(G1335gat));
  INV_X1    g572(.A(new_n652_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n609_), .A2(new_n774_), .ZN(new_n775_));
  NOR3_X1   g574(.A1(new_n626_), .A2(new_n266_), .A3(new_n664_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(G85gat), .B1(new_n778_), .B2(new_n657_), .ZN(new_n779_));
  XOR2_X1   g578(.A(new_n779_), .B(KEYINPUT114), .Z(new_n780_));
  AND2_X1   g579(.A1(new_n714_), .A2(new_n776_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n657_), .A2(G85gat), .ZN(new_n782_));
  XOR2_X1   g581(.A(new_n782_), .B(KEYINPUT115), .Z(new_n783_));
  AOI21_X1  g582(.A(new_n780_), .B1(new_n781_), .B2(new_n783_), .ZN(G1336gat));
  AOI21_X1  g583(.A(G92gat), .B1(new_n778_), .B2(new_n672_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n383_), .A2(new_n359_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n785_), .B1(new_n781_), .B2(new_n786_), .ZN(G1337gat));
  NAND2_X1  g586(.A1(new_n781_), .A2(new_n693_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(G99gat), .ZN(new_n789_));
  OR3_X1    g588(.A1(new_n777_), .A2(new_n238_), .A3(new_n566_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  OR2_X1    g590(.A1(new_n791_), .A2(KEYINPUT116), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(KEYINPUT116), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n792_), .A2(KEYINPUT51), .A3(new_n793_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(KEYINPUT117), .B(KEYINPUT51), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n789_), .A2(new_n790_), .A3(new_n795_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT118), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n794_), .A2(new_n797_), .ZN(G1338gat));
  OR3_X1    g597(.A1(new_n777_), .A2(G106gat), .A3(new_n553_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n781_), .A2(new_n499_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT52), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n800_), .A2(new_n801_), .A3(G106gat), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n801_), .B1(new_n800_), .B2(G106gat), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n799_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g604(.A1(new_n658_), .A2(new_n672_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n807_), .A2(new_n566_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n257_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n247_), .A2(new_n252_), .A3(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n810_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n249_), .A2(new_n251_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n203_), .B1(new_n245_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n251_), .ZN(new_n814_));
  AOI21_X1  g613(.A(KEYINPUT12), .B1(new_n242_), .B2(new_n243_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n816_), .A2(KEYINPUT55), .A3(new_n202_), .A4(new_n250_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n252_), .A2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n813_), .A2(new_n817_), .A3(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT119), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n813_), .A2(new_n817_), .A3(KEYINPUT119), .A4(new_n819_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n822_), .A2(new_n257_), .A3(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT56), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n822_), .A2(KEYINPUT56), .A3(new_n257_), .A4(new_n823_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n811_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n585_), .A2(new_n587_), .ZN(new_n829_));
  MUX2_X1   g628(.A(new_n829_), .B(new_n592_), .S(new_n589_), .Z(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n596_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n599_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n262_), .A2(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n774_), .B1(new_n828_), .B2(new_n833_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(KEYINPUT57), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT58), .ZN(new_n836_));
  INV_X1    g635(.A(new_n827_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n826_), .A2(KEYINPUT120), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT120), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n824_), .A2(new_n839_), .A3(new_n825_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n837_), .B1(new_n838_), .B2(new_n840_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n831_), .A2(new_n599_), .A3(new_n810_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n836_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n840_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n839_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n827_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n842_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n846_), .A2(KEYINPUT58), .A3(new_n847_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n843_), .A2(new_n848_), .A3(new_n653_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n626_), .B1(new_n835_), .B2(new_n849_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n711_), .A2(new_n626_), .A3(new_n266_), .A4(new_n605_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n851_), .B(new_n852_), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n553_), .B(new_n808_), .C1(new_n850_), .C2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(G113gat), .B1(new_n855_), .B2(new_n664_), .ZN(new_n856_));
  AND3_X1   g655(.A1(new_n843_), .A2(new_n653_), .A3(new_n848_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n834_), .B(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n627_), .B1(new_n857_), .B2(new_n859_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n851_), .B(KEYINPUT54), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n499_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT59), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n862_), .A2(new_n863_), .A3(new_n808_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n854_), .A2(KEYINPUT59), .ZN(new_n865_));
  AND3_X1   g664(.A1(new_n864_), .A2(KEYINPUT121), .A3(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(KEYINPUT121), .B1(new_n864_), .B2(new_n865_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n605_), .A2(new_n391_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n856_), .B1(new_n868_), .B2(new_n869_), .ZN(G1340gat));
  NOR2_X1   g669(.A1(new_n266_), .A2(G120gat), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n855_), .B1(KEYINPUT60), .B2(new_n871_), .ZN(new_n872_));
  AND4_X1   g671(.A1(new_n267_), .A2(new_n872_), .A3(new_n865_), .A4(new_n864_), .ZN(new_n873_));
  OAI22_X1  g672(.A1(new_n873_), .A2(new_n384_), .B1(KEYINPUT60), .B2(new_n872_), .ZN(G1341gat));
  NAND2_X1  g673(.A1(new_n862_), .A2(new_n626_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n876_), .A2(new_n385_), .A3(new_n808_), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n866_), .A2(new_n867_), .A3(new_n627_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n878_), .B2(new_n385_), .ZN(G1342gat));
  AOI21_X1  g678(.A(G134gat), .B1(new_n855_), .B2(new_n652_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n711_), .A2(new_n386_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n880_), .B1(new_n868_), .B2(new_n881_), .ZN(G1343gat));
  NOR2_X1   g681(.A1(new_n693_), .A2(new_n553_), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n806_), .B(new_n883_), .C1(new_n850_), .C2(new_n853_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(new_n602_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(new_n403_), .ZN(G1344gat));
  NOR2_X1   g685(.A1(new_n884_), .A2(new_n266_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(KEYINPUT122), .B(G148gat), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n887_), .B(new_n888_), .ZN(G1345gat));
  OAI21_X1  g688(.A(KEYINPUT123), .B1(new_n884_), .B2(new_n627_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n807_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT123), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n891_), .A2(new_n892_), .A3(new_n626_), .A4(new_n883_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT61), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n890_), .A2(new_n893_), .A3(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n894_), .B1(new_n890_), .B2(new_n893_), .ZN(new_n897_));
  NOR3_X1   g696(.A1(new_n896_), .A2(new_n897_), .A3(new_n425_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n890_), .A2(new_n893_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(KEYINPUT61), .ZN(new_n900_));
  AOI21_X1  g699(.A(G155gat), .B1(new_n900_), .B2(new_n895_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n898_), .A2(new_n901_), .ZN(G1346gat));
  NOR3_X1   g701(.A1(new_n884_), .A2(new_n426_), .A3(new_n711_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n891_), .A2(new_n652_), .A3(new_n883_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n903_), .B1(new_n426_), .B2(new_n904_), .ZN(G1347gat));
  NAND2_X1  g704(.A1(new_n860_), .A2(new_n861_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n693_), .A2(new_n658_), .A3(new_n672_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(KEYINPUT124), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n906_), .A2(new_n696_), .A3(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n664_), .A2(new_n345_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(KEYINPUT126), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n910_), .A2(new_n912_), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT125), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n914_), .B1(new_n909_), .B2(new_n602_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n699_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n916_));
  NAND4_X1  g715(.A1(new_n916_), .A2(KEYINPUT125), .A3(new_n664_), .A4(new_n908_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n915_), .A2(G169gat), .A3(new_n917_), .ZN(new_n918_));
  AND2_X1   g717(.A1(new_n918_), .A2(KEYINPUT62), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n918_), .A2(KEYINPUT62), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n913_), .B1(new_n919_), .B2(new_n920_), .ZN(G1348gat));
  NAND4_X1  g720(.A1(new_n916_), .A2(new_n315_), .A3(new_n267_), .A4(new_n908_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n862_), .A2(new_n267_), .A3(new_n908_), .ZN(new_n923_));
  INV_X1    g722(.A(new_n923_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n922_), .B1(new_n924_), .B2(new_n315_), .ZN(G1349gat));
  NOR3_X1   g724(.A1(new_n909_), .A2(new_n627_), .A3(new_n341_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n876_), .A2(new_n908_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n926_), .B1(new_n927_), .B2(new_n304_), .ZN(G1350gat));
  NAND3_X1  g727(.A1(new_n910_), .A2(new_n652_), .A3(new_n338_), .ZN(new_n929_));
  OAI21_X1  g728(.A(G190gat), .B1(new_n909_), .B2(new_n711_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n929_), .A2(new_n930_), .ZN(G1351gat));
  AOI21_X1  g730(.A(new_n383_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n883_), .A2(new_n658_), .ZN(new_n933_));
  XOR2_X1   g732(.A(new_n933_), .B(KEYINPUT127), .Z(new_n934_));
  NAND2_X1  g733(.A1(new_n932_), .A2(new_n934_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n935_), .A2(new_n602_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n936_), .B(new_n279_), .ZN(G1352gat));
  NOR2_X1   g736(.A1(new_n935_), .A2(new_n266_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(new_n256_), .ZN(G1353gat));
  NOR2_X1   g738(.A1(new_n935_), .A2(new_n627_), .ZN(new_n940_));
  NOR3_X1   g739(.A1(new_n940_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n941_));
  XOR2_X1   g740(.A(KEYINPUT63), .B(G211gat), .Z(new_n942_));
  AOI21_X1  g741(.A(new_n941_), .B1(new_n940_), .B2(new_n942_), .ZN(G1354gat));
  NOR3_X1   g742(.A1(new_n935_), .A2(new_n273_), .A3(new_n711_), .ZN(new_n944_));
  NAND3_X1  g743(.A1(new_n932_), .A2(new_n652_), .A3(new_n934_), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n944_), .B1(new_n273_), .B2(new_n945_), .ZN(G1355gat));
endmodule


