//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 1 1 1 0 1 1 1 0 0 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 1 0 0 0 0 0 0 0 0 1 0 1 1 0 1 1 1 0 0 1 1 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n735_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n780_, new_n781_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n894_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n925_, new_n926_, new_n928_, new_n929_, new_n930_,
    new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_,
    new_n937_, new_n939_, new_n940_, new_n941_, new_n943_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n952_,
    new_n953_;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n203_), .A2(KEYINPUT88), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT28), .ZN(new_n205_));
  NOR2_X1   g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT3), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G141gat), .A2(G148gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT2), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n207_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n210_), .A2(new_n211_), .A3(new_n213_), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n212_), .B1(KEYINPUT1), .B2(new_n211_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n215_), .B1(KEYINPUT1), .B2(new_n211_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n206_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n216_), .A2(new_n217_), .A3(new_n208_), .ZN(new_n218_));
  AND2_X1   g017(.A1(new_n214_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT29), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n205_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n214_), .A2(new_n218_), .ZN(new_n222_));
  NOR3_X1   g021(.A1(new_n222_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G22gat), .B(G50gat), .ZN(new_n224_));
  NOR3_X1   g023(.A1(new_n221_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n224_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n219_), .A2(new_n205_), .A3(new_n220_), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT28), .B1(new_n222_), .B2(KEYINPUT29), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n226_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n204_), .B1(new_n225_), .B2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(G197gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(G204gat), .ZN(new_n232_));
  INV_X1    g031(.A(G204gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(G197gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n232_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(G218gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(G211gat), .ZN(new_n237_));
  INV_X1    g036(.A(G211gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(G218gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n235_), .A2(new_n240_), .A3(KEYINPUT21), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n231_), .A2(KEYINPUT86), .A3(G204gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT21), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT86), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G197gat), .B(G204gat), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n243_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G211gat), .B(G218gat), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n247_), .B1(new_n235_), .B2(KEYINPUT21), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n241_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n249_));
  XOR2_X1   g048(.A(KEYINPUT87), .B(KEYINPUT29), .Z(new_n250_));
  OAI21_X1  g049(.A(new_n249_), .B1(new_n219_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(G228gat), .ZN(new_n252_));
  INV_X1    g051(.A(G233gat), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n253_), .A2(KEYINPUT85), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(KEYINPUT85), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n252_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n251_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT21), .ZN(new_n258_));
  NOR3_X1   g057(.A1(new_n245_), .A2(new_n247_), .A3(new_n258_), .ZN(new_n259_));
  OAI211_X1 g058(.A(KEYINPUT21), .B(new_n242_), .C1(new_n235_), .C2(KEYINPUT86), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n240_), .B1(new_n258_), .B2(new_n245_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n259_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n262_), .A2(new_n256_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n263_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n257_), .A2(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n224_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n227_), .A2(new_n228_), .A3(new_n226_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n266_), .A2(new_n203_), .A3(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n230_), .A2(new_n265_), .A3(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n265_), .B1(new_n230_), .B2(new_n268_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  XOR2_X1   g072(.A(G127gat), .B(G134gat), .Z(new_n274_));
  XOR2_X1   g073(.A(G113gat), .B(G120gat), .Z(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n222_), .A2(new_n277_), .ZN(new_n278_));
  OR2_X1    g077(.A1(new_n278_), .A2(KEYINPUT4), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n214_), .A2(new_n276_), .A3(new_n218_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n278_), .A2(KEYINPUT4), .A3(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G225gat), .A2(G233gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT95), .ZN(new_n283_));
  XOR2_X1   g082(.A(new_n283_), .B(KEYINPUT96), .Z(new_n284_));
  NAND3_X1  g083(.A1(new_n279_), .A2(new_n281_), .A3(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n283_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n278_), .A2(new_n280_), .A3(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G1gat), .B(G29gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(G85gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT0), .B(G57gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n285_), .A2(new_n287_), .A3(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT33), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  AND3_X1   g094(.A1(new_n279_), .A2(new_n286_), .A3(new_n281_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n278_), .A2(new_n280_), .A3(new_n284_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(new_n291_), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT33), .B1(new_n296_), .B2(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n295_), .B1(new_n293_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(G183gat), .ZN(new_n301_));
  INV_X1    g100(.A(G190gat), .ZN(new_n302_));
  OAI21_X1  g101(.A(KEYINPUT23), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT23), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n304_), .A2(G183gat), .A3(G190gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT24), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(KEYINPUT91), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT91), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT24), .ZN(new_n310_));
  NOR2_X1   g109(.A1(G169gat), .A2(G176gat), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n308_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n308_), .A2(new_n310_), .ZN(new_n313_));
  INV_X1    g112(.A(G169gat), .ZN(new_n314_));
  INV_X1    g113(.A(G176gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G169gat), .A2(G176gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n306_), .B(new_n312_), .C1(new_n313_), .C2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n301_), .A2(KEYINPUT25), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT25), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(G183gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT90), .ZN(new_n324_));
  NAND2_X1  g123(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n324_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT26), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(new_n302_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n330_), .A2(KEYINPUT90), .A3(new_n325_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n323_), .B1(new_n328_), .B2(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n319_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT22), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n334_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n335_));
  OAI21_X1  g134(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n304_), .B1(G183gat), .B2(G190gat), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT83), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n305_), .A2(new_n340_), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n304_), .A2(KEYINPUT83), .A3(G183gat), .A4(G190gat), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n339_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(G183gat), .A2(G190gat), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n338_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT92), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  OAI211_X1 g146(.A(KEYINPUT92), .B(new_n338_), .C1(new_n343_), .C2(new_n344_), .ZN(new_n348_));
  AOI211_X1 g147(.A(new_n249_), .B(new_n333_), .C1(new_n347_), .C2(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G226gat), .A2(G233gat), .ZN(new_n351_));
  XOR2_X1   g150(.A(new_n350_), .B(new_n351_), .Z(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT81), .B(G190gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(new_n301_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n337_), .B1(new_n354_), .B2(new_n306_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n330_), .B1(new_n353_), .B2(new_n329_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(KEYINPUT80), .A2(G183gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(new_n321_), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n359_));
  AND2_X1   g158(.A1(G169gat), .A2(G176gat), .ZN(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT82), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT82), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n316_), .A2(new_n362_), .A3(KEYINPUT24), .A4(new_n317_), .ZN(new_n363_));
  AOI22_X1  g162(.A1(new_n356_), .A2(new_n358_), .B1(new_n361_), .B2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n341_), .A2(new_n342_), .ZN(new_n365_));
  AOI22_X1  g164(.A1(new_n365_), .A2(new_n303_), .B1(new_n307_), .B2(new_n311_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n355_), .B1(new_n364_), .B2(new_n366_), .ZN(new_n367_));
  OAI211_X1 g166(.A(KEYINPUT20), .B(new_n352_), .C1(new_n367_), .C2(new_n262_), .ZN(new_n368_));
  OAI21_X1  g167(.A(KEYINPUT93), .B1(new_n349_), .B2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n347_), .A2(new_n348_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n323_), .ZN(new_n371_));
  NOR3_X1   g170(.A1(new_n326_), .A2(new_n327_), .A3(new_n324_), .ZN(new_n372_));
  AOI21_X1  g171(.A(KEYINPUT90), .B1(new_n330_), .B2(new_n325_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n371_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n308_), .A2(new_n310_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n375_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n374_), .A2(new_n306_), .A3(new_n312_), .A4(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n370_), .A2(new_n262_), .A3(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT20), .ZN(new_n379_));
  INV_X1    g178(.A(new_n355_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n365_), .A2(new_n303_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n311_), .A2(new_n307_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n361_), .A2(new_n363_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n302_), .A2(KEYINPUT81), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT81), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(G190gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n385_), .A2(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n327_), .B1(new_n388_), .B2(KEYINPUT26), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n357_), .B(KEYINPUT25), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n384_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n380_), .B1(new_n383_), .B2(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n379_), .B1(new_n392_), .B2(new_n249_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT93), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n378_), .A2(new_n393_), .A3(new_n394_), .A4(new_n352_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n352_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n379_), .B1(new_n367_), .B2(new_n262_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n333_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n397_), .B1(new_n262_), .B2(new_n398_), .ZN(new_n399_));
  AOI22_X1  g198(.A1(new_n369_), .A2(new_n395_), .B1(new_n396_), .B2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G8gat), .B(G36gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT18), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G64gat), .B(G92gat), .ZN(new_n403_));
  XOR2_X1   g202(.A(new_n402_), .B(new_n403_), .Z(new_n404_));
  NAND3_X1  g203(.A1(new_n400_), .A2(KEYINPUT94), .A3(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n369_), .A2(new_n395_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n399_), .A2(new_n396_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n404_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n406_), .A2(new_n404_), .A3(new_n407_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT94), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n300_), .A2(new_n405_), .A3(new_n410_), .A4(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n292_), .B1(new_n285_), .B2(new_n287_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(new_n293_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n377_), .A2(new_n262_), .A3(new_n345_), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n418_), .B(KEYINPUT20), .C1(new_n367_), .C2(new_n262_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(new_n396_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(KEYINPUT97), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n397_), .B(new_n352_), .C1(new_n262_), .C2(new_n398_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT97), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n419_), .A2(new_n423_), .A3(new_n396_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n421_), .A2(new_n422_), .A3(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n404_), .A2(KEYINPUT32), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n425_), .A2(new_n427_), .ZN(new_n428_));
  OAI211_X1 g227(.A(new_n417_), .B(new_n428_), .C1(new_n427_), .C2(new_n408_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n273_), .B1(new_n414_), .B2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n424_), .A2(new_n422_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n423_), .B1(new_n419_), .B2(new_n396_), .ZN(new_n432_));
  OAI211_X1 g231(.A(KEYINPUT98), .B(new_n409_), .C1(new_n431_), .C2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(KEYINPUT98), .B1(new_n425_), .B2(new_n409_), .ZN(new_n435_));
  OAI21_X1  g234(.A(KEYINPUT27), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT99), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n411_), .A2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n400_), .A2(KEYINPUT99), .A3(new_n404_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(KEYINPUT100), .B1(new_n436_), .B2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT27), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n409_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT98), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n443_), .B1(new_n446_), .B2(new_n433_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT100), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n447_), .A2(new_n448_), .A3(new_n440_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n442_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n293_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n451_), .A2(new_n415_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n452_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n413_), .A2(new_n405_), .A3(new_n410_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n453_), .B1(new_n443_), .B2(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n430_), .B1(new_n450_), .B2(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n367_), .B(KEYINPUT30), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(KEYINPUT84), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G71gat), .B(G99gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(G43gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G227gat), .A2(G233gat), .ZN(new_n461_));
  INV_X1    g260(.A(G15gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n460_), .B(new_n463_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n458_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n464_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT84), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n466_), .B1(new_n457_), .B2(new_n467_), .ZN(new_n468_));
  XOR2_X1   g267(.A(new_n276_), .B(KEYINPUT31), .Z(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  OR3_X1    g269(.A1(new_n465_), .A2(new_n468_), .A3(new_n470_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n470_), .B1(new_n465_), .B2(new_n468_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT101), .B1(new_n456_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n473_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n475_), .A2(new_n417_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n454_), .A2(new_n443_), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n476_), .A2(new_n450_), .A3(new_n272_), .A4(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT101), .ZN(new_n479_));
  INV_X1    g278(.A(new_n271_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n417_), .B1(new_n480_), .B2(new_n269_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n477_), .A2(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n482_), .B1(new_n442_), .B2(new_n449_), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n479_), .B(new_n475_), .C1(new_n483_), .C2(new_n430_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n474_), .A2(new_n478_), .A3(new_n484_), .ZN(new_n485_));
  XOR2_X1   g284(.A(G29gat), .B(G36gat), .Z(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT72), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G43gat), .B(G50gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT15), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT8), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G99gat), .A2(G106gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(KEYINPUT6), .ZN(new_n494_));
  OR2_X1    g293(.A1(new_n494_), .A2(KEYINPUT66), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(KEYINPUT66), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT7), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(KEYINPUT65), .ZN(new_n498_));
  NOR2_X1   g297(.A1(G99gat), .A2(G106gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n495_), .A2(new_n496_), .A3(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G85gat), .B(G92gat), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n492_), .B1(new_n501_), .B2(new_n503_), .ZN(new_n504_));
  AOI211_X1 g303(.A(KEYINPUT8), .B(new_n502_), .C1(new_n500_), .C2(new_n494_), .ZN(new_n505_));
  OR2_X1    g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT9), .ZN(new_n507_));
  XNOR2_X1  g306(.A(KEYINPUT10), .B(G99gat), .ZN(new_n508_));
  OAI22_X1  g307(.A1(new_n507_), .A2(new_n502_), .B1(new_n508_), .B2(G106gat), .ZN(new_n509_));
  INV_X1    g308(.A(new_n494_), .ZN(new_n510_));
  INV_X1    g309(.A(G85gat), .ZN(new_n511_));
  INV_X1    g310(.A(G92gat), .ZN(new_n512_));
  NOR3_X1   g311(.A1(new_n511_), .A2(new_n512_), .A3(KEYINPUT9), .ZN(new_n513_));
  NOR3_X1   g312(.A1(new_n509_), .A2(new_n510_), .A3(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT64), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n506_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n491_), .A2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G232gat), .A2(G233gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT35), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n489_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n506_), .A2(new_n524_), .A3(new_n515_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n517_), .A2(new_n523_), .A3(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n521_), .A2(new_n522_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT73), .ZN(new_n529_));
  INV_X1    g328(.A(new_n527_), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n517_), .A2(new_n530_), .A3(new_n523_), .A4(new_n525_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n528_), .A2(new_n529_), .A3(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G190gat), .B(G218gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G134gat), .B(G162gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n532_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT36), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n528_), .A2(new_n535_), .A3(new_n531_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT36), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n532_), .A2(new_n540_), .A3(new_n536_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n538_), .A2(new_n539_), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT103), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n538_), .A2(KEYINPUT103), .A3(new_n539_), .A4(new_n541_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  AND2_X1   g346(.A1(new_n485_), .A2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G57gat), .B(G64gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT67), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT11), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  XOR2_X1   g351(.A(G71gat), .B(G78gat), .Z(new_n553_));
  NOR2_X1   g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  AND2_X1   g353(.A1(new_n552_), .A2(new_n553_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n550_), .A2(new_n551_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n554_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n516_), .A2(new_n557_), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n558_), .A2(KEYINPUT68), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n516_), .A2(new_n557_), .ZN(new_n560_));
  OR2_X1    g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G230gat), .A2(G233gat), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n559_), .A2(new_n560_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n561_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n560_), .A2(KEYINPUT12), .A3(new_n558_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT12), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n516_), .A2(new_n567_), .A3(new_n557_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n566_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(new_n562_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n565_), .A2(new_n570_), .ZN(new_n571_));
  XOR2_X1   g370(.A(G120gat), .B(G148gat), .Z(new_n572_));
  XNOR2_X1  g371(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G176gat), .B(G204gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  XOR2_X1   g375(.A(new_n576_), .B(KEYINPUT70), .Z(new_n577_));
  NAND2_X1  g376(.A1(new_n571_), .A2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n565_), .A2(new_n570_), .A3(new_n576_), .ZN(new_n579_));
  AND3_X1   g378(.A1(new_n578_), .A2(KEYINPUT13), .A3(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(KEYINPUT13), .B1(new_n578_), .B2(new_n579_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  XOR2_X1   g382(.A(G15gat), .B(G22gat), .Z(new_n584_));
  XNOR2_X1  g383(.A(KEYINPUT74), .B(G8gat), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(G1gat), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n584_), .B1(new_n586_), .B2(KEYINPUT14), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT75), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G1gat), .B(G8gat), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT75), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n587_), .B(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n589_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n590_), .A2(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(new_n524_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(G229gat), .A2(G233gat), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n596_), .A2(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n491_), .A2(new_n590_), .A3(new_n594_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n595_), .A2(new_n524_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n600_), .A2(new_n601_), .A3(new_n597_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n599_), .A2(new_n602_), .ZN(new_n603_));
  XOR2_X1   g402(.A(G113gat), .B(G141gat), .Z(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT79), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G169gat), .B(G197gat), .ZN(new_n606_));
  XOR2_X1   g405(.A(new_n605_), .B(new_n606_), .Z(new_n607_));
  OR2_X1    g406(.A1(new_n603_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n603_), .A2(new_n607_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(G231gat), .A2(G233gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n595_), .B(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(new_n557_), .ZN(new_n613_));
  XOR2_X1   g412(.A(G127gat), .B(G155gat), .Z(new_n614_));
  XNOR2_X1  g413(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G183gat), .B(G211gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(KEYINPUT17), .ZN(new_n620_));
  OR2_X1    g419(.A1(new_n619_), .A2(KEYINPUT17), .ZN(new_n621_));
  AND3_X1   g420(.A1(new_n613_), .A2(new_n620_), .A3(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n613_), .A2(new_n620_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NOR3_X1   g424(.A1(new_n583_), .A2(new_n610_), .A3(new_n625_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n548_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(G1gat), .B1(new_n628_), .B2(new_n452_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT37), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n542_), .A2(new_n631_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n538_), .A2(KEYINPUT37), .A3(new_n539_), .A4(new_n541_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n634_), .A2(KEYINPUT77), .A3(new_n624_), .ZN(new_n635_));
  AOI21_X1  g434(.A(KEYINPUT77), .B1(new_n634_), .B2(new_n624_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(new_n582_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT78), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n608_), .A2(new_n609_), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n485_), .A2(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n452_), .A2(G1gat), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n639_), .A2(new_n641_), .A3(new_n642_), .ZN(new_n643_));
  AND3_X1   g442(.A1(new_n643_), .A2(KEYINPUT104), .A3(new_n630_), .ZN(new_n644_));
  AOI21_X1  g443(.A(KEYINPUT104), .B1(new_n643_), .B2(new_n630_), .ZN(new_n645_));
  OAI221_X1 g444(.A(new_n629_), .B1(new_n630_), .B2(new_n643_), .C1(new_n644_), .C2(new_n645_), .ZN(G1324gat));
  NAND2_X1  g445(.A1(new_n450_), .A2(new_n477_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n627_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(G8gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT39), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n639_), .A2(new_n641_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n647_), .ZN(new_n652_));
  OR3_X1    g451(.A1(new_n651_), .A2(new_n585_), .A3(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n650_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT40), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n650_), .A2(new_n653_), .A3(KEYINPUT40), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(G1325gat));
  NAND2_X1  g457(.A1(new_n627_), .A2(new_n473_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(G15gat), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(KEYINPUT105), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT105), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n659_), .A2(new_n662_), .A3(G15gat), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n661_), .A2(KEYINPUT41), .A3(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT41), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n662_), .B1(new_n659_), .B2(G15gat), .ZN(new_n666_));
  AOI211_X1 g465(.A(KEYINPUT105), .B(new_n462_), .C1(new_n627_), .C2(new_n473_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n665_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n639_), .A2(new_n462_), .A3(new_n473_), .A4(new_n641_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n664_), .A2(new_n668_), .A3(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT106), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n664_), .A2(new_n668_), .A3(KEYINPUT106), .A4(new_n669_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1326gat));
  INV_X1    g473(.A(G22gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n675_), .B1(new_n627_), .B2(new_n273_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT42), .Z(new_n677_));
  NAND2_X1  g476(.A1(new_n273_), .A2(new_n675_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n677_), .B1(new_n651_), .B2(new_n678_), .ZN(G1327gat));
  INV_X1    g478(.A(KEYINPUT43), .ZN(new_n680_));
  INV_X1    g479(.A(new_n634_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n484_), .A2(new_n478_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n446_), .A2(new_n433_), .ZN(new_n683_));
  AND4_X1   g482(.A1(new_n448_), .A2(new_n683_), .A3(KEYINPUT27), .A4(new_n440_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n448_), .B1(new_n447_), .B2(new_n440_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n455_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n414_), .A2(new_n429_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(new_n272_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n479_), .B1(new_n689_), .B2(new_n475_), .ZN(new_n690_));
  OAI211_X1 g489(.A(new_n680_), .B(new_n681_), .C1(new_n682_), .C2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(KEYINPUT108), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT108), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n485_), .A2(new_n693_), .A3(new_n680_), .A4(new_n681_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n681_), .B1(new_n682_), .B2(new_n690_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(KEYINPUT43), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n692_), .A2(new_n694_), .A3(new_n696_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n582_), .A2(new_n640_), .A3(new_n625_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT107), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n697_), .A2(KEYINPUT44), .A3(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(KEYINPUT44), .B1(new_n697_), .B2(new_n699_), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n700_), .A2(new_n701_), .A3(new_n452_), .ZN(new_n702_));
  INV_X1    g501(.A(G29gat), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n583_), .A2(new_n624_), .A3(new_n547_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n641_), .A2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n417_), .A2(new_n703_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT109), .ZN(new_n707_));
  OAI22_X1  g506(.A1(new_n702_), .A2(new_n703_), .B1(new_n705_), .B2(new_n707_), .ZN(G1328gat));
  INV_X1    g507(.A(G36gat), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n641_), .A2(new_n709_), .A3(new_n647_), .A4(new_n704_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT45), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n710_), .B(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n700_), .A2(new_n701_), .A3(new_n652_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n713_), .B1(new_n714_), .B2(new_n709_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT110), .ZN(new_n716_));
  AOI21_X1  g515(.A(KEYINPUT46), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n697_), .A2(new_n699_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n697_), .A2(new_n699_), .A3(KEYINPUT44), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n720_), .A2(new_n647_), .A3(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n712_), .B1(new_n722_), .B2(G36gat), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT46), .ZN(new_n724_));
  NOR3_X1   g523(.A1(new_n723_), .A2(KEYINPUT110), .A3(new_n724_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n717_), .A2(new_n725_), .ZN(G1329gat));
  NOR2_X1   g525(.A1(new_n700_), .A2(new_n701_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n727_), .A2(G43gat), .A3(new_n473_), .ZN(new_n728_));
  INV_X1    g527(.A(G43gat), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n729_), .B1(new_n705_), .B2(new_n475_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n731_));
  AND3_X1   g530(.A1(new_n728_), .A2(new_n730_), .A3(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n731_), .B1(new_n728_), .B2(new_n730_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1330gat));
  INV_X1    g533(.A(new_n705_), .ZN(new_n735_));
  AOI21_X1  g534(.A(G50gat), .B1(new_n735_), .B2(new_n273_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n273_), .A2(G50gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n727_), .B2(new_n737_), .ZN(G1331gat));
  NOR2_X1   g537(.A1(new_n582_), .A2(new_n640_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n485_), .A2(new_n739_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n740_), .A2(new_n637_), .ZN(new_n741_));
  INV_X1    g540(.A(G57gat), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n741_), .A2(new_n742_), .A3(new_n417_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n548_), .A2(new_n624_), .A3(new_n739_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT112), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n744_), .B(new_n745_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n746_), .A2(new_n417_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n743_), .B1(new_n747_), .B2(new_n742_), .ZN(G1332gat));
  INV_X1    g547(.A(G64gat), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n741_), .A2(new_n749_), .A3(new_n647_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n746_), .A2(new_n647_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(G64gat), .ZN(new_n752_));
  XOR2_X1   g551(.A(KEYINPUT113), .B(KEYINPUT48), .Z(new_n753_));
  AND2_X1   g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n752_), .A2(new_n753_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n750_), .B1(new_n754_), .B2(new_n755_), .ZN(G1333gat));
  INV_X1    g555(.A(G71gat), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n741_), .A2(new_n757_), .A3(new_n473_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n746_), .A2(new_n473_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(G71gat), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n760_), .A2(KEYINPUT49), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n760_), .A2(KEYINPUT49), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n758_), .B1(new_n761_), .B2(new_n762_), .ZN(G1334gat));
  INV_X1    g562(.A(G78gat), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n741_), .A2(new_n764_), .A3(new_n273_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n746_), .A2(new_n273_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(G78gat), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n767_), .A2(KEYINPUT50), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n767_), .A2(KEYINPUT50), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n765_), .B1(new_n768_), .B2(new_n769_), .ZN(G1335gat));
  AND3_X1   g569(.A1(new_n740_), .A2(new_n625_), .A3(new_n546_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n771_), .A2(new_n511_), .A3(new_n417_), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n582_), .A2(new_n640_), .A3(new_n624_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n697_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT114), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n697_), .A2(KEYINPUT114), .A3(new_n773_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n452_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n772_), .B1(new_n778_), .B2(new_n511_), .ZN(G1336gat));
  NAND3_X1  g578(.A1(new_n771_), .A2(new_n512_), .A3(new_n647_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n652_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n780_), .B1(new_n781_), .B2(new_n512_), .ZN(G1337gat));
  INV_X1    g581(.A(KEYINPUT117), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n475_), .A2(new_n508_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n771_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT115), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT115), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n771_), .A2(new_n787_), .A3(new_n784_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n475_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n790_));
  INV_X1    g589(.A(G99gat), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n783_), .B(new_n789_), .C1(new_n790_), .C2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT116), .ZN(new_n793_));
  NAND2_X1  g592(.A1(KEYINPUT116), .A2(KEYINPUT51), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n789_), .B(new_n794_), .C1(new_n790_), .C2(new_n791_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT51), .ZN(new_n796_));
  AOI22_X1  g595(.A1(new_n793_), .A2(new_n795_), .B1(new_n796_), .B2(new_n792_), .ZN(G1338gat));
  OAI21_X1  g596(.A(G106gat), .B1(new_n774_), .B2(new_n272_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT118), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  OAI211_X1 g599(.A(KEYINPUT118), .B(G106gat), .C1(new_n774_), .C2(new_n272_), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n800_), .A2(KEYINPUT52), .A3(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n798_), .A2(new_n799_), .A3(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(G106gat), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n771_), .A2(new_n805_), .A3(new_n273_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(KEYINPUT53), .B1(new_n802_), .B2(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n800_), .A2(KEYINPUT52), .A3(new_n801_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT53), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n809_), .A2(new_n810_), .A3(new_n804_), .A4(new_n806_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n808_), .A2(new_n811_), .ZN(G1339gat));
  NAND2_X1  g611(.A1(new_n624_), .A2(new_n610_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT119), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n813_), .B(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n582_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT120), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n634_), .B1(new_n816_), .B2(KEYINPUT120), .ZN(new_n819_));
  OAI21_X1  g618(.A(KEYINPUT54), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  OR2_X1    g619(.A1(new_n816_), .A2(KEYINPUT120), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n821_), .A2(new_n822_), .A3(new_n634_), .A4(new_n817_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT56), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n569_), .A2(new_n562_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n563_), .B1(new_n566_), .B2(new_n568_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n827_));
  NOR3_X1   g626(.A1(new_n825_), .A2(new_n826_), .A3(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n577_), .B1(new_n570_), .B2(KEYINPUT55), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n824_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n577_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n831_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n570_), .A2(KEYINPUT55), .ZN(new_n833_));
  OAI211_X1 g632(.A(KEYINPUT56), .B(new_n832_), .C1(new_n833_), .C2(new_n825_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n830_), .A2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n596_), .A2(new_n597_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n600_), .A2(new_n601_), .A3(new_n598_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n836_), .A2(new_n837_), .A3(new_n607_), .ZN(new_n838_));
  AND3_X1   g637(.A1(new_n579_), .A2(new_n608_), .A3(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n835_), .A2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT58), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n835_), .A2(KEYINPUT58), .A3(new_n839_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n842_), .A2(new_n681_), .A3(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT57), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n579_), .A2(new_n640_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n846_), .B1(new_n830_), .B2(new_n834_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n608_), .A2(new_n838_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n848_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n847_), .A2(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n845_), .B1(new_n850_), .B2(new_n546_), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n547_), .B(KEYINPUT57), .C1(new_n849_), .C2(new_n847_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n844_), .A2(new_n851_), .A3(new_n852_), .ZN(new_n853_));
  AOI22_X1  g652(.A1(new_n820_), .A2(new_n823_), .B1(new_n625_), .B2(new_n853_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n647_), .A2(new_n273_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n855_), .A2(new_n473_), .A3(new_n417_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n854_), .A2(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(G113gat), .B1(new_n857_), .B2(new_n640_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n853_), .A2(new_n625_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT121), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n853_), .A2(KEYINPUT121), .A3(new_n625_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n820_), .A2(new_n823_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n856_), .A2(KEYINPUT59), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  OAI21_X1  g666(.A(KEYINPUT59), .B1(new_n854_), .B2(new_n856_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(G113gat), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n871_), .B1(new_n640_), .B2(KEYINPUT122), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n872_), .B1(KEYINPUT122), .B2(new_n871_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n858_), .B1(new_n870_), .B2(new_n873_), .ZN(G1340gat));
  OAI21_X1  g673(.A(G120gat), .B1(new_n869_), .B2(new_n582_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n582_), .A2(KEYINPUT60), .ZN(new_n876_));
  MUX2_X1   g675(.A(new_n876_), .B(KEYINPUT60), .S(G120gat), .Z(new_n877_));
  NAND2_X1  g676(.A1(new_n857_), .A2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n875_), .A2(new_n878_), .ZN(G1341gat));
  OAI21_X1  g678(.A(G127gat), .B1(new_n869_), .B2(new_n625_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n857_), .ZN(new_n881_));
  OR3_X1    g680(.A1(new_n881_), .A2(G127gat), .A3(new_n625_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n882_), .ZN(G1342gat));
  OAI21_X1  g682(.A(G134gat), .B1(new_n869_), .B2(new_n634_), .ZN(new_n884_));
  OR3_X1    g683(.A1(new_n881_), .A2(G134gat), .A3(new_n547_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(G1343gat));
  NAND2_X1  g685(.A1(new_n864_), .A2(new_n859_), .ZN(new_n887_));
  NOR4_X1   g686(.A1(new_n647_), .A2(new_n473_), .A3(new_n272_), .A4(new_n452_), .ZN(new_n888_));
  AND2_X1   g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(new_n640_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n583_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g692(.A1(new_n887_), .A2(new_n888_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n894_), .A2(new_n625_), .ZN(new_n895_));
  XOR2_X1   g694(.A(KEYINPUT61), .B(G155gat), .Z(new_n896_));
  XNOR2_X1  g695(.A(new_n895_), .B(new_n896_), .ZN(G1346gat));
  INV_X1    g696(.A(G162gat), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n898_), .B1(new_n889_), .B2(new_n681_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n546_), .A2(new_n898_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n894_), .A2(new_n900_), .ZN(new_n901_));
  OAI21_X1  g700(.A(KEYINPUT123), .B1(new_n899_), .B2(new_n901_), .ZN(new_n902_));
  OAI21_X1  g701(.A(G162gat), .B1(new_n894_), .B2(new_n634_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT123), .ZN(new_n904_));
  OAI211_X1 g703(.A(new_n903_), .B(new_n904_), .C1(new_n894_), .C2(new_n900_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n902_), .A2(new_n905_), .ZN(G1347gat));
  NAND3_X1  g705(.A1(new_n647_), .A2(new_n272_), .A3(new_n476_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n907_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n908_), .A2(new_n334_), .A3(new_n640_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(KEYINPUT62), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT62), .ZN(new_n911_));
  INV_X1    g710(.A(new_n907_), .ZN(new_n912_));
  NAND4_X1  g711(.A1(new_n865_), .A2(new_n911_), .A3(new_n640_), .A4(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(G169gat), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n910_), .A2(new_n914_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n909_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(G1348gat));
  AOI21_X1  g716(.A(G176gat), .B1(new_n908_), .B2(new_n583_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n854_), .A2(new_n907_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n919_), .A2(G176gat), .A3(new_n583_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT124), .ZN(new_n921_));
  OR2_X1    g720(.A1(new_n920_), .A2(new_n921_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n920_), .A2(new_n921_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n918_), .B1(new_n922_), .B2(new_n923_), .ZN(G1349gat));
  AOI21_X1  g723(.A(G183gat), .B1(new_n919_), .B2(new_n624_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n625_), .A2(new_n371_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n925_), .B1(new_n908_), .B2(new_n926_), .ZN(G1350gat));
  OAI21_X1  g726(.A(new_n546_), .B1(new_n373_), .B2(new_n372_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(KEYINPUT125), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n908_), .A2(new_n929_), .ZN(new_n930_));
  INV_X1    g729(.A(new_n930_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n302_), .B1(new_n908_), .B2(new_n681_), .ZN(new_n932_));
  OAI21_X1  g731(.A(KEYINPUT126), .B1(new_n931_), .B2(new_n932_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n865_), .A2(new_n681_), .A3(new_n912_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(G190gat), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT126), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n935_), .A2(new_n936_), .A3(new_n930_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n933_), .A2(new_n937_), .ZN(G1351gat));
  NOR3_X1   g737(.A1(new_n652_), .A2(new_n473_), .A3(new_n453_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n887_), .A2(new_n939_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n940_), .A2(new_n610_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(new_n231_), .ZN(G1352gat));
  NOR2_X1   g741(.A1(new_n940_), .A2(new_n582_), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n943_), .B(new_n233_), .ZN(G1353gat));
  AND2_X1   g743(.A1(new_n887_), .A2(new_n939_), .ZN(new_n945_));
  AOI211_X1 g744(.A(KEYINPUT63), .B(G211gat), .C1(new_n945_), .C2(new_n624_), .ZN(new_n946_));
  XOR2_X1   g745(.A(KEYINPUT63), .B(G211gat), .Z(new_n947_));
  NAND4_X1  g746(.A1(new_n887_), .A2(new_n624_), .A3(new_n939_), .A4(new_n947_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n948_), .A2(KEYINPUT127), .ZN(new_n949_));
  AND2_X1   g748(.A1(new_n948_), .A2(KEYINPUT127), .ZN(new_n950_));
  NOR3_X1   g749(.A1(new_n946_), .A2(new_n949_), .A3(new_n950_), .ZN(G1354gat));
  NAND3_X1  g750(.A1(new_n945_), .A2(new_n236_), .A3(new_n546_), .ZN(new_n952_));
  OAI21_X1  g751(.A(G218gat), .B1(new_n940_), .B2(new_n634_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n952_), .A2(new_n953_), .ZN(G1355gat));
endmodule


