//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 1 1 1 0 0 1 1 0 0 0 1 0 0 1 0 0 1 0 1 1 1 0 1 1 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n713_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n860_, new_n861_, new_n862_, new_n864_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n890_, new_n891_, new_n893_, new_n894_,
    new_n895_, new_n897_, new_n898_, new_n900_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_;
  XNOR2_X1  g000(.A(KEYINPUT74), .B(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(G8gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G15gat), .B(G22gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G1gat), .B(G8gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G231gat), .A2(G233gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT76), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G57gat), .B(G64gat), .ZN(new_n212_));
  OR2_X1    g011(.A1(new_n212_), .A2(KEYINPUT11), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(KEYINPUT11), .ZN(new_n214_));
  XOR2_X1   g013(.A(G71gat), .B(G78gat), .Z(new_n215_));
  NAND3_X1  g014(.A1(new_n213_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  OR2_X1    g015(.A1(new_n214_), .A2(new_n215_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  XOR2_X1   g017(.A(new_n218_), .B(KEYINPUT75), .Z(new_n219_));
  XNOR2_X1  g018(.A(new_n211_), .B(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G127gat), .B(G155gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n221_), .B(G211gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT16), .B(G183gat), .ZN(new_n223_));
  XOR2_X1   g022(.A(new_n222_), .B(new_n223_), .Z(new_n224_));
  INV_X1    g023(.A(KEYINPUT17), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT77), .ZN(new_n228_));
  OR2_X1    g027(.A1(new_n227_), .A2(KEYINPUT77), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n220_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT78), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n230_), .B(new_n231_), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n224_), .A2(new_n225_), .ZN(new_n233_));
  NOR3_X1   g032(.A1(new_n220_), .A2(new_n226_), .A3(new_n233_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n232_), .A2(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NOR3_X1   g036(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G99gat), .A2(G106gat), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n241_), .A2(KEYINPUT6), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT6), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n243_), .A2(KEYINPUT67), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n240_), .B1(new_n242_), .B2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(KEYINPUT67), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n241_), .A2(KEYINPUT6), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n246_), .A2(new_n247_), .A3(G99gat), .A4(G106gat), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n239_), .A2(new_n245_), .A3(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(G85gat), .ZN(new_n250_));
  INV_X1    g049(.A(G92gat), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(G85gat), .A2(G92gat), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n249_), .A2(KEYINPUT8), .A3(new_n254_), .ZN(new_n255_));
  OR2_X1    g054(.A1(new_n254_), .A2(KEYINPUT8), .ZN(new_n256_));
  NOR3_X1   g055(.A1(new_n237_), .A2(new_n238_), .A3(KEYINPUT8), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n250_), .A2(KEYINPUT65), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT65), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(G85gat), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n258_), .A2(new_n260_), .A3(G92gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n264_), .B1(G85gat), .B2(G92gat), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n263_), .A2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT10), .B(G99gat), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n268_), .A2(G106gat), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n257_), .B1(new_n267_), .B2(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(KEYINPUT66), .B(KEYINPUT6), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(new_n240_), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n255_), .B(new_n256_), .C1(new_n271_), .C2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n218_), .ZN(new_n275_));
  AOI21_X1  g074(.A(KEYINPUT12), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT68), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT9), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT64), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT64), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(KEYINPUT9), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n279_), .A2(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT65), .B(G85gat), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n282_), .B1(G92gat), .B2(new_n283_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n270_), .B1(new_n284_), .B2(new_n265_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n257_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n273_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n255_), .A2(new_n256_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n277_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n265_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n286_), .B1(new_n290_), .B2(new_n269_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n273_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND4_X1  g092(.A1(new_n293_), .A2(KEYINPUT68), .A3(new_n255_), .A4(new_n256_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n289_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n275_), .A2(KEYINPUT12), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n276_), .B1(new_n295_), .B2(new_n297_), .ZN(new_n298_));
  NAND4_X1  g097(.A1(new_n293_), .A2(new_n218_), .A3(new_n255_), .A4(new_n256_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G230gat), .A2(G233gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n298_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n274_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n304_), .A2(new_n218_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n299_), .ZN(new_n306_));
  OAI211_X1 g105(.A(G230gat), .B(G233gat), .C1(new_n305_), .C2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n303_), .A2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G176gat), .B(G204gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G120gat), .B(G148gat), .ZN(new_n312_));
  XOR2_X1   g111(.A(new_n311_), .B(new_n312_), .Z(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT69), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n308_), .B(new_n315_), .ZN(new_n316_));
  OR2_X1    g115(.A1(new_n316_), .A2(KEYINPUT13), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(KEYINPUT13), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G190gat), .B(G218gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G134gat), .B(G162gat), .ZN(new_n322_));
  XOR2_X1   g121(.A(new_n321_), .B(new_n322_), .Z(new_n323_));
  INV_X1    g122(.A(KEYINPUT36), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G232gat), .A2(G233gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT34), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT35), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT72), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n331_), .A2(KEYINPUT72), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT15), .ZN(new_n336_));
  XOR2_X1   g135(.A(G43gat), .B(G50gat), .Z(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT71), .ZN(new_n338_));
  XOR2_X1   g137(.A(G29gat), .B(G36gat), .Z(new_n339_));
  XNOR2_X1  g138(.A(G43gat), .B(G50gat), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT71), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  AND3_X1   g141(.A1(new_n338_), .A2(new_n339_), .A3(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n339_), .B1(new_n338_), .B2(new_n342_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n336_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n338_), .A2(new_n342_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n339_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n338_), .A2(new_n339_), .A3(new_n342_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n348_), .A2(KEYINPUT15), .A3(new_n349_), .ZN(new_n350_));
  AND2_X1   g149(.A1(new_n345_), .A2(new_n350_), .ZN(new_n351_));
  AOI22_X1  g150(.A1(new_n295_), .A2(new_n351_), .B1(new_n330_), .B2(new_n329_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n348_), .A2(new_n349_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n304_), .A2(new_n353_), .ZN(new_n354_));
  AOI211_X1 g153(.A(new_n334_), .B(new_n335_), .C1(new_n352_), .C2(new_n354_), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n352_), .A2(KEYINPUT72), .A3(new_n331_), .A4(new_n354_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n326_), .B1(new_n355_), .B2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT37), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n352_), .A2(new_n354_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n334_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n335_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n360_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n323_), .B(KEYINPUT36), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n363_), .A2(new_n364_), .A3(new_n356_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n358_), .A2(new_n359_), .A3(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n364_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT73), .ZN(new_n368_));
  OR2_X1    g167(.A1(new_n367_), .A2(KEYINPUT73), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n363_), .A2(new_n356_), .A3(new_n368_), .A4(new_n369_), .ZN(new_n370_));
  AND2_X1   g169(.A1(new_n358_), .A2(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n366_), .B1(new_n371_), .B2(new_n359_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n235_), .A2(new_n320_), .A3(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT79), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n208_), .A2(new_n345_), .A3(new_n350_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n207_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n206_), .B(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(new_n353_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G229gat), .A2(G233gat), .ZN(new_n379_));
  XOR2_X1   g178(.A(new_n379_), .B(KEYINPUT80), .Z(new_n380_));
  NAND3_X1  g179(.A1(new_n375_), .A2(new_n378_), .A3(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(KEYINPUT81), .ZN(new_n382_));
  AND2_X1   g181(.A1(new_n377_), .A2(new_n353_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n377_), .A2(new_n353_), .ZN(new_n384_));
  OAI211_X1 g183(.A(G229gat), .B(G233gat), .C1(new_n383_), .C2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT81), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n375_), .A2(new_n378_), .A3(new_n386_), .A4(new_n380_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G113gat), .B(G141gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G169gat), .B(G197gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n382_), .A2(new_n385_), .A3(new_n387_), .A4(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT82), .ZN(new_n393_));
  OR2_X1    g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n392_), .A2(new_n393_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n382_), .A2(new_n385_), .A3(new_n387_), .ZN(new_n396_));
  AOI22_X1  g195(.A1(new_n394_), .A2(new_n395_), .B1(new_n396_), .B2(new_n390_), .ZN(new_n397_));
  OR4_X1    g196(.A1(KEYINPUT92), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT2), .ZN(new_n399_));
  INV_X1    g198(.A(G141gat), .ZN(new_n400_));
  INV_X1    g199(.A(G148gat), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n399_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n403_));
  OAI22_X1  g202(.A1(KEYINPUT92), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n398_), .A2(new_n402_), .A3(new_n403_), .A4(new_n404_), .ZN(new_n405_));
  AND2_X1   g204(.A1(G155gat), .A2(G162gat), .ZN(new_n406_));
  NOR2_X1   g205(.A1(G155gat), .A2(G162gat), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n405_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT1), .ZN(new_n410_));
  AOI22_X1  g209(.A1(new_n408_), .A2(new_n410_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n411_));
  AOI22_X1  g210(.A1(new_n406_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n409_), .A2(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(G50gat), .B1(new_n414_), .B2(KEYINPUT29), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(KEYINPUT28), .B(G22gat), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NOR3_X1   g217(.A1(new_n414_), .A2(KEYINPUT29), .A3(G50gat), .ZN(new_n419_));
  OR3_X1    g218(.A1(new_n416_), .A2(new_n418_), .A3(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n418_), .B1(new_n416_), .B2(new_n419_), .ZN(new_n421_));
  XOR2_X1   g220(.A(G197gat), .B(G204gat), .Z(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT21), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G211gat), .B(G218gat), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n425_), .A2(KEYINPUT93), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT93), .ZN(new_n427_));
  NOR3_X1   g226(.A1(new_n423_), .A2(new_n427_), .A3(new_n424_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n422_), .A2(KEYINPUT21), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n423_), .A2(new_n424_), .ZN(new_n430_));
  OAI22_X1  g229(.A1(new_n426_), .A2(new_n428_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n414_), .A2(KEYINPUT29), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n433_), .A2(G228gat), .A3(G233gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G228gat), .A2(G233gat), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n431_), .A2(new_n435_), .A3(new_n432_), .ZN(new_n436_));
  XOR2_X1   g235(.A(G78gat), .B(G106gat), .Z(new_n437_));
  NAND3_X1  g236(.A1(new_n434_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n437_), .B1(new_n434_), .B2(new_n436_), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n420_), .B(new_n421_), .C1(new_n439_), .C2(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(KEYINPUT94), .B1(new_n421_), .B2(new_n420_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n440_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(new_n438_), .A3(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n440_), .A2(KEYINPUT94), .ZN(new_n445_));
  AND3_X1   g244(.A1(new_n441_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT23), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n447_), .A2(G183gat), .A3(G190gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(KEYINPUT84), .ZN(new_n449_));
  INV_X1    g248(.A(G183gat), .ZN(new_n450_));
  INV_X1    g249(.A(G190gat), .ZN(new_n451_));
  OAI21_X1  g250(.A(KEYINPUT23), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n449_), .A2(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n453_), .B1(G183gat), .B2(G190gat), .ZN(new_n454_));
  XOR2_X1   g253(.A(KEYINPUT86), .B(G176gat), .Z(new_n455_));
  XNOR2_X1  g254(.A(KEYINPUT22), .B(G169gat), .ZN(new_n456_));
  AOI22_X1  g255(.A1(new_n455_), .A2(new_n456_), .B1(G169gat), .B2(G176gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n454_), .A2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(KEYINPUT26), .B(G190gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(KEYINPUT25), .B(G183gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  OR2_X1    g260(.A1(G169gat), .A2(G176gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G169gat), .A2(G176gat), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n462_), .A2(KEYINPUT24), .A3(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n461_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT95), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n452_), .A2(new_n448_), .ZN(new_n468_));
  OR2_X1    g267(.A1(new_n462_), .A2(KEYINPUT24), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n461_), .A2(KEYINPUT95), .A3(new_n464_), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n467_), .A2(new_n468_), .A3(new_n469_), .A4(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n458_), .A2(new_n471_), .ZN(new_n472_));
  OAI21_X1  g271(.A(KEYINPUT20), .B1(new_n472_), .B2(new_n431_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G226gat), .A2(G233gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT19), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n473_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n453_), .A2(new_n469_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT85), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT83), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n480_), .B1(new_n451_), .B2(KEYINPUT26), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n481_), .B(new_n460_), .C1(new_n459_), .C2(new_n480_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n453_), .A2(KEYINPUT85), .A3(new_n469_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n479_), .A2(new_n482_), .A3(new_n483_), .A4(new_n464_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n468_), .B1(G183gat), .B2(G190gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n457_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n484_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT96), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n487_), .A2(new_n488_), .A3(new_n431_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n488_), .B1(new_n487_), .B2(new_n431_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n476_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n472_), .A2(new_n431_), .ZN(new_n492_));
  OAI211_X1 g291(.A(new_n492_), .B(KEYINPUT20), .C1(new_n487_), .C2(new_n431_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(new_n475_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n491_), .A2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G64gat), .B(G92gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G8gat), .B(G36gat), .ZN(new_n499_));
  XOR2_X1   g298(.A(new_n498_), .B(new_n499_), .Z(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(KEYINPUT98), .B1(new_n495_), .B2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT98), .ZN(new_n503_));
  AOI211_X1 g302(.A(new_n503_), .B(new_n500_), .C1(new_n491_), .C2(new_n494_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n491_), .A2(new_n494_), .A3(new_n500_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NOR3_X1   g305(.A1(new_n502_), .A2(new_n504_), .A3(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G1gat), .B(G29gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(new_n250_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(KEYINPUT0), .B(G57gat), .ZN(new_n510_));
  XOR2_X1   g309(.A(new_n509_), .B(new_n510_), .Z(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G127gat), .B(G134gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G113gat), .B(G120gat), .ZN(new_n514_));
  OR2_X1    g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT90), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n513_), .A2(new_n514_), .ZN(new_n517_));
  XOR2_X1   g316(.A(new_n517_), .B(KEYINPUT89), .Z(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT91), .B1(new_n516_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT90), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n515_), .B(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT91), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n517_), .B(KEYINPUT89), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n521_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n519_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(new_n414_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT4), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n515_), .A2(new_n517_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT100), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n530_), .A2(new_n414_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT99), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n526_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n525_), .A2(KEYINPUT99), .A3(new_n414_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n531_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n528_), .B1(new_n535_), .B2(new_n527_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G225gat), .A2(G233gat), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n512_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n531_), .ZN(new_n539_));
  AND3_X1   g338(.A1(new_n525_), .A2(KEYINPUT99), .A3(new_n414_), .ZN(new_n540_));
  AOI21_X1  g339(.A(KEYINPUT99), .B1(new_n525_), .B2(new_n414_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n539_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n538_), .B1(new_n537_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n537_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n536_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n535_), .A2(new_n537_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT33), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(KEYINPUT101), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n545_), .A2(new_n512_), .A3(new_n546_), .A4(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n528_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n550_), .B1(new_n542_), .B2(KEYINPUT4), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n512_), .B(new_n546_), .C1(new_n551_), .C2(new_n537_), .ZN(new_n552_));
  XOR2_X1   g351(.A(KEYINPUT101), .B(KEYINPUT33), .Z(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n507_), .A2(new_n543_), .A3(new_n549_), .A4(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n475_), .ZN(new_n556_));
  OR2_X1    g355(.A1(new_n489_), .A2(new_n490_), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n473_), .B(KEYINPUT102), .Z(new_n558_));
  AOI21_X1  g357(.A(new_n556_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n493_), .A2(new_n475_), .ZN(new_n560_));
  OAI211_X1 g359(.A(KEYINPUT32), .B(new_n500_), .C1(new_n559_), .C2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n500_), .A2(KEYINPUT32), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n491_), .A2(new_n494_), .A3(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n512_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n552_), .ZN(new_n565_));
  OAI211_X1 g364(.A(new_n561_), .B(new_n563_), .C1(new_n564_), .C2(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n446_), .B1(new_n555_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT88), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT30), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n484_), .A2(new_n569_), .A3(new_n486_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n569_), .B1(new_n484_), .B2(new_n486_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n568_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n572_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n574_), .A2(KEYINPUT88), .A3(new_n570_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G15gat), .B(G43gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G71gat), .B(G99gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G227gat), .A2(G233gat), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n579_), .B(KEYINPUT87), .Z(new_n580_));
  XOR2_X1   g379(.A(new_n578_), .B(new_n580_), .Z(new_n581_));
  NAND3_X1  g380(.A1(new_n573_), .A2(new_n575_), .A3(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n581_), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n574_), .A2(KEYINPUT88), .A3(new_n570_), .A4(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n525_), .B(KEYINPUT31), .Z(new_n585_));
  NAND3_X1  g384(.A1(new_n582_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n585_), .B1(new_n582_), .B2(new_n584_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n495_), .A2(new_n501_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(new_n503_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n495_), .A2(KEYINPUT98), .A3(new_n501_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n591_), .A2(new_n505_), .A3(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT27), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n582_), .A2(new_n584_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n585_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n446_), .A2(new_n598_), .A3(new_n586_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n441_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n600_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n501_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n603_), .A2(KEYINPUT27), .A3(new_n505_), .ZN(new_n604_));
  AND3_X1   g403(.A1(new_n595_), .A2(new_n602_), .A3(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n564_), .A2(new_n565_), .ZN(new_n606_));
  AOI22_X1  g405(.A1(new_n567_), .A2(new_n589_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  NOR3_X1   g406(.A1(new_n374_), .A2(new_n397_), .A3(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n606_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n608_), .A2(new_n609_), .A3(new_n202_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT38), .ZN(new_n611_));
  INV_X1    g410(.A(new_n607_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n319_), .A2(new_n397_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n235_), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n363_), .A2(new_n364_), .A3(new_n356_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n325_), .B1(new_n363_), .B2(new_n356_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n614_), .A2(new_n617_), .ZN(new_n618_));
  AND3_X1   g417(.A1(new_n612_), .A2(new_n613_), .A3(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  OAI21_X1  g419(.A(G1gat), .B1(new_n620_), .B2(new_n606_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n611_), .A2(new_n621_), .ZN(G1324gat));
  AND2_X1   g421(.A1(new_n595_), .A2(new_n604_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n203_), .B1(new_n619_), .B2(new_n624_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT39), .Z(new_n626_));
  NAND3_X1  g425(.A1(new_n608_), .A2(new_n203_), .A3(new_n624_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT40), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n628_), .B(new_n629_), .ZN(G1325gat));
  INV_X1    g429(.A(G15gat), .ZN(new_n631_));
  INV_X1    g430(.A(new_n589_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n631_), .B1(new_n619_), .B2(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT41), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n608_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(G1326gat));
  INV_X1    g435(.A(G22gat), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n637_), .B1(new_n619_), .B2(new_n446_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n638_), .B(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n608_), .A2(new_n637_), .A3(new_n446_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(G1327gat));
  OR2_X1    g441(.A1(KEYINPUT104), .A2(KEYINPUT43), .ZN(new_n643_));
  NAND2_X1  g442(.A1(KEYINPUT104), .A2(KEYINPUT43), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n615_), .A2(new_n616_), .A3(KEYINPUT37), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n359_), .B1(new_n358_), .B2(new_n370_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT105), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n643_), .B(new_n644_), .C1(new_n607_), .C2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT43), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n605_), .A2(new_n606_), .ZN(new_n651_));
  AOI211_X1 g450(.A(new_n632_), .B(new_n446_), .C1(new_n555_), .C2(new_n566_), .ZN(new_n652_));
  OAI211_X1 g451(.A(new_n650_), .B(new_n647_), .C1(new_n651_), .C2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n649_), .A2(new_n653_), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n235_), .A2(new_n397_), .A3(new_n319_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT44), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n656_), .A2(KEYINPUT106), .A3(new_n657_), .ZN(new_n658_));
  XOR2_X1   g457(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n659_));
  OAI21_X1  g458(.A(new_n658_), .B1(new_n656_), .B2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT107), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n660_), .A2(new_n661_), .A3(new_n609_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n656_), .A2(new_n659_), .ZN(new_n663_));
  AND4_X1   g462(.A1(KEYINPUT106), .A2(new_n654_), .A3(new_n657_), .A4(new_n655_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n609_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(KEYINPUT107), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n662_), .A2(new_n666_), .A3(G29gat), .ZN(new_n667_));
  INV_X1    g466(.A(new_n617_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n607_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(new_n655_), .ZN(new_n670_));
  OR2_X1    g469(.A1(new_n606_), .A2(G29gat), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n667_), .B1(new_n670_), .B2(new_n671_), .ZN(G1328gat));
  NOR2_X1   g471(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n673_));
  INV_X1    g472(.A(G36gat), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n674_), .B1(new_n660_), .B2(new_n624_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n670_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n676_), .A2(new_n674_), .A3(new_n624_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT45), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n673_), .B1(new_n675_), .B2(new_n679_), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n656_), .A2(new_n659_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n623_), .B1(new_n681_), .B2(new_n658_), .ZN(new_n682_));
  OAI221_X1 g481(.A(new_n678_), .B1(KEYINPUT108), .B2(KEYINPUT46), .C1(new_n682_), .C2(new_n674_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n680_), .A2(new_n683_), .ZN(G1329gat));
  INV_X1    g483(.A(KEYINPUT47), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n632_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(G43gat), .ZN(new_n687_));
  NOR3_X1   g486(.A1(new_n670_), .A2(G43gat), .A3(new_n589_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n685_), .B1(new_n687_), .B2(new_n689_), .ZN(new_n690_));
  AOI211_X1 g489(.A(KEYINPUT47), .B(new_n688_), .C1(new_n686_), .C2(G43gat), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1330gat));
  NAND3_X1  g491(.A1(new_n660_), .A2(KEYINPUT109), .A3(new_n446_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n446_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT109), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n693_), .A2(new_n696_), .A3(G50gat), .ZN(new_n697_));
  OR3_X1    g496(.A1(new_n670_), .A2(G50gat), .A3(new_n600_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(G1331gat));
  XNOR2_X1  g498(.A(new_n392_), .B(new_n393_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n396_), .A2(new_n390_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n607_), .A2(new_n702_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n614_), .A2(new_n320_), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n703_), .A2(new_n372_), .A3(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(G57gat), .B1(new_n705_), .B2(new_n609_), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n703_), .A2(new_n668_), .A3(new_n704_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n609_), .A2(G57gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n706_), .B1(new_n707_), .B2(new_n708_), .ZN(G1332gat));
  INV_X1    g508(.A(G64gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n710_), .B1(new_n707_), .B2(new_n624_), .ZN(new_n711_));
  XOR2_X1   g510(.A(new_n711_), .B(KEYINPUT48), .Z(new_n712_));
  NAND3_X1  g511(.A1(new_n705_), .A2(new_n710_), .A3(new_n624_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1333gat));
  INV_X1    g513(.A(G71gat), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n705_), .A2(new_n715_), .A3(new_n632_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n715_), .B1(new_n707_), .B2(new_n632_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(KEYINPUT110), .B(KEYINPUT49), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n717_), .A2(new_n718_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n716_), .B1(new_n719_), .B2(new_n720_), .ZN(G1334gat));
  INV_X1    g520(.A(G78gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n722_), .B1(new_n707_), .B2(new_n446_), .ZN(new_n723_));
  XOR2_X1   g522(.A(new_n723_), .B(KEYINPUT50), .Z(new_n724_));
  NAND3_X1  g523(.A1(new_n705_), .A2(new_n722_), .A3(new_n446_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(G1335gat));
  NAND3_X1  g525(.A1(new_n614_), .A2(new_n397_), .A3(new_n319_), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n727_), .A2(new_n607_), .A3(new_n668_), .ZN(new_n728_));
  AOI21_X1  g527(.A(G85gat), .B1(new_n728_), .B2(new_n609_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n727_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n654_), .A2(new_n730_), .ZN(new_n731_));
  OR2_X1    g530(.A1(new_n731_), .A2(KEYINPUT111), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(KEYINPUT111), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n609_), .A2(new_n283_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n729_), .B1(new_n734_), .B2(new_n735_), .ZN(G1336gat));
  NAND3_X1  g535(.A1(new_n728_), .A2(new_n251_), .A3(new_n624_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n623_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n737_), .B1(new_n738_), .B2(new_n251_), .ZN(G1337gat));
  OAI21_X1  g538(.A(G99gat), .B1(new_n731_), .B2(new_n589_), .ZN(new_n740_));
  AOI21_X1  g539(.A(KEYINPUT113), .B1(KEYINPUT112), .B2(KEYINPUT51), .ZN(new_n741_));
  INV_X1    g540(.A(new_n268_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n728_), .A2(new_n742_), .A3(new_n632_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n740_), .A2(new_n741_), .A3(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n740_), .A2(new_n743_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(KEYINPUT113), .B2(KEYINPUT51), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n744_), .B1(new_n746_), .B2(new_n741_), .ZN(G1338gat));
  INV_X1    g546(.A(G106gat), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n728_), .A2(new_n748_), .A3(new_n446_), .ZN(new_n749_));
  AOI211_X1 g548(.A(new_n600_), .B(new_n727_), .C1(new_n649_), .C2(new_n653_), .ZN(new_n750_));
  OAI21_X1  g549(.A(KEYINPUT114), .B1(new_n750_), .B2(new_n748_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT114), .ZN(new_n752_));
  OAI211_X1 g551(.A(new_n752_), .B(G106gat), .C1(new_n731_), .C2(new_n600_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT52), .ZN(new_n754_));
  AND3_X1   g553(.A1(new_n751_), .A2(new_n753_), .A3(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n751_), .B2(new_n753_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n749_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(KEYINPUT53), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT53), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n759_), .B(new_n749_), .C1(new_n755_), .C2(new_n756_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(G1339gat));
  NOR2_X1   g560(.A1(new_n624_), .A2(new_n606_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n601_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT117), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT56), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n300_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n767_));
  AOI21_X1  g566(.A(KEYINPUT55), .B1(new_n298_), .B2(new_n302_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n296_), .B1(new_n289_), .B2(new_n294_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT55), .ZN(new_n770_));
  NOR4_X1   g569(.A1(new_n769_), .A2(new_n276_), .A3(new_n301_), .A4(new_n770_), .ZN(new_n771_));
  NOR3_X1   g570(.A1(new_n767_), .A2(new_n768_), .A3(new_n771_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n766_), .B1(new_n772_), .B2(new_n313_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n303_), .A2(new_n770_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n771_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  OAI211_X1 g575(.A(KEYINPUT56), .B(new_n314_), .C1(new_n776_), .C2(new_n767_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n773_), .A2(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n380_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n375_), .A2(new_n378_), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n779_), .B(new_n390_), .C1(new_n780_), .C2(new_n380_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n303_), .A2(new_n307_), .A3(new_n313_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n700_), .A2(new_n781_), .A3(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(KEYINPUT58), .B1(new_n778_), .B2(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n765_), .B1(new_n785_), .B2(new_n372_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n783_), .B1(new_n773_), .B2(new_n777_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(KEYINPUT58), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n647_), .B(KEYINPUT117), .C1(new_n787_), .C2(KEYINPUT58), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n786_), .A2(new_n788_), .A3(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT118), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT118), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n786_), .A2(new_n789_), .A3(new_n792_), .A4(new_n788_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n791_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n782_), .ZN(new_n795_));
  OAI21_X1  g594(.A(KEYINPUT115), .B1(new_n397_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n702_), .A2(new_n797_), .A3(new_n782_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n796_), .A2(new_n798_), .A3(new_n778_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n700_), .A2(new_n781_), .ZN(new_n800_));
  OR2_X1    g599(.A1(new_n800_), .A2(new_n316_), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n799_), .A2(new_n801_), .ZN(new_n802_));
  OAI211_X1 g601(.A(KEYINPUT116), .B(KEYINPUT57), .C1(new_n802_), .C2(new_n617_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT57), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n617_), .B1(new_n799_), .B2(new_n801_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT116), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n804_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n803_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n794_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT119), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n794_), .A2(KEYINPUT119), .A3(new_n808_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n811_), .A2(new_n614_), .A3(new_n812_), .ZN(new_n813_));
  OR3_X1    g612(.A1(new_n373_), .A2(KEYINPUT54), .A3(new_n702_), .ZN(new_n814_));
  OAI21_X1  g613(.A(KEYINPUT54), .B1(new_n373_), .B2(new_n702_), .ZN(new_n815_));
  AND2_X1   g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n764_), .B1(new_n813_), .B2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(G113gat), .B1(new_n818_), .B2(new_n702_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n818_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n235_), .B1(new_n808_), .B2(new_n790_), .ZN(new_n821_));
  OR2_X1    g620(.A1(new_n816_), .A2(new_n821_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n764_), .A2(KEYINPUT59), .ZN(new_n823_));
  AOI22_X1  g622(.A1(new_n820_), .A2(KEYINPUT59), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n702_), .A2(G113gat), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n825_), .B(KEYINPUT120), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n819_), .B1(new_n824_), .B2(new_n826_), .ZN(G1340gat));
  NAND2_X1  g626(.A1(new_n822_), .A2(new_n823_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT59), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n319_), .B(new_n828_), .C1(new_n818_), .C2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT60), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n831_), .B1(new_n320_), .B2(G120gat), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n818_), .A2(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(G120gat), .B1(new_n830_), .B2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n831_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(G1341gat));
  INV_X1    g635(.A(G127gat), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n614_), .A2(new_n837_), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n828_), .B(new_n838_), .C1(new_n818_), .C2(new_n829_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n764_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n816_), .A2(new_n235_), .A3(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n837_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n839_), .A2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(KEYINPUT121), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT121), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n839_), .A2(new_n845_), .A3(new_n842_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n846_), .ZN(G1342gat));
  NAND2_X1  g646(.A1(new_n813_), .A2(new_n817_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n848_), .A2(new_n617_), .A3(new_n840_), .ZN(new_n849_));
  INV_X1    g648(.A(G134gat), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  XOR2_X1   g650(.A(KEYINPUT122), .B(G134gat), .Z(new_n852_));
  NOR2_X1   g651(.A1(new_n372_), .A2(new_n852_), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n828_), .B(new_n853_), .C1(new_n818_), .C2(new_n829_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n851_), .A2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT123), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n851_), .A2(new_n854_), .A3(KEYINPUT123), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(G1343gat));
  INV_X1    g658(.A(new_n599_), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n848_), .A2(new_n860_), .A3(new_n762_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n702_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n319_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g664(.A1(new_n861_), .A2(new_n235_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(KEYINPUT61), .B(G155gat), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n866_), .B(new_n867_), .ZN(G1346gat));
  AOI21_X1  g667(.A(G162gat), .B1(new_n861_), .B2(new_n617_), .ZN(new_n869_));
  INV_X1    g668(.A(G162gat), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n648_), .A2(new_n870_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(KEYINPUT124), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n869_), .B1(new_n861_), .B2(new_n872_), .ZN(G1347gat));
  NOR2_X1   g672(.A1(new_n623_), .A2(new_n609_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n875_), .A2(new_n601_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n822_), .A2(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(G169gat), .B1(new_n877_), .B2(new_n397_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT62), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n877_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n881_), .A2(new_n702_), .A3(new_n456_), .ZN(new_n882_));
  AND2_X1   g681(.A1(new_n882_), .A2(new_n878_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n880_), .B1(new_n883_), .B2(new_n879_), .ZN(G1348gat));
  OAI21_X1  g683(.A(new_n455_), .B1(new_n877_), .B2(new_n320_), .ZN(new_n885_));
  NAND4_X1  g684(.A1(new_n848_), .A2(G176gat), .A3(new_n319_), .A4(new_n876_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT125), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n887_), .B(new_n888_), .ZN(G1349gat));
  NOR2_X1   g688(.A1(new_n614_), .A2(new_n460_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n816_), .A2(new_n235_), .A3(new_n876_), .ZN(new_n891_));
  AOI22_X1  g690(.A1(new_n881_), .A2(new_n890_), .B1(new_n450_), .B2(new_n891_), .ZN(G1350gat));
  NAND3_X1  g691(.A1(new_n881_), .A2(new_n459_), .A3(new_n617_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n881_), .A2(new_n647_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n893_), .B1(new_n895_), .B2(new_n451_), .ZN(G1351gat));
  AOI211_X1 g695(.A(new_n599_), .B(new_n875_), .C1(new_n813_), .C2(new_n817_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n702_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g698(.A1(new_n897_), .A2(new_n319_), .ZN(new_n900_));
  INV_X1    g699(.A(G204gat), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n901_), .A2(KEYINPUT126), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n900_), .B(new_n902_), .ZN(G1353gat));
  NOR2_X1   g702(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n904_), .B1(new_n897_), .B2(new_n235_), .ZN(new_n905_));
  AND3_X1   g704(.A1(new_n794_), .A2(KEYINPUT119), .A3(new_n808_), .ZN(new_n906_));
  AOI21_X1  g705(.A(KEYINPUT119), .B1(new_n794_), .B2(new_n808_), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n906_), .A2(new_n907_), .A3(new_n235_), .ZN(new_n908_));
  OAI211_X1 g707(.A(new_n860_), .B(new_n874_), .C1(new_n908_), .C2(new_n816_), .ZN(new_n909_));
  XOR2_X1   g708(.A(KEYINPUT63), .B(G211gat), .Z(new_n910_));
  NOR3_X1   g709(.A1(new_n909_), .A2(new_n614_), .A3(new_n910_), .ZN(new_n911_));
  OAI21_X1  g710(.A(KEYINPUT127), .B1(new_n905_), .B2(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n910_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n897_), .A2(new_n235_), .A3(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT127), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n909_), .A2(new_n614_), .ZN(new_n916_));
  OAI211_X1 g715(.A(new_n914_), .B(new_n915_), .C1(new_n916_), .C2(new_n904_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n912_), .A2(new_n917_), .ZN(G1354gat));
  AND3_X1   g717(.A1(new_n897_), .A2(G218gat), .A3(new_n647_), .ZN(new_n919_));
  AOI21_X1  g718(.A(G218gat), .B1(new_n897_), .B2(new_n617_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n919_), .A2(new_n920_), .ZN(G1355gat));
endmodule


