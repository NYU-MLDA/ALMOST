//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 0 1 0 1 0 1 0 0 1 1 0 0 0 1 0 1 1 0 1 1 0 1 0 0 1 0 0 0 0 0 1 1 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 1 0 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n795_, new_n796_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n902_, new_n903_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n910_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n947_, new_n948_, new_n949_, new_n951_, new_n952_, new_n953_,
    new_n955_, new_n956_, new_n958_, new_n959_, new_n960_, new_n962_,
    new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_,
    new_n969_, new_n970_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n977_, new_n978_, new_n979_;
  INV_X1    g000(.A(KEYINPUT100), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G1gat), .B(G29gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(G85gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT0), .B(G57gat), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  INV_X1    g005(.A(KEYINPUT33), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT98), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G225gat), .A2(G233gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210_));
  INV_X1    g009(.A(G141gat), .ZN(new_n211_));
  INV_X1    g010(.A(G148gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT87), .B1(new_n214_), .B2(KEYINPUT1), .ZN(new_n215_));
  OR2_X1    g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(KEYINPUT1), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  NOR3_X1   g017(.A1(new_n214_), .A2(KEYINPUT87), .A3(KEYINPUT1), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n210_), .B(new_n213_), .C1(new_n218_), .C2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT3), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT2), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n210_), .A2(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n222_), .A2(new_n224_), .A3(new_n225_), .A4(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT88), .ZN(new_n228_));
  AND2_X1   g027(.A1(new_n216_), .A2(new_n214_), .ZN(new_n229_));
  AND3_X1   g028(.A1(new_n227_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n228_), .B1(new_n227_), .B2(new_n229_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n220_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT97), .ZN(new_n233_));
  XOR2_X1   g032(.A(G127gat), .B(G134gat), .Z(new_n234_));
  XOR2_X1   g033(.A(G113gat), .B(G120gat), .Z(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n232_), .A2(new_n233_), .A3(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n227_), .A2(new_n229_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(KEYINPUT88), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n227_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n242_), .A2(new_n220_), .A3(new_n236_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n238_), .A2(KEYINPUT4), .A3(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT4), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n232_), .A2(new_n237_), .A3(new_n233_), .A4(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n209_), .B1(new_n244_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n209_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n232_), .A2(new_n237_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n248_), .B1(new_n249_), .B2(new_n243_), .ZN(new_n250_));
  OAI211_X1 g049(.A(new_n206_), .B(new_n208_), .C1(new_n247_), .C2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT99), .ZN(new_n252_));
  AOI21_X1  g051(.A(KEYINPUT98), .B1(new_n252_), .B2(new_n207_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n251_), .A2(new_n254_), .ZN(new_n255_));
  XOR2_X1   g054(.A(G8gat), .B(G36gat), .Z(new_n256_));
  XNOR2_X1  g055(.A(G64gat), .B(G92gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G226gat), .A2(G233gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT19), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT20), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT91), .ZN(new_n265_));
  INV_X1    g064(.A(G204gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(KEYINPUT91), .A2(G204gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT90), .B(G197gat), .ZN(new_n271_));
  AOI22_X1  g070(.A1(new_n270_), .A2(G197gat), .B1(new_n271_), .B2(G204gat), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT21), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G211gat), .B(G218gat), .ZN(new_n274_));
  OR3_X1    g073(.A1(new_n272_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n274_), .ZN(new_n276_));
  INV_X1    g075(.A(G197gat), .ZN(new_n277_));
  AND2_X1   g076(.A1(KEYINPUT91), .A2(G204gat), .ZN(new_n278_));
  NOR2_X1   g077(.A1(KEYINPUT91), .A2(G204gat), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n277_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n280_), .B1(new_n271_), .B2(G204gat), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n276_), .B1(new_n281_), .B2(KEYINPUT21), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n277_), .A2(KEYINPUT90), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT90), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(G197gat), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n283_), .A2(new_n285_), .A3(G204gat), .ZN(new_n286_));
  OAI211_X1 g085(.A(new_n286_), .B(new_n273_), .C1(new_n269_), .C2(new_n277_), .ZN(new_n287_));
  AOI21_X1  g086(.A(KEYINPUT92), .B1(new_n282_), .B2(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(G204gat), .B1(new_n283_), .B2(new_n285_), .ZN(new_n289_));
  AOI21_X1  g088(.A(G197gat), .B1(new_n267_), .B2(new_n268_), .ZN(new_n290_));
  OAI21_X1  g089(.A(KEYINPUT21), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  AND4_X1   g090(.A1(KEYINPUT92), .A2(new_n291_), .A3(new_n287_), .A4(new_n274_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n275_), .B1(new_n288_), .B2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT95), .B(KEYINPUT24), .ZN(new_n294_));
  NOR2_X1   g093(.A1(G169gat), .A2(G176gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n295_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G169gat), .A2(G176gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n296_), .B1(new_n299_), .B2(new_n294_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT25), .B(G183gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT26), .B(G190gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G183gat), .A2(G190gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT23), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT23), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n306_), .A2(G183gat), .A3(G190gat), .ZN(new_n307_));
  AOI22_X1  g106(.A1(new_n302_), .A2(new_n303_), .B1(new_n305_), .B2(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(G183gat), .A2(G190gat), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n309_), .B1(new_n306_), .B2(new_n304_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n310_), .B1(new_n306_), .B2(new_n304_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n298_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT22), .B(G169gat), .ZN(new_n313_));
  INV_X1    g112(.A(G176gat), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n312_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  AOI22_X1  g114(.A1(new_n301_), .A2(new_n308_), .B1(new_n311_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n264_), .B1(new_n293_), .B2(new_n317_), .ZN(new_n318_));
  NOR3_X1   g117(.A1(new_n272_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n291_), .A2(new_n287_), .A3(new_n274_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT92), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n291_), .A2(new_n287_), .A3(KEYINPUT92), .A4(new_n274_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n319_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(G183gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(KEYINPUT25), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT25), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(G183gat), .ZN(new_n328_));
  INV_X1    g127(.A(G190gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT26), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT26), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(G190gat), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n326_), .A2(new_n328_), .A3(new_n330_), .A4(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT82), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n297_), .A2(KEYINPUT24), .A3(new_n298_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT24), .ZN(new_n336_));
  AOI22_X1  g135(.A1(new_n305_), .A2(new_n307_), .B1(new_n336_), .B2(new_n295_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT82), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n302_), .A2(new_n303_), .A3(new_n338_), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n334_), .A2(new_n335_), .A3(new_n337_), .A4(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT83), .ZN(new_n341_));
  INV_X1    g140(.A(G169gat), .ZN(new_n342_));
  OAI21_X1  g141(.A(KEYINPUT22), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  OR2_X1    g142(.A1(new_n342_), .A2(KEYINPUT22), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n314_), .B(new_n343_), .C1(new_n344_), .C2(new_n341_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n311_), .A2(new_n345_), .A3(new_n298_), .ZN(new_n346_));
  AND2_X1   g145(.A1(new_n340_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n324_), .A2(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n263_), .B1(new_n318_), .B2(new_n348_), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n275_), .B(new_n316_), .C1(new_n288_), .C2(new_n292_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT20), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n322_), .A2(new_n323_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n347_), .B1(new_n352_), .B2(new_n275_), .ZN(new_n353_));
  NOR3_X1   g152(.A1(new_n351_), .A2(new_n353_), .A3(new_n262_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n260_), .B1(new_n349_), .B2(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(KEYINPUT20), .B1(new_n324_), .B2(new_n316_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n340_), .A2(new_n346_), .ZN(new_n357_));
  AOI211_X1 g156(.A(new_n319_), .B(new_n357_), .C1(new_n322_), .C2(new_n323_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n262_), .B1(new_n356_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n260_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n264_), .B1(new_n324_), .B2(new_n316_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n293_), .A2(new_n357_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n361_), .A2(new_n263_), .A3(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n359_), .A2(new_n360_), .A3(new_n363_), .ZN(new_n364_));
  AND3_X1   g163(.A1(new_n255_), .A2(new_n355_), .A3(new_n364_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n206_), .B1(new_n247_), .B2(new_n250_), .ZN(new_n366_));
  AND2_X1   g165(.A1(new_n249_), .A2(new_n243_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n206_), .B1(new_n367_), .B2(new_n248_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n244_), .A2(new_n246_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n368_), .B1(new_n369_), .B2(new_n248_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n254_), .B1(new_n366_), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n360_), .A2(KEYINPUT32), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n359_), .A2(new_n363_), .A3(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n262_), .B1(new_n351_), .B2(new_n353_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n318_), .A2(new_n263_), .A3(new_n348_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n373_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n369_), .A2(new_n248_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n250_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n206_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n379_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  AOI22_X1  g181(.A1(new_n377_), .A2(new_n378_), .B1(new_n382_), .B2(new_n366_), .ZN(new_n383_));
  AOI22_X1  g182(.A1(new_n365_), .A2(new_n372_), .B1(new_n374_), .B2(new_n383_), .ZN(new_n384_));
  XOR2_X1   g183(.A(G78gat), .B(G106gat), .Z(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT29), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n387_), .B(new_n220_), .C1(new_n230_), .C2(new_n231_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT28), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT28), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n242_), .A2(new_n390_), .A3(new_n387_), .A4(new_n220_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G22gat), .B(G50gat), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n392_), .A2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n389_), .A2(new_n391_), .A3(new_n393_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT94), .ZN(new_n398_));
  NAND2_X1  g197(.A1(KEYINPUT89), .A2(G233gat), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(KEYINPUT89), .A2(G233gat), .ZN(new_n401_));
  OAI21_X1  g200(.A(G228gat), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n387_), .B1(new_n242_), .B2(new_n220_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n403_), .B1(new_n324_), .B2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT93), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  OAI211_X1 g206(.A(KEYINPUT93), .B(new_n403_), .C1(new_n324_), .C2(new_n404_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT94), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n395_), .A2(new_n410_), .A3(new_n396_), .ZN(new_n411_));
  NOR3_X1   g210(.A1(new_n324_), .A2(new_n404_), .A3(new_n403_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  AND4_X1   g212(.A1(new_n398_), .A2(new_n409_), .A3(new_n411_), .A4(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n412_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n398_), .B1(new_n415_), .B2(new_n411_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n386_), .B1(new_n414_), .B2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n409_), .A2(new_n413_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n418_), .A2(KEYINPUT94), .A3(new_n397_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n415_), .A2(new_n398_), .A3(new_n411_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n419_), .A2(new_n385_), .A3(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n417_), .A2(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n202_), .B1(new_n384_), .B2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n377_), .A2(new_n378_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n382_), .A2(new_n366_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n424_), .A2(new_n425_), .A3(new_n374_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n255_), .A2(new_n355_), .A3(new_n364_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n426_), .B1(new_n427_), .B2(new_n371_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n428_), .A2(KEYINPUT100), .A3(new_n421_), .A4(new_n417_), .ZN(new_n429_));
  AOI21_X1  g228(.A(KEYINPUT27), .B1(new_n355_), .B2(new_n364_), .ZN(new_n430_));
  NOR3_X1   g229(.A1(new_n356_), .A2(new_n358_), .A3(new_n262_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n263_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n260_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT101), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT101), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n377_), .A2(new_n435_), .A3(new_n260_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n364_), .A2(KEYINPUT27), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n430_), .B1(new_n437_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n425_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n422_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n423_), .A2(new_n429_), .A3(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G15gat), .B(G43gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT84), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n445_), .B(KEYINPUT30), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(KEYINPUT31), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G227gat), .A2(G233gat), .ZN(new_n448_));
  INV_X1    g247(.A(G71gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  XOR2_X1   g249(.A(new_n450_), .B(G99gat), .Z(new_n451_));
  XNOR2_X1  g250(.A(new_n357_), .B(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n447_), .B(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(KEYINPUT85), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(new_n237_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT85), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n453_), .B(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(new_n236_), .ZN(new_n458_));
  AND3_X1   g257(.A1(new_n455_), .A2(new_n458_), .A3(KEYINPUT86), .ZN(new_n459_));
  AOI21_X1  g258(.A(KEYINPUT86), .B1(new_n455_), .B2(new_n458_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n440_), .A2(KEYINPUT102), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT102), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n438_), .B1(new_n434_), .B2(new_n436_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n463_), .B1(new_n464_), .B2(new_n430_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n422_), .B1(new_n462_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n455_), .A2(new_n458_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n467_), .A2(new_n425_), .ZN(new_n468_));
  AOI22_X1  g267(.A1(new_n443_), .A2(new_n461_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT15), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G29gat), .B(G36gat), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT72), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G43gat), .B(G50gat), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n471_), .B(KEYINPUT72), .ZN(new_n476_));
  INV_X1    g275(.A(new_n474_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n470_), .B1(new_n475_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n473_), .A2(new_n474_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n476_), .A2(new_n477_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n480_), .A2(new_n481_), .A3(KEYINPUT15), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G1gat), .B(G8gat), .ZN(new_n483_));
  OR2_X1    g282(.A1(new_n483_), .A2(KEYINPUT76), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(KEYINPUT76), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G15gat), .B(G22gat), .ZN(new_n487_));
  INV_X1    g286(.A(G1gat), .ZN(new_n488_));
  INV_X1    g287(.A(G8gat), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT14), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n487_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n486_), .A2(new_n491_), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n484_), .A2(new_n490_), .A3(new_n487_), .A4(new_n485_), .ZN(new_n493_));
  AND2_X1   g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n479_), .A2(new_n482_), .A3(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G229gat), .A2(G233gat), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n492_), .A2(new_n493_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n480_), .A2(new_n481_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n497_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n495_), .A2(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n498_), .A2(new_n499_), .ZN(new_n502_));
  AOI22_X1  g301(.A1(new_n480_), .A2(new_n481_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n497_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  XOR2_X1   g303(.A(G113gat), .B(G141gat), .Z(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT79), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G169gat), .B(G197gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n501_), .A2(new_n504_), .A3(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT80), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT81), .ZN(new_n511_));
  AND3_X1   g310(.A1(new_n509_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n511_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n501_), .A2(new_n504_), .ZN(new_n514_));
  OAI22_X1  g313(.A1(new_n512_), .A2(new_n513_), .B1(new_n514_), .B2(new_n508_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n509_), .A2(new_n510_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT81), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n514_), .A2(new_n508_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n509_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n517_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  AND2_X1   g319(.A1(new_n515_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n469_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G232gat), .A2(G233gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT34), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n525_), .A2(KEYINPUT35), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n525_), .A2(KEYINPUT35), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n479_), .A2(new_n482_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT67), .ZN(new_n530_));
  INV_X1    g329(.A(G85gat), .ZN(new_n531_));
  INV_X1    g330(.A(G92gat), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G85gat), .A2(G92gat), .ZN(new_n534_));
  AND2_X1   g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G99gat), .A2(G106gat), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT6), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(G99gat), .A2(G106gat), .ZN(new_n539_));
  NOR2_X1   g338(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  OAI22_X1  g340(.A1(KEYINPUT66), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  OAI211_X1 g342(.A(new_n530_), .B(new_n535_), .C1(new_n538_), .C2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT8), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n544_), .A2(KEYINPUT68), .A3(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(G106gat), .ZN(new_n547_));
  XOR2_X1   g346(.A(KEYINPUT10), .B(G99gat), .Z(new_n548_));
  AOI21_X1  g347(.A(new_n538_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT9), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n534_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT65), .ZN(new_n552_));
  NAND3_X1  g351(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n553_));
  AOI22_X1  g352(.A1(new_n551_), .A2(KEYINPUT64), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n554_), .B1(KEYINPUT64), .B2(new_n551_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n552_), .B1(new_n533_), .B2(new_n553_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n549_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n544_), .A2(KEYINPUT68), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n535_), .B1(new_n538_), .B2(new_n543_), .ZN(new_n559_));
  OAI21_X1  g358(.A(KEYINPUT8), .B1(new_n559_), .B2(KEYINPUT68), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n546_), .B(new_n557_), .C1(new_n558_), .C2(new_n560_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n529_), .A2(new_n561_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n499_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n528_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT75), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n562_), .A2(new_n563_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(new_n526_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT74), .ZN(new_n569_));
  OAI211_X1 g368(.A(KEYINPUT75), .B(new_n528_), .C1(new_n562_), .C2(new_n563_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n566_), .A2(new_n568_), .A3(new_n569_), .A4(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G190gat), .B(G218gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT73), .ZN(new_n573_));
  XOR2_X1   g372(.A(G134gat), .B(G162gat), .Z(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n576_), .A2(KEYINPUT36), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n571_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n528_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n563_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n529_), .A2(new_n561_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n580_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  AOI22_X1  g382(.A1(new_n583_), .A2(KEYINPUT75), .B1(new_n567_), .B2(new_n526_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n584_), .A2(new_n569_), .A3(new_n566_), .A4(new_n577_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n579_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(new_n566_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n587_), .A2(KEYINPUT36), .A3(new_n576_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n586_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(KEYINPUT37), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G57gat), .B(G64gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G71gat), .B(G78gat), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n591_), .A2(new_n592_), .A3(KEYINPUT11), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(KEYINPUT11), .ZN(new_n594_));
  INV_X1    g393(.A(new_n592_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n591_), .A2(KEYINPUT11), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n593_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(G231gat), .A2(G233gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT77), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n598_), .B(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(new_n498_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  XOR2_X1   g402(.A(G127gat), .B(G155gat), .Z(new_n604_));
  XNOR2_X1  g403(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G183gat), .B(G211gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT69), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n609_), .A2(new_n610_), .A3(KEYINPUT17), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n603_), .A2(new_n611_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n611_), .B1(KEYINPUT17), .B2(new_n609_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(new_n602_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT37), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n586_), .A2(new_n616_), .A3(new_n588_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n590_), .A2(new_n615_), .A3(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n598_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n561_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT12), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n598_), .A2(new_n610_), .ZN(new_n622_));
  OAI211_X1 g421(.A(KEYINPUT69), .B(new_n593_), .C1(new_n596_), .C2(new_n597_), .ZN(new_n623_));
  AND3_X1   g422(.A1(new_n622_), .A2(KEYINPUT12), .A3(new_n623_), .ZN(new_n624_));
  AOI22_X1  g423(.A1(new_n620_), .A2(new_n621_), .B1(new_n561_), .B2(new_n624_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n546_), .A2(new_n557_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n544_), .A2(KEYINPUT68), .ZN(new_n627_));
  OAI211_X1 g426(.A(new_n627_), .B(KEYINPUT8), .C1(KEYINPUT68), .C2(new_n559_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n626_), .A2(new_n628_), .A3(new_n598_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT70), .ZN(new_n630_));
  NAND2_X1  g429(.A1(G230gat), .A2(G233gat), .ZN(new_n631_));
  AND3_X1   g430(.A1(new_n629_), .A2(new_n630_), .A3(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n630_), .B1(new_n629_), .B2(new_n631_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n625_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT71), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n631_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n629_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n598_), .B1(new_n626_), .B2(new_n628_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n637_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n625_), .B(KEYINPUT71), .C1(new_n632_), .C2(new_n633_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n636_), .A2(new_n640_), .A3(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(G120gat), .B(G148gat), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT5), .ZN(new_n644_));
  XNOR2_X1  g443(.A(G176gat), .B(G204gat), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n644_), .B(new_n645_), .Z(new_n646_));
  NAND2_X1  g445(.A1(new_n642_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n646_), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n636_), .A2(new_n640_), .A3(new_n641_), .A4(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT13), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n650_), .B(new_n651_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n618_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n523_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n655_), .A2(new_n488_), .A3(new_n425_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT38), .ZN(new_n657_));
  INV_X1    g456(.A(new_n615_), .ZN(new_n658_));
  NOR3_X1   g457(.A1(new_n652_), .A2(new_n522_), .A3(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT103), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n443_), .A2(new_n461_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n466_), .A2(new_n468_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT104), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n589_), .B(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n663_), .A2(KEYINPUT105), .A3(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT105), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n668_), .B1(new_n469_), .B2(new_n665_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n660_), .B1(new_n667_), .B2(new_n669_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n670_), .A2(new_n425_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n657_), .B1(new_n671_), .B2(new_n488_), .ZN(G1324gat));
  NAND2_X1  g471(.A1(new_n462_), .A2(new_n465_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n655_), .A2(new_n489_), .A3(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT39), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n670_), .A2(new_n674_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n676_), .B1(new_n677_), .B2(G8gat), .ZN(new_n678_));
  AOI211_X1 g477(.A(KEYINPUT39), .B(new_n489_), .C1(new_n670_), .C2(new_n674_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n675_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT40), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n680_), .B(new_n681_), .ZN(G1325gat));
  INV_X1    g481(.A(new_n461_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n670_), .A2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(G15gat), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(KEYINPUT106), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT106), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n684_), .A2(new_n687_), .A3(G15gat), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT41), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  OR3_X1    g490(.A1(new_n654_), .A2(G15gat), .A3(new_n461_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n686_), .A2(KEYINPUT41), .A3(new_n688_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n691_), .A2(new_n692_), .A3(new_n693_), .ZN(G1326gat));
  INV_X1    g493(.A(G22gat), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n655_), .A2(new_n695_), .A3(new_n422_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT42), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n670_), .A2(new_n422_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n697_), .B1(new_n698_), .B2(G22gat), .ZN(new_n699_));
  AOI211_X1 g498(.A(KEYINPUT42), .B(new_n695_), .C1(new_n670_), .C2(new_n422_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n696_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT107), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n701_), .B(new_n702_), .ZN(G1327gat));
  NOR3_X1   g502(.A1(new_n652_), .A2(new_n522_), .A3(new_n615_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT43), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n586_), .A2(new_n616_), .A3(new_n588_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n616_), .B1(new_n586_), .B2(new_n588_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n705_), .B1(new_n663_), .B2(new_n709_), .ZN(new_n710_));
  NOR3_X1   g509(.A1(new_n469_), .A2(KEYINPUT43), .A3(new_n708_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n704_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n663_), .A2(new_n705_), .A3(new_n709_), .ZN(new_n715_));
  OAI21_X1  g514(.A(KEYINPUT43), .B1(new_n469_), .B2(new_n708_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n717_), .A2(KEYINPUT44), .A3(new_n704_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n714_), .A2(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(G29gat), .B1(new_n719_), .B2(new_n441_), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n666_), .A2(new_n652_), .A3(new_n615_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n523_), .A2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(G29gat), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n425_), .A2(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n720_), .B1(new_n723_), .B2(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT108), .ZN(G1328gat));
  NOR2_X1   g526(.A1(new_n673_), .A2(G36gat), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n722_), .A2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(KEYINPUT45), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT45), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n722_), .A2(new_n731_), .A3(new_n728_), .ZN(new_n732_));
  AND3_X1   g531(.A1(new_n730_), .A2(KEYINPUT110), .A3(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(KEYINPUT110), .A2(G36gat), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n714_), .A2(new_n674_), .A3(new_n718_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT109), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n734_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n714_), .A2(KEYINPUT109), .A3(new_n674_), .A4(new_n718_), .ZN(new_n738_));
  AOI211_X1 g537(.A(KEYINPUT46), .B(new_n733_), .C1(new_n737_), .C2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT46), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n735_), .A2(new_n736_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n734_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n741_), .A2(new_n738_), .A3(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n733_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n740_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n739_), .A2(new_n745_), .ZN(G1329gat));
  INV_X1    g545(.A(G43gat), .ZN(new_n747_));
  OR3_X1    g546(.A1(new_n719_), .A2(new_n747_), .A3(new_n467_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n747_), .B1(new_n723_), .B2(new_n461_), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n748_), .A2(KEYINPUT47), .A3(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(KEYINPUT47), .B1(new_n748_), .B2(new_n749_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n750_), .A2(new_n751_), .ZN(G1330gat));
  INV_X1    g551(.A(G50gat), .ZN(new_n753_));
  INV_X1    g552(.A(new_n422_), .ZN(new_n754_));
  NOR3_X1   g553(.A1(new_n719_), .A2(new_n753_), .A3(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(G50gat), .B1(new_n722_), .B2(new_n422_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n755_), .A2(new_n756_), .ZN(G1331gat));
  INV_X1    g556(.A(G57gat), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n469_), .A2(new_n521_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n650_), .B(KEYINPUT13), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n618_), .A2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n758_), .B1(new_n762_), .B2(new_n441_), .ZN(new_n763_));
  XOR2_X1   g562(.A(new_n763_), .B(KEYINPUT111), .Z(new_n764_));
  NAND3_X1  g563(.A1(new_n652_), .A2(new_n522_), .A3(new_n615_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n765_), .B1(new_n667_), .B2(new_n669_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n441_), .A2(new_n758_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n764_), .B1(new_n766_), .B2(new_n767_), .ZN(G1332gat));
  OR3_X1    g567(.A1(new_n762_), .A2(G64gat), .A3(new_n673_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n766_), .ZN(new_n770_));
  OAI21_X1  g569(.A(G64gat), .B1(new_n770_), .B2(new_n673_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n771_), .A2(KEYINPUT48), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n771_), .A2(KEYINPUT48), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n769_), .B1(new_n772_), .B2(new_n773_), .ZN(G1333gat));
  OAI21_X1  g573(.A(G71gat), .B1(new_n770_), .B2(new_n461_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n775_), .A2(KEYINPUT49), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n775_), .A2(KEYINPUT49), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n683_), .A2(new_n449_), .ZN(new_n778_));
  OAI22_X1  g577(.A1(new_n776_), .A2(new_n777_), .B1(new_n762_), .B2(new_n778_), .ZN(G1334gat));
  INV_X1    g578(.A(KEYINPUT50), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n766_), .A2(new_n422_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n780_), .B1(new_n781_), .B2(G78gat), .ZN(new_n782_));
  INV_X1    g581(.A(G78gat), .ZN(new_n783_));
  AOI211_X1 g582(.A(KEYINPUT50), .B(new_n783_), .C1(new_n766_), .C2(new_n422_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n422_), .A2(new_n783_), .ZN(new_n785_));
  OAI22_X1  g584(.A1(new_n782_), .A2(new_n784_), .B1(new_n762_), .B2(new_n785_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT112), .ZN(G1335gat));
  NAND3_X1  g586(.A1(new_n652_), .A2(new_n522_), .A3(new_n658_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n717_), .A2(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(G85gat), .B1(new_n790_), .B2(new_n441_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n759_), .A2(new_n665_), .A3(new_n652_), .A4(new_n658_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n425_), .A2(new_n531_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n791_), .B1(new_n792_), .B2(new_n793_), .ZN(G1336gat));
  OAI21_X1  g593(.A(G92gat), .B1(new_n790_), .B2(new_n673_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n674_), .A2(new_n532_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n795_), .B1(new_n792_), .B2(new_n796_), .ZN(G1337gat));
  OAI21_X1  g596(.A(G99gat), .B1(new_n790_), .B2(new_n461_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n548_), .ZN(new_n799_));
  OR3_X1    g598(.A1(new_n792_), .A2(new_n467_), .A3(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n798_), .A2(new_n800_), .A3(KEYINPUT114), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT113), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT51), .ZN(new_n803_));
  NOR3_X1   g602(.A1(new_n801_), .A2(new_n802_), .A3(new_n803_), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n801_), .A2(new_n803_), .ZN(new_n805_));
  AOI21_X1  g604(.A(KEYINPUT113), .B1(new_n798_), .B2(new_n800_), .ZN(new_n806_));
  NOR3_X1   g605(.A1(new_n804_), .A2(new_n805_), .A3(new_n806_), .ZN(G1338gat));
  NOR3_X1   g606(.A1(new_n792_), .A2(G106gat), .A3(new_n754_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT115), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n808_), .B(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n788_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n547_), .B1(new_n811_), .B2(new_n422_), .ZN(new_n812_));
  OR2_X1    g611(.A1(new_n812_), .A2(KEYINPUT52), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(KEYINPUT52), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n810_), .A2(new_n813_), .A3(new_n814_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n815_), .B(new_n817_), .ZN(G1339gat));
  INV_X1    g617(.A(KEYINPUT117), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n708_), .A2(new_n760_), .A3(new_n522_), .A4(new_n615_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n819_), .B1(new_n820_), .B2(KEYINPUT54), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n653_), .A2(KEYINPUT117), .A3(new_n822_), .A4(new_n522_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n820_), .A2(KEYINPUT54), .ZN(new_n824_));
  AND3_X1   g623(.A1(new_n821_), .A2(new_n823_), .A3(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT57), .ZN(new_n826_));
  OR2_X1    g625(.A1(new_n502_), .A2(new_n503_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n508_), .B1(new_n827_), .B2(new_n496_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n503_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n495_), .A2(new_n829_), .A3(new_n497_), .ZN(new_n830_));
  AOI22_X1  g629(.A1(new_n514_), .A2(new_n508_), .B1(new_n828_), .B2(new_n830_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n650_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT55), .ZN(new_n833_));
  AND3_X1   g632(.A1(new_n636_), .A2(new_n833_), .A3(new_n641_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n624_), .A2(new_n561_), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n835_), .B(new_n629_), .C1(new_n639_), .C2(KEYINPUT12), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n637_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(KEYINPUT118), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT118), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n836_), .A2(new_n839_), .A3(new_n637_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n840_), .ZN(new_n841_));
  OAI211_X1 g640(.A(KEYINPUT55), .B(new_n625_), .C1(new_n632_), .C2(new_n633_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n646_), .B1(new_n834_), .B2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT56), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT119), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n636_), .A2(new_n833_), .A3(new_n641_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n848_), .A2(new_n842_), .A3(new_n841_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n849_), .A2(KEYINPUT56), .A3(new_n646_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n846_), .A2(new_n847_), .A3(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n521_), .A2(new_n649_), .ZN(new_n852_));
  AOI21_X1  g651(.A(KEYINPUT56), .B1(new_n849_), .B2(new_n646_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n852_), .B1(new_n853_), .B2(KEYINPUT119), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n832_), .B1(new_n851_), .B2(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n826_), .B1(new_n855_), .B2(new_n665_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT120), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  OAI211_X1 g657(.A(KEYINPUT120), .B(new_n826_), .C1(new_n855_), .C2(new_n665_), .ZN(new_n859_));
  OR3_X1    g658(.A1(new_n855_), .A2(new_n826_), .A3(new_n665_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT58), .ZN(new_n861_));
  AND2_X1   g660(.A1(new_n846_), .A2(new_n850_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n649_), .A2(new_n831_), .ZN(new_n863_));
  OAI211_X1 g662(.A(KEYINPUT121), .B(new_n861_), .C1(new_n862_), .C2(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n863_), .B1(new_n846_), .B2(new_n850_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT121), .ZN(new_n866_));
  OAI21_X1  g665(.A(KEYINPUT58), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n864_), .A2(new_n709_), .A3(new_n867_), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n858_), .A2(new_n859_), .A3(new_n860_), .A4(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n825_), .B1(new_n869_), .B2(new_n658_), .ZN(new_n870_));
  NOR4_X1   g669(.A1(new_n674_), .A2(new_n441_), .A3(new_n422_), .A4(new_n467_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(KEYINPUT59), .B1(new_n870_), .B2(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n821_), .A2(new_n823_), .A3(new_n824_), .ZN(new_n874_));
  AND3_X1   g673(.A1(new_n860_), .A2(new_n856_), .A3(new_n868_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n875_), .B2(new_n615_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT59), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n876_), .A2(new_n877_), .A3(new_n871_), .ZN(new_n878_));
  INV_X1    g677(.A(G113gat), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n522_), .A2(new_n879_), .ZN(new_n880_));
  AND3_X1   g679(.A1(new_n873_), .A2(new_n878_), .A3(new_n880_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n870_), .A2(new_n872_), .ZN(new_n882_));
  AOI21_X1  g681(.A(G113gat), .B1(new_n882_), .B2(new_n521_), .ZN(new_n883_));
  OAI21_X1  g682(.A(KEYINPUT122), .B1(new_n881_), .B2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n869_), .A2(new_n658_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n874_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(new_n871_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n879_), .B1(new_n887_), .B2(new_n522_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT122), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n873_), .A2(new_n878_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n880_), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n888_), .B(new_n889_), .C1(new_n890_), .C2(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n884_), .A2(new_n892_), .ZN(G1340gat));
  OAI21_X1  g692(.A(G120gat), .B1(new_n890_), .B2(new_n760_), .ZN(new_n894_));
  INV_X1    g693(.A(G120gat), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n895_), .B1(new_n760_), .B2(KEYINPUT60), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n896_), .B1(KEYINPUT60), .B2(new_n895_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n894_), .B1(new_n887_), .B2(new_n897_), .ZN(G1341gat));
  OAI21_X1  g697(.A(G127gat), .B1(new_n890_), .B2(new_n658_), .ZN(new_n899_));
  OR2_X1    g698(.A1(new_n658_), .A2(G127gat), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n899_), .B1(new_n887_), .B2(new_n900_), .ZN(G1342gat));
  OAI21_X1  g700(.A(G134gat), .B1(new_n890_), .B2(new_n708_), .ZN(new_n902_));
  OR2_X1    g701(.A1(new_n666_), .A2(G134gat), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n902_), .B1(new_n887_), .B2(new_n903_), .ZN(G1343gat));
  NOR2_X1   g703(.A1(new_n683_), .A2(new_n754_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n905_), .A2(new_n673_), .A3(new_n425_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n870_), .A2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(new_n521_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g708(.A1(new_n907_), .A2(new_n652_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g710(.A(KEYINPUT61), .B(G155gat), .ZN(new_n912_));
  INV_X1    g711(.A(new_n912_), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT123), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n907_), .A2(new_n914_), .A3(new_n615_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n914_), .B1(new_n907_), .B2(new_n615_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n913_), .B1(new_n916_), .B2(new_n917_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n906_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n886_), .A2(new_n919_), .ZN(new_n920_));
  OAI21_X1  g719(.A(KEYINPUT123), .B1(new_n920_), .B2(new_n658_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n921_), .A2(new_n915_), .A3(new_n912_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n918_), .A2(new_n922_), .ZN(G1346gat));
  OAI21_X1  g722(.A(G162gat), .B1(new_n920_), .B2(new_n708_), .ZN(new_n924_));
  INV_X1    g723(.A(G162gat), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n665_), .A2(new_n925_), .ZN(new_n926_));
  OAI211_X1 g725(.A(new_n924_), .B(KEYINPUT124), .C1(new_n920_), .C2(new_n926_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT124), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n920_), .A2(new_n926_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n925_), .B1(new_n907_), .B2(new_n709_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n928_), .B1(new_n929_), .B2(new_n930_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n927_), .A2(new_n931_), .ZN(G1347gat));
  AND2_X1   g731(.A1(new_n876_), .A2(new_n754_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n673_), .A2(new_n425_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n683_), .A2(new_n934_), .ZN(new_n935_));
  INV_X1    g734(.A(new_n935_), .ZN(new_n936_));
  AND2_X1   g735(.A1(new_n933_), .A2(new_n936_), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n937_), .A2(new_n313_), .A3(new_n521_), .ZN(new_n938_));
  OAI21_X1  g737(.A(KEYINPUT125), .B1(new_n935_), .B2(new_n522_), .ZN(new_n939_));
  INV_X1    g738(.A(KEYINPUT125), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n936_), .A2(new_n940_), .A3(new_n521_), .ZN(new_n941_));
  NAND4_X1  g740(.A1(new_n876_), .A2(new_n754_), .A3(new_n939_), .A4(new_n941_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n942_), .A2(G169gat), .ZN(new_n943_));
  AND2_X1   g742(.A1(new_n943_), .A2(KEYINPUT62), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n943_), .A2(KEYINPUT62), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n938_), .B1(new_n944_), .B2(new_n945_), .ZN(G1348gat));
  NAND2_X1  g745(.A1(new_n937_), .A2(new_n652_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n870_), .A2(new_n422_), .ZN(new_n948_));
  NOR3_X1   g747(.A1(new_n935_), .A2(new_n314_), .A3(new_n760_), .ZN(new_n949_));
  AOI22_X1  g748(.A1(new_n947_), .A2(new_n314_), .B1(new_n948_), .B2(new_n949_), .ZN(G1349gat));
  NOR2_X1   g749(.A1(new_n935_), .A2(new_n658_), .ZN(new_n951_));
  AOI21_X1  g750(.A(G183gat), .B1(new_n948_), .B2(new_n951_), .ZN(new_n952_));
  NOR3_X1   g751(.A1(new_n935_), .A2(new_n302_), .A3(new_n658_), .ZN(new_n953_));
  AOI21_X1  g752(.A(new_n952_), .B1(new_n933_), .B2(new_n953_), .ZN(G1350gat));
  NAND3_X1  g753(.A1(new_n937_), .A2(new_n303_), .A3(new_n665_), .ZN(new_n955_));
  AND3_X1   g754(.A1(new_n933_), .A2(new_n709_), .A3(new_n936_), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n955_), .B1(new_n329_), .B2(new_n956_), .ZN(G1351gat));
  NAND2_X1  g756(.A1(new_n905_), .A2(new_n934_), .ZN(new_n958_));
  NOR2_X1   g757(.A1(new_n870_), .A2(new_n958_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n959_), .A2(new_n521_), .ZN(new_n960_));
  XNOR2_X1  g759(.A(new_n960_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g760(.A1(new_n959_), .A2(new_n269_), .A3(new_n652_), .ZN(new_n962_));
  INV_X1    g761(.A(new_n962_), .ZN(new_n963_));
  AOI21_X1  g762(.A(G204gat), .B1(new_n959_), .B2(new_n652_), .ZN(new_n964_));
  OAI21_X1  g763(.A(KEYINPUT126), .B1(new_n963_), .B2(new_n964_), .ZN(new_n965_));
  INV_X1    g764(.A(new_n958_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n886_), .A2(new_n966_), .ZN(new_n967_));
  OAI21_X1  g766(.A(new_n266_), .B1(new_n967_), .B2(new_n760_), .ZN(new_n968_));
  INV_X1    g767(.A(KEYINPUT126), .ZN(new_n969_));
  NAND3_X1  g768(.A1(new_n968_), .A2(new_n969_), .A3(new_n962_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n965_), .A2(new_n970_), .ZN(G1353gat));
  NAND2_X1  g770(.A1(new_n959_), .A2(new_n615_), .ZN(new_n972_));
  NOR2_X1   g771(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n973_));
  AND2_X1   g772(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n974_));
  NOR3_X1   g773(.A1(new_n972_), .A2(new_n973_), .A3(new_n974_), .ZN(new_n975_));
  AOI21_X1  g774(.A(new_n975_), .B1(new_n972_), .B2(new_n973_), .ZN(G1354gat));
  NAND2_X1  g775(.A1(new_n959_), .A2(new_n665_), .ZN(new_n977_));
  XNOR2_X1  g776(.A(KEYINPUT127), .B(G218gat), .ZN(new_n978_));
  NOR2_X1   g777(.A1(new_n708_), .A2(new_n978_), .ZN(new_n979_));
  AOI22_X1  g778(.A1(new_n977_), .A2(new_n978_), .B1(new_n959_), .B2(new_n979_), .ZN(G1355gat));
endmodule


