//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 1 0 1 1 0 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n701_, new_n702_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n838_, new_n839_, new_n840_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n854_, new_n855_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_, new_n884_, new_n886_, new_n887_,
    new_n889_, new_n890_, new_n892_, new_n893_, new_n894_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G29gat), .B(G36gat), .ZN(new_n203_));
  AND2_X1   g002(.A1(new_n203_), .A2(KEYINPUT71), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n203_), .A2(KEYINPUT71), .ZN(new_n205_));
  XOR2_X1   g004(.A(G43gat), .B(G50gat), .Z(new_n206_));
  OR3_X1    g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n206_), .B1(new_n204_), .B2(new_n205_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G15gat), .B(G22gat), .ZN(new_n210_));
  INV_X1    g009(.A(G8gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G1gat), .B(G8gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n209_), .A2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(KEYINPUT76), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G229gat), .A2(G233gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT15), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n209_), .A2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n207_), .A2(new_n208_), .A3(KEYINPUT15), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n221_), .A2(new_n215_), .A3(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT77), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT77), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n221_), .A2(new_n225_), .A3(new_n215_), .A4(new_n222_), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n218_), .A2(new_n219_), .A3(new_n224_), .A4(new_n226_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n217_), .A2(KEYINPUT76), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT76), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n229_), .B1(new_n209_), .B2(new_n216_), .ZN(new_n230_));
  OAI22_X1  g029(.A1(new_n228_), .A2(new_n230_), .B1(new_n216_), .B2(new_n209_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n219_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n227_), .A2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G113gat), .B(G141gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G169gat), .B(G197gat), .ZN(new_n236_));
  XOR2_X1   g035(.A(new_n235_), .B(new_n236_), .Z(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n234_), .A2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n227_), .A2(new_n233_), .A3(new_n237_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G120gat), .B(G148gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT5), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G176gat), .B(G204gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G99gat), .A2(G106gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(KEYINPUT6), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT6), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n249_), .A2(G99gat), .A3(G106gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT9), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n252_), .A2(G85gat), .A3(G92gat), .ZN(new_n253_));
  AND2_X1   g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  XOR2_X1   g053(.A(G85gat), .B(G92gat), .Z(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT9), .ZN(new_n256_));
  XOR2_X1   g055(.A(KEYINPUT10), .B(G99gat), .Z(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT64), .B(G106gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n254_), .A2(new_n256_), .A3(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT65), .ZN(new_n261_));
  INV_X1    g060(.A(G99gat), .ZN(new_n262_));
  INV_X1    g061(.A(G106gat), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n261_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT7), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT7), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n261_), .A2(new_n266_), .A3(new_n262_), .A4(new_n263_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n265_), .A2(new_n251_), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT8), .ZN(new_n269_));
  AND3_X1   g068(.A1(new_n268_), .A2(new_n269_), .A3(new_n255_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n269_), .B1(new_n268_), .B2(new_n255_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n260_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT66), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  OAI211_X1 g073(.A(KEYINPUT66), .B(new_n260_), .C1(new_n270_), .C2(new_n271_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G57gat), .B(G64gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G71gat), .B(G78gat), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n276_), .A2(new_n277_), .A3(KEYINPUT11), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n276_), .A2(KEYINPUT11), .ZN(new_n279_));
  INV_X1    g078(.A(new_n277_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n276_), .A2(KEYINPUT11), .ZN(new_n282_));
  OAI211_X1 g081(.A(KEYINPUT12), .B(new_n278_), .C1(new_n281_), .C2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n274_), .A2(new_n275_), .A3(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G230gat), .A2(G233gat), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT12), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n268_), .A2(new_n255_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT8), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n268_), .A2(new_n269_), .A3(new_n255_), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n256_), .A2(new_n259_), .ZN(new_n291_));
  AOI22_X1  g090(.A1(new_n289_), .A2(new_n290_), .B1(new_n254_), .B2(new_n291_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n278_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n287_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  OAI211_X1 g093(.A(new_n293_), .B(new_n260_), .C1(new_n270_), .C2(new_n271_), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n285_), .A2(new_n286_), .A3(new_n294_), .A4(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n292_), .A2(new_n293_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n295_), .ZN(new_n298_));
  OAI211_X1 g097(.A(G230gat), .B(G233gat), .C1(new_n297_), .C2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n296_), .A2(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n246_), .B1(new_n300_), .B2(KEYINPUT67), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT67), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n296_), .A2(new_n302_), .A3(new_n299_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n296_), .A2(new_n299_), .A3(new_n246_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT68), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT68), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n296_), .A2(new_n307_), .A3(new_n299_), .A4(new_n246_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n304_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n311_));
  OR2_X1    g110(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n310_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  AND2_X1   g112(.A1(new_n310_), .A2(new_n312_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G228gat), .A2(G233gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT89), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT94), .ZN(new_n318_));
  OR2_X1    g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G22gat), .B(G50gat), .ZN(new_n320_));
  XOR2_X1   g119(.A(new_n319_), .B(new_n320_), .Z(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT90), .B(G197gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(G204gat), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT21), .ZN(new_n325_));
  INV_X1    g124(.A(G197gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT91), .B(G204gat), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n324_), .B(new_n325_), .C1(new_n326_), .C2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT92), .ZN(new_n329_));
  INV_X1    g128(.A(new_n327_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(G197gat), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT92), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n331_), .A2(new_n332_), .A3(new_n325_), .A4(new_n324_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n329_), .A2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G211gat), .B(G218gat), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  OAI22_X1  g135(.A1(new_n330_), .A2(G197gat), .B1(new_n323_), .B2(G204gat), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n336_), .B1(new_n337_), .B2(KEYINPUT21), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n334_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT93), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n324_), .B(new_n340_), .C1(new_n326_), .C2(new_n327_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n335_), .A2(new_n325_), .ZN(new_n342_));
  AND2_X1   g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n331_), .A2(new_n324_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT93), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n339_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n317_), .A2(new_n318_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(G155gat), .A2(G162gat), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G155gat), .A2(G162gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT1), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT1), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n353_), .A2(G155gat), .A3(G162gat), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n350_), .A2(new_n352_), .A3(new_n354_), .ZN(new_n355_));
  XOR2_X1   g154(.A(G141gat), .B(G148gat), .Z(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(KEYINPUT86), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT86), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n355_), .A2(new_n359_), .A3(new_n356_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(G141gat), .A2(G148gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT3), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G141gat), .A2(G148gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT2), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  AND2_X1   g164(.A1(new_n350_), .A2(new_n351_), .ZN(new_n366_));
  AOI22_X1  g165(.A1(new_n358_), .A2(new_n360_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT29), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n348_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(G78gat), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n347_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  AOI22_X1  g171(.A1(new_n334_), .A2(new_n338_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n373_));
  OAI21_X1  g172(.A(G78gat), .B1(new_n373_), .B2(new_n369_), .ZN(new_n374_));
  AND3_X1   g173(.A1(new_n372_), .A2(new_n374_), .A3(G106gat), .ZN(new_n375_));
  AOI21_X1  g174(.A(G106gat), .B1(new_n372_), .B2(new_n374_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n358_), .A2(new_n360_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n365_), .A2(new_n366_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(KEYINPUT87), .B1(new_n379_), .B2(KEYINPUT29), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT87), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n367_), .A2(new_n381_), .A3(new_n368_), .ZN(new_n382_));
  XOR2_X1   g181(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  AND3_X1   g183(.A1(new_n380_), .A2(new_n382_), .A3(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n384_), .B1(new_n380_), .B2(new_n382_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NOR3_X1   g186(.A1(new_n375_), .A2(new_n376_), .A3(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n386_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n380_), .A2(new_n382_), .A3(new_n384_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n371_), .B1(new_n347_), .B2(new_n370_), .ZN(new_n392_));
  NOR3_X1   g191(.A1(new_n373_), .A2(new_n369_), .A3(G78gat), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n263_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n372_), .A2(new_n374_), .A3(G106gat), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n391_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n322_), .B1(new_n388_), .B2(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n387_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n394_), .A2(new_n395_), .A3(new_n391_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n398_), .A2(new_n399_), .A3(new_n321_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n397_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G226gat), .A2(G233gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(KEYINPUT19), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT23), .ZN(new_n406_));
  INV_X1    g205(.A(G183gat), .ZN(new_n407_));
  INV_X1    g206(.A(G190gat), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n406_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n409_), .B(new_n410_), .C1(G183gat), .C2(G190gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G169gat), .A2(G176gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT22), .B(G169gat), .ZN(new_n413_));
  INV_X1    g212(.A(G176gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  AND3_X1   g214(.A1(new_n411_), .A2(new_n412_), .A3(new_n415_), .ZN(new_n416_));
  OR2_X1    g215(.A1(new_n416_), .A2(KEYINPUT97), .ZN(new_n417_));
  NOR2_X1   g216(.A1(G169gat), .A2(G176gat), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT24), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n409_), .A2(new_n420_), .A3(new_n410_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT96), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT25), .B(G183gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(KEYINPUT26), .B(G190gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n412_), .A2(KEYINPUT24), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n418_), .B1(new_n427_), .B2(KEYINPUT95), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n428_), .B1(KEYINPUT95), .B2(new_n427_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n423_), .A2(new_n426_), .A3(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n416_), .A2(KEYINPUT97), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n417_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n432_));
  OAI211_X1 g231(.A(KEYINPUT20), .B(new_n405_), .C1(new_n347_), .C2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  AND2_X1   g233(.A1(new_n411_), .A2(new_n412_), .ZN(new_n435_));
  INV_X1    g234(.A(G169gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT22), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(KEYINPUT78), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n414_), .B(new_n438_), .C1(new_n413_), .C2(KEYINPUT78), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(KEYINPUT79), .ZN(new_n440_));
  AOI21_X1  g239(.A(G176gat), .B1(new_n437_), .B2(KEYINPUT78), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT79), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n441_), .B(new_n442_), .C1(KEYINPUT78), .C2(new_n413_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n435_), .A2(new_n440_), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT80), .ZN(new_n445_));
  INV_X1    g244(.A(new_n421_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n446_), .B(new_n426_), .C1(new_n418_), .C2(new_n427_), .ZN(new_n447_));
  AND3_X1   g246(.A1(new_n444_), .A2(new_n445_), .A3(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n445_), .B1(new_n444_), .B2(new_n447_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NOR3_X1   g249(.A1(new_n450_), .A2(KEYINPUT98), .A3(new_n373_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT98), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n444_), .A2(new_n447_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT80), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n444_), .A2(new_n445_), .A3(new_n447_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n452_), .B1(new_n456_), .B2(new_n347_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n434_), .B1(new_n451_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n347_), .A2(new_n432_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT20), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n456_), .A2(new_n347_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n404_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  XOR2_X1   g261(.A(G8gat), .B(G36gat), .Z(new_n463_));
  XNOR2_X1  g262(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G64gat), .B(G92gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n465_), .B(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n458_), .A2(new_n462_), .A3(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n450_), .A2(new_n373_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT20), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n470_), .B1(new_n347_), .B2(new_n432_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n469_), .A2(new_n471_), .A3(new_n405_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n416_), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n430_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(new_n373_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT20), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n478_), .B1(new_n451_), .B2(new_n457_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n473_), .B1(new_n479_), .B2(new_n404_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n467_), .B(KEYINPUT105), .ZN(new_n481_));
  OAI211_X1 g280(.A(KEYINPUT27), .B(new_n468_), .C1(new_n480_), .C2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT27), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n467_), .B1(new_n458_), .B2(new_n462_), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT98), .B1(new_n450_), .B2(new_n373_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n456_), .A2(new_n452_), .A3(new_n347_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n433_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n405_), .B1(new_n469_), .B2(new_n471_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n467_), .ZN(new_n489_));
  NOR3_X1   g288(.A1(new_n487_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n483_), .B1(new_n484_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n482_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G225gat), .A2(G233gat), .ZN(new_n493_));
  XOR2_X1   g292(.A(new_n493_), .B(KEYINPUT102), .Z(new_n494_));
  XNOR2_X1  g293(.A(G127gat), .B(G134gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT83), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G113gat), .B(G120gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT83), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n495_), .B(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n497_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n498_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n379_), .A2(new_n503_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n494_), .B1(new_n504_), .B2(KEYINPUT4), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n367_), .A2(new_n498_), .A3(new_n502_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n504_), .A2(new_n506_), .A3(KEYINPUT4), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT101), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT101), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n504_), .A2(new_n506_), .A3(new_n509_), .A4(KEYINPUT4), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n505_), .B1(new_n508_), .B2(new_n510_), .ZN(new_n511_));
  AND3_X1   g310(.A1(new_n504_), .A2(new_n506_), .A3(new_n493_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G1gat), .B(G29gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(G85gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(KEYINPUT0), .B(G57gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n513_), .B(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n402_), .B1(new_n492_), .B2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT30), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n456_), .A2(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n454_), .A2(KEYINPUT30), .A3(new_n455_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G71gat), .B(G99gat), .ZN(new_n524_));
  INV_X1    g323(.A(G43gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G227gat), .A2(G233gat), .ZN(new_n527_));
  INV_X1    g326(.A(G15gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n526_), .B(new_n529_), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n522_), .A2(KEYINPUT81), .A3(new_n523_), .A4(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n522_), .A2(KEYINPUT81), .A3(new_n523_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n530_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(KEYINPUT81), .B1(new_n522_), .B2(new_n523_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n531_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  XOR2_X1   g335(.A(new_n503_), .B(KEYINPUT31), .Z(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT82), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n537_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT84), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n538_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT85), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n536_), .A2(new_n542_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n544_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n546_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n542_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n549_));
  OAI21_X1  g348(.A(KEYINPUT85), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n547_), .A2(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n477_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n472_), .B1(new_n552_), .B2(new_n405_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n467_), .A2(KEYINPUT32), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT104), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(new_n519_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n458_), .A2(new_n462_), .A3(new_n554_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n557_), .B1(new_n556_), .B2(new_n560_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n401_), .B1(new_n559_), .B2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n513_), .A2(KEYINPUT33), .A3(new_n518_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT100), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n564_), .B1(new_n484_), .B2(new_n490_), .ZN(new_n565_));
  AOI21_X1  g364(.A(KEYINPUT33), .B1(new_n513_), .B2(new_n518_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n493_), .B1(new_n504_), .B2(KEYINPUT4), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n567_), .B1(new_n508_), .B2(new_n510_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n504_), .A2(new_n506_), .A3(new_n494_), .ZN(new_n569_));
  AOI21_X1  g368(.A(KEYINPUT103), .B1(new_n569_), .B2(new_n517_), .ZN(new_n570_));
  AND3_X1   g369(.A1(new_n569_), .A2(KEYINPUT103), .A3(new_n517_), .ZN(new_n571_));
  NOR3_X1   g370(.A1(new_n568_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n566_), .A2(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n489_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n468_), .A2(new_n574_), .A3(KEYINPUT100), .ZN(new_n575_));
  AND4_X1   g374(.A1(new_n563_), .A2(new_n565_), .A3(new_n573_), .A4(new_n575_), .ZN(new_n576_));
  OAI211_X1 g375(.A(new_n520_), .B(new_n551_), .C1(new_n562_), .C2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n401_), .A2(new_n482_), .A3(new_n491_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT106), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n513_), .B(new_n517_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n401_), .A2(new_n482_), .A3(KEYINPUT106), .A4(new_n491_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n544_), .A2(new_n546_), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n580_), .A2(new_n581_), .A3(new_n582_), .A4(new_n583_), .ZN(new_n584_));
  AOI211_X1 g383(.A(new_n242_), .B(new_n315_), .C1(new_n577_), .C2(new_n584_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n274_), .A2(new_n222_), .A3(new_n221_), .A4(new_n275_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(G232gat), .A2(G233gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT34), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n588_), .A2(KEYINPUT35), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n589_), .B1(new_n292_), .B2(new_n209_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(KEYINPUT35), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n591_), .B(KEYINPUT70), .Z(new_n592_));
  AND3_X1   g391(.A1(new_n586_), .A2(new_n590_), .A3(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n592_), .B1(new_n586_), .B2(new_n590_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G190gat), .B(G218gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G134gat), .B(G162gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n598_), .A2(KEYINPUT36), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n595_), .A2(new_n599_), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n598_), .B(KEYINPUT36), .Z(new_n601_));
  OAI21_X1  g400(.A(new_n601_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n603_), .A2(KEYINPUT37), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n600_), .A2(KEYINPUT72), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT72), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n595_), .A2(new_n606_), .A3(new_n599_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n601_), .B(KEYINPUT73), .ZN(new_n608_));
  OAI211_X1 g407(.A(new_n605_), .B(new_n607_), .C1(new_n595_), .C2(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n604_), .B1(new_n609_), .B2(KEYINPUT37), .ZN(new_n610_));
  XOR2_X1   g409(.A(G127gat), .B(G155gat), .Z(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT16), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G183gat), .B(G211gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT17), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n614_), .B(KEYINPUT17), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n215_), .B(new_n293_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(G231gat), .A2(G233gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  MUX2_X1   g419(.A(new_n616_), .B(new_n617_), .S(new_n620_), .Z(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT74), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n610_), .A2(new_n622_), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(KEYINPUT75), .Z(new_n624_));
  AND4_X1   g423(.A1(new_n202_), .A2(new_n585_), .A3(new_n519_), .A4(new_n624_), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n625_), .A2(KEYINPUT38), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(KEYINPUT38), .ZN(new_n627_));
  INV_X1    g426(.A(new_n603_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n628_), .A2(new_n621_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n585_), .A2(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(G1gat), .B1(new_n630_), .B2(new_n581_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n626_), .A2(new_n627_), .A3(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT107), .ZN(G1324gat));
  AND2_X1   g432(.A1(new_n585_), .A2(new_n624_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n634_), .A2(new_n211_), .A3(new_n492_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n492_), .ZN(new_n636_));
  OAI21_X1  g435(.A(G8gat), .B1(new_n630_), .B2(new_n636_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n637_), .A2(KEYINPUT39), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(KEYINPUT39), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n635_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT40), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  OAI211_X1 g441(.A(KEYINPUT40), .B(new_n635_), .C1(new_n638_), .C2(new_n639_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(G1325gat));
  INV_X1    g443(.A(new_n551_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n634_), .A2(new_n528_), .A3(new_n645_), .ZN(new_n646_));
  XOR2_X1   g445(.A(KEYINPUT108), .B(KEYINPUT41), .Z(new_n647_));
  INV_X1    g446(.A(KEYINPUT109), .ZN(new_n648_));
  INV_X1    g447(.A(new_n630_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(new_n645_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n648_), .B1(new_n650_), .B2(G15gat), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  AOI211_X1 g451(.A(KEYINPUT109), .B(new_n528_), .C1(new_n649_), .C2(new_n645_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n647_), .B1(new_n652_), .B2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n647_), .ZN(new_n656_));
  NOR3_X1   g455(.A1(new_n651_), .A2(new_n653_), .A3(new_n656_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n646_), .B1(new_n655_), .B2(new_n657_), .ZN(G1326gat));
  OAI21_X1  g457(.A(G22gat), .B1(new_n630_), .B2(new_n401_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT42), .ZN(new_n660_));
  INV_X1    g459(.A(G22gat), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n634_), .A2(new_n661_), .A3(new_n402_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n662_), .ZN(G1327gat));
  INV_X1    g462(.A(new_n622_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n664_), .A2(new_n603_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n585_), .A2(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(G29gat), .B1(new_n666_), .B2(new_n519_), .ZN(new_n667_));
  OR2_X1    g466(.A1(new_n313_), .A2(new_n314_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n668_), .A2(new_n241_), .A3(new_n622_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT110), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT43), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n671_), .B1(new_n610_), .B2(KEYINPUT111), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n577_), .A2(new_n584_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n673_), .B1(new_n674_), .B2(new_n610_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n610_), .ZN(new_n676_));
  AOI211_X1 g475(.A(new_n676_), .B(new_n672_), .C1(new_n577_), .C2(new_n584_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n670_), .B1(new_n675_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT44), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  OAI211_X1 g479(.A(KEYINPUT44), .B(new_n670_), .C1(new_n675_), .C2(new_n677_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n519_), .A2(G29gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n667_), .B1(new_n682_), .B2(new_n683_), .ZN(G1328gat));
  NAND3_X1  g483(.A1(new_n680_), .A2(new_n492_), .A3(new_n681_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(G36gat), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n636_), .A2(G36gat), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n585_), .A2(new_n665_), .A3(new_n687_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT45), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n686_), .A2(new_n689_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(KEYINPUT112), .B(KEYINPUT46), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n690_), .A2(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n686_), .A2(new_n689_), .A3(new_n691_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(G1329gat));
  NAND4_X1  g494(.A1(new_n680_), .A2(G43gat), .A3(new_n583_), .A4(new_n681_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n666_), .A2(new_n645_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(new_n525_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n698_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g499(.A(G50gat), .B1(new_n666_), .B2(new_n402_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n402_), .A2(G50gat), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n701_), .B1(new_n682_), .B2(new_n702_), .ZN(G1331gat));
  AOI211_X1 g502(.A(new_n241_), .B(new_n668_), .C1(new_n577_), .C2(new_n584_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n622_), .A2(new_n628_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(G57gat), .B1(new_n707_), .B2(new_n581_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n704_), .A2(new_n624_), .ZN(new_n709_));
  INV_X1    g508(.A(G57gat), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n709_), .A2(new_n710_), .A3(new_n519_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n708_), .A2(new_n711_), .ZN(G1332gat));
  INV_X1    g511(.A(G64gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n713_), .B1(new_n706_), .B2(new_n492_), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT48), .Z(new_n715_));
  NAND3_X1  g514(.A1(new_n709_), .A2(new_n713_), .A3(new_n492_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1333gat));
  INV_X1    g516(.A(G71gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n718_), .B1(new_n706_), .B2(new_n645_), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT49), .Z(new_n720_));
  NAND3_X1  g519(.A1(new_n709_), .A2(new_n718_), .A3(new_n645_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1334gat));
  AOI21_X1  g521(.A(new_n371_), .B1(new_n706_), .B2(new_n402_), .ZN(new_n723_));
  XOR2_X1   g522(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n724_));
  XNOR2_X1  g523(.A(new_n723_), .B(new_n724_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n709_), .A2(new_n371_), .A3(new_n402_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1335gat));
  AND2_X1   g526(.A1(new_n704_), .A2(new_n665_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(new_n519_), .ZN(new_n729_));
  INV_X1    g528(.A(G85gat), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  OR2_X1    g530(.A1(new_n731_), .A2(KEYINPUT114), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(KEYINPUT114), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n675_), .A2(new_n677_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n315_), .A2(new_n242_), .A3(new_n622_), .ZN(new_n735_));
  XOR2_X1   g534(.A(new_n735_), .B(KEYINPUT115), .Z(new_n736_));
  AND2_X1   g535(.A1(new_n734_), .A2(new_n736_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n737_), .A2(G85gat), .A3(new_n519_), .ZN(new_n738_));
  AND3_X1   g537(.A1(new_n732_), .A2(new_n733_), .A3(new_n738_), .ZN(G1336gat));
  AOI21_X1  g538(.A(G92gat), .B1(new_n728_), .B2(new_n492_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n492_), .A2(G92gat), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n741_), .B(KEYINPUT116), .Z(new_n742_));
  AOI21_X1  g541(.A(new_n740_), .B1(new_n737_), .B2(new_n742_), .ZN(G1337gat));
  XNOR2_X1  g542(.A(KEYINPUT118), .B(KEYINPUT51), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT117), .ZN(new_n745_));
  OAI211_X1 g544(.A(new_n736_), .B(new_n645_), .C1(new_n675_), .C2(new_n677_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(new_n746_), .B2(G99gat), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n746_), .A2(new_n745_), .A3(G99gat), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n728_), .A2(new_n257_), .A3(new_n583_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n744_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n749_), .ZN(new_n753_));
  OAI211_X1 g552(.A(new_n751_), .B(new_n744_), .C1(new_n753_), .C2(new_n747_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n752_), .A2(new_n755_), .ZN(G1338gat));
  OAI211_X1 g555(.A(new_n736_), .B(new_n402_), .C1(new_n675_), .C2(new_n677_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(G106gat), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT52), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n402_), .A2(new_n258_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n704_), .A2(new_n665_), .A3(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT119), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n762_), .B(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n757_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n760_), .A2(new_n764_), .A3(new_n765_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(KEYINPUT120), .B(KEYINPUT53), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n766_), .B(new_n767_), .ZN(G1339gat));
  NAND3_X1  g567(.A1(new_n623_), .A2(new_n668_), .A3(new_n242_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT54), .ZN(new_n770_));
  INV_X1    g569(.A(new_n293_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT12), .B1(new_n272_), .B2(new_n771_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n772_), .A2(new_n298_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n286_), .B1(new_n773_), .B2(new_n285_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT55), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n296_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n773_), .A2(KEYINPUT55), .A3(new_n286_), .A4(new_n285_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n246_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT56), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n778_), .A2(KEYINPUT56), .A3(new_n779_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n218_), .A2(new_n232_), .A3(new_n224_), .A4(new_n226_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n231_), .A2(new_n219_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n785_), .A2(new_n238_), .A3(new_n786_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n787_), .A2(new_n240_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n784_), .A2(KEYINPUT58), .A3(new_n309_), .A4(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(KEYINPUT56), .B1(new_n778_), .B2(new_n779_), .ZN(new_n790_));
  AOI211_X1 g589(.A(new_n781_), .B(new_n246_), .C1(new_n776_), .C2(new_n777_), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n309_), .B(new_n788_), .C1(new_n790_), .C2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT58), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n789_), .A2(new_n794_), .A3(new_n610_), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n241_), .B(new_n309_), .C1(new_n790_), .C2(new_n791_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT121), .ZN(new_n797_));
  AOI22_X1  g596(.A1(new_n303_), .A2(new_n301_), .B1(new_n306_), .B2(new_n308_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n787_), .A2(new_n240_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n797_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n306_), .A2(new_n308_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n303_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n302_), .B1(new_n296_), .B2(new_n299_), .ZN(new_n803_));
  NOR3_X1   g602(.A1(new_n802_), .A2(new_n803_), .A3(new_n246_), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n788_), .B(KEYINPUT121), .C1(new_n801_), .C2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n796_), .A2(new_n800_), .A3(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT57), .ZN(new_n807_));
  AND3_X1   g606(.A1(new_n806_), .A2(new_n807_), .A3(new_n603_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n807_), .B1(new_n806_), .B2(new_n603_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n795_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n621_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n770_), .A2(new_n811_), .ZN(new_n812_));
  AND4_X1   g611(.A1(new_n519_), .A2(new_n580_), .A3(new_n582_), .A4(new_n583_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(G113gat), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n814_), .A2(new_n815_), .A3(new_n241_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT59), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n814_), .A2(new_n817_), .ZN(new_n818_));
  AND3_X1   g617(.A1(new_n789_), .A2(new_n794_), .A3(new_n610_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n796_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n800_), .A2(new_n805_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n603_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(KEYINPUT57), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n806_), .A2(new_n807_), .A3(new_n603_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n819_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(KEYINPUT122), .B1(new_n825_), .B2(new_n664_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT122), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n810_), .A2(new_n827_), .A3(new_n622_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n826_), .A2(new_n770_), .A3(new_n828_), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n829_), .A2(new_n817_), .A3(new_n813_), .ZN(new_n830_));
  NOR3_X1   g629(.A1(new_n818_), .A2(new_n830_), .A3(new_n242_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n816_), .B1(new_n831_), .B2(new_n815_), .ZN(G1340gat));
  INV_X1    g631(.A(G120gat), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n833_), .B1(new_n668_), .B2(KEYINPUT60), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n814_), .B(new_n834_), .C1(KEYINPUT60), .C2(new_n833_), .ZN(new_n835_));
  NOR3_X1   g634(.A1(new_n818_), .A2(new_n830_), .A3(new_n668_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n835_), .B1(new_n836_), .B2(new_n833_), .ZN(G1341gat));
  INV_X1    g636(.A(G127gat), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n814_), .A2(new_n838_), .A3(new_n664_), .ZN(new_n839_));
  NOR3_X1   g638(.A1(new_n818_), .A2(new_n830_), .A3(new_n621_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n839_), .B1(new_n840_), .B2(new_n838_), .ZN(G1342gat));
  AOI21_X1  g640(.A(G134gat), .B1(new_n814_), .B2(new_n628_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n818_), .A2(new_n830_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(KEYINPUT123), .B(G134gat), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n676_), .A2(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n842_), .B1(new_n843_), .B2(new_n845_), .ZN(G1343gat));
  NOR2_X1   g645(.A1(new_n645_), .A2(new_n401_), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n812_), .A2(new_n847_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n492_), .A2(new_n581_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n850_), .A2(new_n242_), .ZN(new_n851_));
  INV_X1    g650(.A(G141gat), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n851_), .B(new_n852_), .ZN(G1344gat));
  NOR2_X1   g652(.A1(new_n850_), .A2(new_n668_), .ZN(new_n854_));
  INV_X1    g653(.A(G148gat), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n854_), .B(new_n855_), .ZN(G1345gat));
  NAND4_X1  g655(.A1(new_n812_), .A2(new_n664_), .A3(new_n847_), .A4(new_n849_), .ZN(new_n857_));
  OR2_X1    g656(.A1(new_n857_), .A2(KEYINPUT124), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(KEYINPUT124), .ZN(new_n859_));
  XNOR2_X1  g658(.A(KEYINPUT61), .B(G155gat), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n858_), .A2(new_n859_), .A3(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n860_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n861_), .A2(new_n862_), .ZN(G1346gat));
  INV_X1    g662(.A(new_n850_), .ZN(new_n864_));
  AOI21_X1  g663(.A(G162gat), .B1(new_n864_), .B2(new_n628_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n610_), .A2(G162gat), .ZN(new_n866_));
  XOR2_X1   g665(.A(new_n866_), .B(KEYINPUT125), .Z(new_n867_));
  AOI21_X1  g666(.A(new_n865_), .B1(new_n864_), .B2(new_n867_), .ZN(G1347gat));
  NOR4_X1   g667(.A1(new_n551_), .A2(new_n636_), .A3(new_n519_), .A4(new_n402_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n829_), .A2(new_n241_), .A3(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(G169gat), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(KEYINPUT126), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT126), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n870_), .A2(new_n873_), .A3(G169gat), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n872_), .A2(KEYINPUT62), .A3(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT62), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n871_), .A2(KEYINPUT126), .A3(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n829_), .A2(new_n869_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n879_), .A2(new_n241_), .A3(new_n413_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n875_), .A2(new_n877_), .A3(new_n880_), .ZN(G1348gat));
  NAND4_X1  g680(.A1(new_n812_), .A2(G176gat), .A3(new_n315_), .A4(new_n869_), .ZN(new_n882_));
  XOR2_X1   g681(.A(new_n882_), .B(KEYINPUT127), .Z(new_n883_));
  AOI21_X1  g682(.A(G176gat), .B1(new_n879_), .B2(new_n315_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n883_), .A2(new_n884_), .ZN(G1349gat));
  NOR3_X1   g684(.A1(new_n878_), .A2(new_n424_), .A3(new_n621_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n812_), .A2(new_n664_), .A3(new_n869_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n886_), .B1(new_n407_), .B2(new_n887_), .ZN(G1350gat));
  OAI21_X1  g687(.A(G190gat), .B1(new_n878_), .B2(new_n676_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n628_), .A2(new_n425_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n889_), .B1(new_n878_), .B2(new_n890_), .ZN(G1351gat));
  NOR2_X1   g690(.A1(new_n636_), .A2(new_n519_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n848_), .A2(new_n892_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n893_), .A2(new_n242_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(new_n326_), .ZN(G1352gat));
  NAND3_X1  g694(.A1(new_n848_), .A2(new_n315_), .A3(new_n892_), .ZN(new_n896_));
  MUX2_X1   g695(.A(new_n330_), .B(G204gat), .S(new_n896_), .Z(G1353gat));
  NOR2_X1   g696(.A1(new_n893_), .A2(new_n621_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n899_));
  AND2_X1   g698(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n898_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n901_), .B1(new_n898_), .B2(new_n899_), .ZN(G1354gat));
  OAI21_X1  g701(.A(G218gat), .B1(new_n893_), .B2(new_n676_), .ZN(new_n903_));
  OR2_X1    g702(.A1(new_n603_), .A2(G218gat), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n903_), .B1(new_n893_), .B2(new_n904_), .ZN(G1355gat));
endmodule


