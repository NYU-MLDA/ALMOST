//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 0 0 0 1 1 1 1 0 0 1 1 1 1 0 1 1 1 0 0 1 1 1 0 1 1 1 0 0 0 1 0 0 0 1 1 1 1 1 1 1 0 0 1 0 0 1 0 1 0 0 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n623_,
    new_n624_, new_n625_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n691_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n704_, new_n705_, new_n706_, new_n707_, new_n709_,
    new_n710_, new_n711_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n733_, new_n734_, new_n735_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n809_, new_n810_, new_n811_, new_n813_, new_n814_,
    new_n815_, new_n817_, new_n818_, new_n819_, new_n821_, new_n823_,
    new_n824_, new_n826_, new_n827_, new_n828_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n843_, new_n844_,
    new_n845_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n854_, new_n855_, new_n856_, new_n858_, new_n859_,
    new_n860_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_;
  XOR2_X1   g000(.A(G71gat), .B(G78gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G57gat), .B(G64gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT69), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  OAI21_X1  g004(.A(new_n202_), .B1(new_n205_), .B2(KEYINPUT11), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT70), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(KEYINPUT11), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  OR2_X1    g008(.A1(new_n206_), .A2(KEYINPUT70), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n206_), .A2(KEYINPUT70), .ZN(new_n211_));
  NAND4_X1  g010(.A1(new_n210_), .A2(KEYINPUT11), .A3(new_n205_), .A4(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n209_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT12), .ZN(new_n214_));
  INV_X1    g013(.A(G99gat), .ZN(new_n215_));
  INV_X1    g014(.A(G106gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n215_), .A2(new_n216_), .A3(KEYINPUT67), .ZN(new_n217_));
  XOR2_X1   g016(.A(new_n217_), .B(KEYINPUT7), .Z(new_n218_));
  NAND2_X1  g017(.A1(G99gat), .A2(G106gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT6), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  XOR2_X1   g020(.A(G85gat), .B(G92gat), .Z(new_n222_));
  AND2_X1   g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  OR2_X1    g022(.A1(new_n223_), .A2(KEYINPUT8), .ZN(new_n224_));
  OR2_X1    g023(.A1(new_n218_), .A2(KEYINPUT68), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n218_), .A2(KEYINPUT68), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(new_n226_), .A3(new_n220_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n227_), .A2(KEYINPUT8), .A3(new_n222_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT10), .B(G99gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT64), .ZN(new_n230_));
  XNOR2_X1  g029(.A(KEYINPUT65), .B(G106gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT66), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n222_), .A2(KEYINPUT9), .ZN(new_n234_));
  INV_X1    g033(.A(G85gat), .ZN(new_n235_));
  INV_X1    g034(.A(G92gat), .ZN(new_n236_));
  OR3_X1    g035(.A1(new_n235_), .A2(new_n236_), .A3(KEYINPUT9), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n234_), .A2(new_n220_), .A3(new_n237_), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n224_), .B(new_n228_), .C1(new_n233_), .C2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n213_), .A2(new_n214_), .A3(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n213_), .B(new_n239_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n240_), .B1(new_n241_), .B2(new_n214_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G230gat), .A2(G233gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n241_), .A2(G230gat), .A3(G233gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G120gat), .B(G148gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT5), .ZN(new_n247_));
  XOR2_X1   g046(.A(G176gat), .B(G204gat), .Z(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n244_), .A2(new_n245_), .A3(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT72), .ZN(new_n252_));
  OR2_X1    g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n252_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n244_), .A2(new_n245_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n250_), .B1(new_n256_), .B2(KEYINPUT71), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n257_), .B1(KEYINPUT71), .B2(new_n256_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n255_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT13), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n255_), .A2(new_n258_), .A3(KEYINPUT13), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT73), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G29gat), .B(G36gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT75), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G43gat), .B(G50gat), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  OR2_X1    g067(.A1(new_n266_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n266_), .A2(new_n268_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT82), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(KEYINPUT81), .B(G8gat), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(G1gat), .ZN(new_n276_));
  OAI21_X1  g075(.A(KEYINPUT14), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G15gat), .B(G22gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G1gat), .B(G8gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n273_), .B(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G229gat), .A2(G233gat), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT83), .ZN(new_n287_));
  XOR2_X1   g086(.A(new_n271_), .B(KEYINPUT15), .Z(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(new_n281_), .ZN(new_n289_));
  XOR2_X1   g088(.A(new_n289_), .B(KEYINPUT84), .Z(new_n290_));
  NAND2_X1  g089(.A1(new_n273_), .A2(new_n282_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n290_), .A2(new_n291_), .A3(new_n284_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n287_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G113gat), .B(G141gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G169gat), .B(G197gat), .ZN(new_n295_));
  XOR2_X1   g094(.A(new_n294_), .B(new_n295_), .Z(new_n296_));
  XNOR2_X1  g095(.A(new_n293_), .B(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT97), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G78gat), .B(G106gat), .ZN(new_n299_));
  INV_X1    g098(.A(G228gat), .ZN(new_n300_));
  INV_X1    g099(.A(G233gat), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  XOR2_X1   g102(.A(G211gat), .B(G218gat), .Z(new_n304_));
  INV_X1    g103(.A(G197gat), .ZN(new_n305_));
  INV_X1    g104(.A(G204gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  AND2_X1   g106(.A1(KEYINPUT92), .A2(G204gat), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(KEYINPUT92), .A2(G204gat), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n307_), .B1(new_n313_), .B2(new_n305_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT21), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n304_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n305_), .B1(new_n308_), .B2(new_n310_), .ZN(new_n317_));
  AOI22_X1  g116(.A1(new_n317_), .A2(KEYINPUT93), .B1(G197gat), .B2(new_n306_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT93), .ZN(new_n319_));
  OAI211_X1 g118(.A(new_n319_), .B(new_n305_), .C1(new_n308_), .C2(new_n310_), .ZN(new_n320_));
  AOI211_X1 g119(.A(KEYINPUT94), .B(new_n315_), .C1(new_n318_), .C2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT94), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n317_), .A2(KEYINPUT93), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n306_), .A2(G197gat), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n323_), .A2(new_n320_), .A3(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n322_), .B1(new_n325_), .B2(KEYINPUT21), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n316_), .B1(new_n321_), .B2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT95), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT95), .ZN(new_n329_));
  OAI211_X1 g128(.A(new_n329_), .B(new_n316_), .C1(new_n321_), .C2(new_n326_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n304_), .ZN(new_n332_));
  NOR3_X1   g131(.A1(new_n314_), .A2(new_n315_), .A3(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n331_), .A2(new_n334_), .ZN(new_n335_));
  OR2_X1    g134(.A1(G155gat), .A2(G162gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G155gat), .A2(G162gat), .ZN(new_n337_));
  OR2_X1    g136(.A1(G141gat), .A2(G148gat), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT3), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT91), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n338_), .B(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G141gat), .A2(G148gat), .ZN(new_n342_));
  XOR2_X1   g141(.A(new_n342_), .B(KEYINPUT2), .Z(new_n343_));
  OAI211_X1 g142(.A(new_n336_), .B(new_n337_), .C1(new_n341_), .C2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n337_), .A2(KEYINPUT1), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(new_n336_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n337_), .A2(KEYINPUT1), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n338_), .B(new_n342_), .C1(new_n346_), .C2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n344_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT29), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n303_), .B1(new_n335_), .B2(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n333_), .B1(new_n328_), .B2(new_n330_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n350_), .ZN(new_n353_));
  NOR3_X1   g152(.A1(new_n352_), .A2(new_n302_), .A3(new_n353_), .ZN(new_n354_));
  OAI211_X1 g153(.A(new_n298_), .B(new_n299_), .C1(new_n351_), .C2(new_n354_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n349_), .A2(KEYINPUT29), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(KEYINPUT28), .ZN(new_n357_));
  XOR2_X1   g156(.A(G22gat), .B(G50gat), .Z(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n335_), .A2(new_n303_), .A3(new_n350_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n302_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n299_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n360_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n355_), .A2(new_n359_), .A3(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n360_), .A2(new_n361_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n298_), .B1(new_n365_), .B2(new_n299_), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT98), .B1(new_n364_), .B2(new_n366_), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n363_), .A2(new_n359_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n299_), .B1(new_n351_), .B2(new_n354_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT97), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT98), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n368_), .A2(new_n370_), .A3(new_n371_), .A4(new_n355_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n359_), .B1(new_n369_), .B2(new_n363_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT96), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  AOI211_X1 g174(.A(KEYINPUT96), .B(new_n359_), .C1(new_n369_), .C2(new_n363_), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n367_), .B(new_n372_), .C1(new_n375_), .C2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G1gat), .B(G29gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(G85gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(KEYINPUT0), .B(G57gat), .ZN(new_n381_));
  XOR2_X1   g180(.A(new_n380_), .B(new_n381_), .Z(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G127gat), .B(G134gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G113gat), .B(G120gat), .ZN(new_n385_));
  OR2_X1    g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(new_n385_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n386_), .A2(KEYINPUT90), .A3(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT90), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n384_), .A2(new_n385_), .A3(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n349_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n386_), .A2(new_n387_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n344_), .A2(new_n348_), .A3(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n392_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT4), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT101), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT101), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n392_), .A2(new_n398_), .A3(KEYINPUT4), .A4(new_n394_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n349_), .A2(new_n396_), .A3(new_n391_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n397_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G225gat), .A2(G233gat), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n395_), .A2(new_n402_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n383_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n405_), .ZN(new_n407_));
  AOI211_X1 g206(.A(new_n382_), .B(new_n407_), .C1(new_n401_), .C2(new_n403_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n406_), .A2(new_n408_), .ZN(new_n409_));
  XOR2_X1   g208(.A(new_n409_), .B(KEYINPUT105), .Z(new_n410_));
  INV_X1    g209(.A(G169gat), .ZN(new_n411_));
  INV_X1    g210(.A(G176gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n413_), .A2(KEYINPUT24), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G183gat), .A2(G190gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(KEYINPUT23), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT23), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n417_), .A2(G183gat), .A3(G190gat), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n414_), .B1(new_n416_), .B2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT85), .ZN(new_n420_));
  OR2_X1    g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT25), .B(G183gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT26), .B(G190gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G169gat), .A2(G176gat), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n424_), .A2(KEYINPUT24), .ZN(new_n425_));
  AOI22_X1  g224(.A1(new_n422_), .A2(new_n423_), .B1(new_n425_), .B2(new_n413_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n419_), .A2(new_n420_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n421_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n415_), .A2(new_n417_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n430_));
  OAI211_X1 g229(.A(new_n429_), .B(new_n430_), .C1(G183gat), .C2(G190gat), .ZN(new_n431_));
  OR2_X1    g230(.A1(new_n431_), .A2(KEYINPUT88), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(KEYINPUT88), .ZN(new_n433_));
  XOR2_X1   g232(.A(KEYINPUT87), .B(G176gat), .Z(new_n434_));
  INV_X1    g233(.A(KEYINPUT86), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT22), .ZN(new_n436_));
  OAI21_X1  g235(.A(G169gat), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n411_), .A2(KEYINPUT22), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n434_), .B(new_n437_), .C1(new_n435_), .C2(new_n438_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n432_), .A2(new_n424_), .A3(new_n433_), .A4(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n428_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G227gat), .A2(G233gat), .ZN(new_n442_));
  INV_X1    g241(.A(G71gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(G99gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n441_), .B(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(new_n391_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G15gat), .B(G43gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(KEYINPUT89), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(KEYINPUT30), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(KEYINPUT31), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n447_), .B(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n410_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT106), .ZN(new_n455_));
  INV_X1    g254(.A(new_n441_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n325_), .A2(KEYINPUT21), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT94), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n325_), .A2(new_n322_), .A3(KEYINPUT21), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n329_), .B1(new_n460_), .B2(new_n316_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n330_), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n334_), .B(new_n456_), .C1(new_n461_), .C2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT20), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G226gat), .A2(G233gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(KEYINPUT19), .ZN(new_n466_));
  XOR2_X1   g265(.A(new_n466_), .B(KEYINPUT99), .Z(new_n467_));
  NAND2_X1  g266(.A1(new_n436_), .A2(G169gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n438_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(new_n434_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n471_), .A2(new_n424_), .A3(new_n431_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n419_), .A2(new_n426_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n475_), .B1(new_n331_), .B2(new_n334_), .ZN(new_n476_));
  NOR3_X1   g275(.A1(new_n464_), .A2(new_n467_), .A3(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT103), .ZN(new_n478_));
  AOI211_X1 g277(.A(new_n333_), .B(new_n474_), .C1(new_n328_), .C2(new_n330_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT20), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n478_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n335_), .A2(new_n441_), .ZN(new_n482_));
  OAI211_X1 g281(.A(new_n334_), .B(new_n475_), .C1(new_n461_), .C2(new_n462_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n483_), .A2(KEYINPUT103), .A3(KEYINPUT20), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n481_), .A2(new_n482_), .A3(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n477_), .B1(new_n485_), .B2(new_n466_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G8gat), .B(G36gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(KEYINPUT18), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G64gat), .B(G92gat), .ZN(new_n489_));
  XOR2_X1   g288(.A(new_n488_), .B(new_n489_), .Z(new_n490_));
  OAI21_X1  g289(.A(new_n455_), .B1(new_n486_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n490_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n466_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n483_), .A2(KEYINPUT20), .ZN(new_n494_));
  AOI22_X1  g293(.A1(new_n494_), .A2(new_n478_), .B1(new_n335_), .B2(new_n441_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n493_), .B1(new_n495_), .B2(new_n484_), .ZN(new_n496_));
  OAI211_X1 g295(.A(KEYINPUT106), .B(new_n492_), .C1(new_n496_), .C2(new_n477_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n467_), .B1(new_n464_), .B2(new_n476_), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n482_), .A2(KEYINPUT20), .A3(new_n493_), .A4(new_n483_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n498_), .A2(new_n499_), .A3(new_n490_), .ZN(new_n500_));
  AND2_X1   g299(.A1(new_n500_), .A2(KEYINPUT27), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n491_), .A2(new_n497_), .A3(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT107), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT107), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n491_), .A2(new_n497_), .A3(new_n504_), .A4(new_n501_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n503_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n467_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n476_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n480_), .B1(new_n352_), .B2(new_n456_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n507_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n493_), .B1(new_n352_), .B2(new_n456_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n494_), .A2(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n492_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n513_), .A2(KEYINPUT100), .A3(new_n500_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT100), .ZN(new_n515_));
  OAI211_X1 g314(.A(new_n515_), .B(new_n492_), .C1(new_n510_), .C2(new_n512_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n514_), .A2(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n517_), .A2(KEYINPUT27), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(KEYINPUT108), .B1(new_n506_), .B2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT108), .ZN(new_n521_));
  AOI211_X1 g320(.A(new_n521_), .B(new_n518_), .C1(new_n503_), .C2(new_n505_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n378_), .B(new_n454_), .C1(new_n520_), .C2(new_n522_), .ZN(new_n523_));
  AND2_X1   g322(.A1(new_n367_), .A2(new_n372_), .ZN(new_n524_));
  OR2_X1    g323(.A1(new_n375_), .A2(new_n376_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n410_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  AND3_X1   g325(.A1(new_n506_), .A2(new_n519_), .A3(new_n526_), .ZN(new_n527_));
  OR2_X1    g326(.A1(new_n406_), .A2(KEYINPUT33), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n406_), .A2(KEYINPUT33), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n383_), .B1(new_n395_), .B2(new_n402_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT102), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n531_), .B1(new_n403_), .B2(new_n401_), .ZN(new_n532_));
  AND3_X1   g331(.A1(new_n528_), .A2(new_n529_), .A3(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n517_), .A2(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n510_), .A2(new_n512_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n490_), .A2(KEYINPUT32), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n409_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  OAI211_X1 g336(.A(KEYINPUT32), .B(new_n490_), .C1(new_n496_), .C2(new_n477_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n534_), .A2(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n540_), .A2(new_n378_), .A3(KEYINPUT104), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT104), .ZN(new_n542_));
  AOI22_X1  g341(.A1(new_n517_), .A2(new_n533_), .B1(new_n538_), .B2(new_n537_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n542_), .B1(new_n543_), .B2(new_n377_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n541_), .A2(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n453_), .B1(new_n527_), .B2(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n297_), .B1(new_n523_), .B2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G190gat), .B(G218gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT76), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G134gat), .B(G162gat), .ZN(new_n550_));
  XOR2_X1   g349(.A(new_n549_), .B(new_n550_), .Z(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT36), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT78), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n239_), .A2(new_n288_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT77), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G232gat), .A2(G233gat), .ZN(new_n556_));
  XOR2_X1   g355(.A(new_n556_), .B(KEYINPUT34), .Z(new_n557_));
  XOR2_X1   g356(.A(KEYINPUT74), .B(KEYINPUT35), .Z(new_n558_));
  AOI21_X1  g357(.A(new_n555_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  OAI211_X1 g358(.A(new_n554_), .B(new_n559_), .C1(new_n271_), .C2(new_n239_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n557_), .A2(new_n558_), .ZN(new_n561_));
  OR2_X1    g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n560_), .A2(new_n561_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n553_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT36), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n562_), .A2(new_n566_), .A3(new_n563_), .A4(new_n551_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  XOR2_X1   g368(.A(KEYINPUT80), .B(KEYINPUT37), .Z(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n565_), .A2(KEYINPUT79), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT79), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n567_), .B1(new_n564_), .B2(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(KEYINPUT37), .B1(new_n572_), .B2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n571_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G231gat), .A2(G233gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n213_), .B(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(new_n282_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G127gat), .B(G155gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT16), .ZN(new_n582_));
  XOR2_X1   g381(.A(G183gat), .B(G211gat), .Z(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(KEYINPUT17), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n585_), .A2(KEYINPUT17), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n580_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n580_), .A2(new_n586_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n577_), .A2(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n264_), .A2(new_n547_), .A3(new_n592_), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n410_), .A2(KEYINPUT109), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n410_), .A2(KEYINPUT109), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  OR3_X1    g396(.A1(new_n593_), .A2(G1gat), .A3(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT38), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n569_), .B1(new_n523_), .B2(new_n546_), .ZN(new_n601_));
  NOR3_X1   g400(.A1(new_n263_), .A2(new_n297_), .A3(new_n591_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n410_), .ZN(new_n604_));
  OAI21_X1  g403(.A(G1gat), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n598_), .A2(new_n599_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n600_), .A2(new_n605_), .A3(new_n606_), .ZN(G1324gat));
  NOR2_X1   g406(.A1(new_n520_), .A2(new_n522_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(new_n275_), .ZN(new_n609_));
  OR3_X1    g408(.A1(new_n593_), .A2(KEYINPUT110), .A3(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(KEYINPUT110), .B1(new_n593_), .B2(new_n609_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n608_), .ZN(new_n613_));
  OAI21_X1  g412(.A(G8gat), .B1(new_n603_), .B2(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(KEYINPUT111), .B(KEYINPUT39), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  OR2_X1    g415(.A1(new_n614_), .A2(new_n615_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n612_), .A2(new_n616_), .A3(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT40), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n612_), .A2(KEYINPUT40), .A3(new_n616_), .A4(new_n617_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(G1325gat));
  OAI21_X1  g421(.A(G15gat), .B1(new_n603_), .B2(new_n453_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT41), .ZN(new_n624_));
  NOR3_X1   g423(.A1(new_n593_), .A2(G15gat), .A3(new_n453_), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n624_), .A2(new_n625_), .ZN(G1326gat));
  NAND3_X1  g425(.A1(new_n601_), .A2(new_n602_), .A3(new_n377_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(KEYINPUT112), .B(KEYINPUT42), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n627_), .A2(G22gat), .A3(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n628_), .B1(new_n627_), .B2(G22gat), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n378_), .A2(G22gat), .ZN(new_n631_));
  OAI22_X1  g430(.A1(new_n629_), .A2(new_n630_), .B1(new_n593_), .B2(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT113), .ZN(G1327gat));
  NAND2_X1  g432(.A1(new_n596_), .A2(G29gat), .ZN(new_n634_));
  NOR3_X1   g433(.A1(new_n263_), .A2(new_n297_), .A3(new_n590_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT43), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n523_), .A2(new_n546_), .ZN(new_n637_));
  AND3_X1   g436(.A1(new_n571_), .A2(new_n575_), .A3(KEYINPUT114), .ZN(new_n638_));
  AOI21_X1  g437(.A(KEYINPUT114), .B1(new_n571_), .B2(new_n575_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n636_), .B1(new_n637_), .B2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n577_), .A2(new_n636_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n642_), .B1(new_n523_), .B2(new_n546_), .ZN(new_n643_));
  OAI211_X1 g442(.A(KEYINPUT44), .B(new_n635_), .C1(new_n641_), .C2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n635_), .B1(new_n641_), .B2(new_n643_), .ZN(new_n646_));
  AOI21_X1  g445(.A(KEYINPUT44), .B1(new_n646_), .B2(KEYINPUT115), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT115), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n648_), .B(new_n635_), .C1(new_n641_), .C2(new_n643_), .ZN(new_n649_));
  AOI211_X1 g448(.A(new_n634_), .B(new_n645_), .C1(new_n647_), .C2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n591_), .A2(new_n569_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n263_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n547_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(KEYINPUT116), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT116), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n547_), .A2(new_n655_), .A3(new_n652_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n654_), .A2(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(G29gat), .B1(new_n657_), .B2(new_n410_), .ZN(new_n658_));
  OAI21_X1  g457(.A(KEYINPUT117), .B1(new_n650_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n658_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT117), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n646_), .A2(KEYINPUT115), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT44), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n662_), .A2(new_n663_), .A3(new_n649_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(new_n644_), .ZN(new_n665_));
  OAI211_X1 g464(.A(new_n660_), .B(new_n661_), .C1(new_n665_), .C2(new_n634_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n659_), .A2(new_n666_), .ZN(G1328gat));
  INV_X1    g466(.A(KEYINPUT46), .ZN(new_n668_));
  INV_X1    g467(.A(G36gat), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n644_), .A2(new_n608_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n669_), .B1(new_n664_), .B2(new_n671_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n654_), .A2(new_n608_), .A3(new_n669_), .A4(new_n656_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT45), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n673_), .B(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n668_), .B1(new_n672_), .B2(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n673_), .B(KEYINPUT45), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n670_), .B1(new_n647_), .B2(new_n649_), .ZN(new_n678_));
  OAI211_X1 g477(.A(new_n677_), .B(KEYINPUT46), .C1(new_n669_), .C2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n676_), .A2(new_n679_), .ZN(G1329gat));
  NAND2_X1  g479(.A1(new_n452_), .A2(G43gat), .ZN(new_n681_));
  AOI211_X1 g480(.A(new_n681_), .B(new_n645_), .C1(new_n647_), .C2(new_n649_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n657_), .A2(new_n452_), .ZN(new_n683_));
  XOR2_X1   g482(.A(KEYINPUT118), .B(G43gat), .Z(new_n684_));
  AND2_X1   g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(KEYINPUT47), .B1(new_n682_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT47), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n683_), .A2(new_n684_), .ZN(new_n688_));
  OAI211_X1 g487(.A(new_n687_), .B(new_n688_), .C1(new_n665_), .C2(new_n681_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n686_), .A2(new_n689_), .ZN(G1330gat));
  AOI21_X1  g489(.A(G50gat), .B1(new_n657_), .B2(new_n377_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n665_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n377_), .A2(G50gat), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n691_), .B1(new_n692_), .B2(new_n693_), .ZN(G1331gat));
  INV_X1    g493(.A(new_n264_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n297_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n696_), .A2(new_n591_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n695_), .A2(new_n601_), .A3(new_n697_), .ZN(new_n698_));
  OAI21_X1  g497(.A(G57gat), .B1(new_n698_), .B2(new_n604_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n696_), .B1(new_n523_), .B2(new_n546_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n700_), .A2(new_n263_), .A3(new_n592_), .ZN(new_n701_));
  OR2_X1    g500(.A1(new_n597_), .A2(G57gat), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n699_), .B1(new_n701_), .B2(new_n702_), .ZN(G1332gat));
  OAI21_X1  g502(.A(G64gat), .B1(new_n698_), .B2(new_n613_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT48), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n613_), .A2(G64gat), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT119), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n705_), .B1(new_n701_), .B2(new_n707_), .ZN(G1333gat));
  OAI21_X1  g507(.A(G71gat), .B1(new_n698_), .B2(new_n453_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT49), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n452_), .A2(new_n443_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n710_), .B1(new_n701_), .B2(new_n711_), .ZN(G1334gat));
  OR3_X1    g511(.A1(new_n701_), .A2(G78gat), .A3(new_n378_), .ZN(new_n713_));
  OR2_X1    g512(.A1(new_n698_), .A2(new_n378_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(KEYINPUT120), .B(KEYINPUT50), .ZN(new_n715_));
  AND3_X1   g514(.A1(new_n714_), .A2(G78gat), .A3(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n715_), .B1(new_n714_), .B2(G78gat), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n713_), .B1(new_n716_), .B2(new_n717_), .ZN(G1335gat));
  NOR2_X1   g517(.A1(new_n641_), .A2(new_n643_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n263_), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n720_), .A2(new_n696_), .A3(new_n590_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n719_), .A2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(new_n410_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(G85gat), .ZN(new_n725_));
  AND4_X1   g524(.A1(new_n695_), .A2(new_n591_), .A3(new_n569_), .A4(new_n700_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n726_), .A2(new_n235_), .A3(new_n596_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(KEYINPUT121), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT121), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n725_), .A2(new_n730_), .A3(new_n727_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(G1336gat));
  NAND3_X1  g531(.A1(new_n726_), .A2(new_n236_), .A3(new_n608_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n723_), .A2(new_n608_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n733_), .B1(new_n735_), .B2(new_n236_), .ZN(G1337gat));
  NAND2_X1  g535(.A1(new_n723_), .A2(new_n452_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(G99gat), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n726_), .A2(new_n452_), .A3(new_n230_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT51), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT51), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n738_), .A2(new_n742_), .A3(new_n739_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(G1338gat));
  NAND3_X1  g543(.A1(new_n726_), .A2(new_n377_), .A3(new_n231_), .ZN(new_n745_));
  OAI211_X1 g544(.A(new_n377_), .B(new_n721_), .C1(new_n641_), .C2(new_n643_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT52), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n746_), .A2(new_n747_), .A3(G106gat), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n746_), .B2(G106gat), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n745_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g550(.A1(new_n597_), .A2(new_n453_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT57), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n290_), .A2(new_n291_), .A3(new_n285_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n296_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n296_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n757_), .B1(new_n293_), .B2(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n759_), .B1(new_n255_), .B2(new_n258_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n242_), .A2(KEYINPUT55), .ZN(new_n761_));
  NAND3_X1  g560(.A1(KEYINPUT122), .A2(G230gat), .A3(G233gat), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n763_), .A2(new_n250_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n242_), .A2(new_n243_), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n761_), .B(new_n762_), .C1(new_n765_), .C2(KEYINPUT55), .ZN(new_n766_));
  AOI21_X1  g565(.A(KEYINPUT56), .B1(new_n764_), .B2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n764_), .A2(new_n766_), .A3(KEYINPUT56), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n297_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n760_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n754_), .B1(new_n772_), .B2(new_n569_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n255_), .A2(new_n696_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n774_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n775_));
  OAI211_X1 g574(.A(KEYINPUT57), .B(new_n568_), .C1(new_n775_), .C2(new_n760_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n759_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n770_), .A2(KEYINPUT58), .A3(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n769_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n777_), .B1(new_n779_), .B2(new_n767_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT58), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n778_), .A2(new_n782_), .A3(new_n577_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n773_), .A2(new_n776_), .A3(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(new_n591_), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n261_), .A2(new_n576_), .A3(new_n262_), .A4(new_n697_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT54), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n753_), .B1(new_n785_), .B2(new_n787_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n608_), .A2(new_n377_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(G113gat), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n790_), .A2(new_n791_), .A3(new_n696_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n785_), .A2(new_n787_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT123), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n793_), .A2(new_n794_), .A3(new_n789_), .A4(new_n752_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT59), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n788_), .A2(new_n794_), .A3(KEYINPUT59), .A4(new_n789_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n297_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n792_), .B1(new_n799_), .B2(new_n791_), .ZN(G1340gat));
  NOR2_X1   g599(.A1(new_n720_), .A2(KEYINPUT60), .ZN(new_n801_));
  INV_X1    g600(.A(G120gat), .ZN(new_n802_));
  MUX2_X1   g601(.A(KEYINPUT60), .B(new_n801_), .S(new_n802_), .Z(new_n803_));
  NAND4_X1  g602(.A1(new_n793_), .A2(new_n789_), .A3(new_n752_), .A4(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT124), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n804_), .B(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n264_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n806_), .B1(new_n807_), .B2(new_n802_), .ZN(G1341gat));
  INV_X1    g607(.A(G127gat), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n790_), .A2(new_n809_), .A3(new_n590_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n591_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n810_), .B1(new_n811_), .B2(new_n809_), .ZN(G1342gat));
  INV_X1    g611(.A(G134gat), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n790_), .A2(new_n813_), .A3(new_n569_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n576_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n814_), .B1(new_n815_), .B2(new_n813_), .ZN(G1343gat));
  NAND3_X1  g615(.A1(new_n596_), .A2(new_n377_), .A3(new_n453_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n817_), .B1(new_n785_), .B2(new_n787_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n818_), .A2(new_n613_), .A3(new_n696_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n819_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g619(.A1(new_n818_), .A2(new_n613_), .A3(new_n695_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g621(.A1(new_n818_), .A2(new_n613_), .A3(new_n590_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(KEYINPUT61), .B(G155gat), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n823_), .B(new_n824_), .ZN(G1346gat));
  AND2_X1   g624(.A1(new_n818_), .A2(new_n613_), .ZN(new_n826_));
  AOI21_X1  g625(.A(G162gat), .B1(new_n826_), .B2(new_n569_), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n640_), .A2(G162gat), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n827_), .B1(new_n826_), .B2(new_n828_), .ZN(G1347gat));
  NOR3_X1   g628(.A1(new_n596_), .A2(new_n377_), .A3(new_n453_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n831_), .B1(new_n785_), .B2(new_n787_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n832_), .A2(KEYINPUT125), .A3(new_n608_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(KEYINPUT125), .B1(new_n832_), .B2(new_n608_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n696_), .A2(new_n470_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n832_), .A2(new_n608_), .A3(new_n696_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT62), .ZN(new_n839_));
  AND3_X1   g638(.A1(new_n838_), .A2(new_n839_), .A3(G169gat), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n839_), .B1(new_n838_), .B2(G169gat), .ZN(new_n841_));
  OAI22_X1  g640(.A1(new_n836_), .A2(new_n837_), .B1(new_n840_), .B2(new_n841_), .ZN(G1348gat));
  NAND3_X1  g641(.A1(new_n793_), .A2(new_n608_), .A3(new_n830_), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n843_), .A2(new_n412_), .A3(new_n264_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n263_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n844_), .B1(new_n845_), .B2(new_n434_), .ZN(G1349gat));
  NOR2_X1   g645(.A1(new_n843_), .A2(new_n591_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n847_), .A2(G183gat), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT125), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n843_), .A2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n833_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n591_), .A2(new_n422_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n848_), .B1(new_n851_), .B2(new_n852_), .ZN(G1350gat));
  OAI211_X1 g652(.A(new_n423_), .B(new_n569_), .C1(new_n834_), .C2(new_n835_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n576_), .B1(new_n850_), .B2(new_n833_), .ZN(new_n855_));
  INV_X1    g654(.A(G190gat), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n854_), .B1(new_n855_), .B2(new_n856_), .ZN(G1351gat));
  NAND2_X1  g656(.A1(new_n526_), .A2(new_n453_), .ZN(new_n858_));
  AOI211_X1 g657(.A(new_n613_), .B(new_n858_), .C1(new_n785_), .C2(new_n787_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n696_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g660(.A(new_n858_), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n793_), .A2(new_n608_), .A3(new_n695_), .A4(new_n862_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n863_), .A2(new_n312_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT127), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n863_), .A2(KEYINPUT127), .A3(new_n312_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n863_), .A2(KEYINPUT126), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(G204gat), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n863_), .A2(KEYINPUT126), .ZN(new_n870_));
  OAI22_X1  g669(.A1(new_n866_), .A2(new_n867_), .B1(new_n869_), .B2(new_n870_), .ZN(G1353gat));
  AOI211_X1 g670(.A(KEYINPUT63), .B(G211gat), .C1(new_n859_), .C2(new_n590_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n859_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n873_), .A2(new_n591_), .ZN(new_n874_));
  XOR2_X1   g673(.A(KEYINPUT63), .B(G211gat), .Z(new_n875_));
  AOI21_X1  g674(.A(new_n872_), .B1(new_n874_), .B2(new_n875_), .ZN(G1354gat));
  OAI21_X1  g675(.A(G218gat), .B1(new_n873_), .B2(new_n576_), .ZN(new_n877_));
  OR2_X1    g676(.A1(new_n568_), .A2(G218gat), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n873_), .B2(new_n878_), .ZN(G1355gat));
endmodule


