//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 1 0 1 1 0 1 1 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 0 1 0 0 1 0 0 0 1 0 1 0 0 1 1 1 1 1 1 1 1 1 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n674_, new_n675_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n698_, new_n699_, new_n700_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n718_, new_n719_,
    new_n720_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n824_, new_n825_, new_n826_,
    new_n828_, new_n829_, new_n830_, new_n832_, new_n833_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n865_, new_n866_, new_n867_, new_n869_, new_n870_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n896_;
  INV_X1    g000(.A(KEYINPUT98), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G141gat), .A2(G148gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  NOR2_X1   g003(.A1(G141gat), .A2(G148gat), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT82), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT82), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n210_), .A2(G155gat), .A3(G162gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n212_), .A2(KEYINPUT1), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n214_), .B1(new_n212_), .B2(KEYINPUT1), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT83), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n213_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT1), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n218_), .B1(new_n209_), .B2(new_n211_), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT83), .B1(new_n219_), .B2(new_n214_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n207_), .B1(new_n217_), .B2(new_n220_), .ZN(new_n221_));
  AND2_X1   g020(.A1(new_n209_), .A2(new_n211_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT3), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT2), .ZN(new_n224_));
  OAI22_X1  g023(.A1(new_n205_), .A2(new_n223_), .B1(new_n203_), .B2(new_n224_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n225_), .B1(new_n223_), .B2(new_n205_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n203_), .A2(new_n224_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(KEYINPUT84), .ZN(new_n228_));
  AOI211_X1 g027(.A(new_n214_), .B(new_n222_), .C1(new_n226_), .C2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT85), .B1(new_n221_), .B2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n214_), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n216_), .B(new_n231_), .C1(new_n222_), .C2(new_n218_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n213_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n232_), .A2(new_n220_), .A3(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(new_n206_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT85), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n226_), .A2(new_n228_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n237_), .A2(new_n231_), .A3(new_n212_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n235_), .A2(new_n236_), .A3(new_n238_), .ZN(new_n239_));
  XOR2_X1   g038(.A(G127gat), .B(G134gat), .Z(new_n240_));
  XNOR2_X1  g039(.A(G113gat), .B(G120gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n230_), .A2(new_n239_), .A3(new_n242_), .ZN(new_n243_));
  OR3_X1    g042(.A1(new_n221_), .A2(new_n229_), .A3(new_n242_), .ZN(new_n244_));
  AND3_X1   g043(.A1(new_n243_), .A2(KEYINPUT4), .A3(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT4), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n230_), .A2(new_n239_), .A3(new_n246_), .A4(new_n242_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G225gat), .A2(G233gat), .ZN(new_n248_));
  XOR2_X1   g047(.A(new_n248_), .B(KEYINPUT91), .Z(new_n249_));
  NAND2_X1  g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(KEYINPUT92), .B1(new_n245_), .B2(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n243_), .A2(KEYINPUT4), .A3(new_n244_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT92), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n252_), .A2(new_n253_), .A3(new_n249_), .A4(new_n247_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n249_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n243_), .A2(new_n244_), .A3(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n251_), .A2(new_n254_), .A3(new_n256_), .ZN(new_n257_));
  XOR2_X1   g056(.A(G57gat), .B(G85gat), .Z(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT94), .ZN(new_n259_));
  XOR2_X1   g058(.A(G1gat), .B(G29gat), .Z(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n262_));
  XOR2_X1   g061(.A(new_n261_), .B(new_n262_), .Z(new_n263_));
  NAND2_X1  g062(.A1(new_n257_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n263_), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n251_), .A2(new_n265_), .A3(new_n254_), .A4(new_n256_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT86), .ZN(new_n269_));
  INV_X1    g068(.A(G218gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(G211gat), .ZN(new_n271_));
  INV_X1    g070(.A(G211gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(G218gat), .ZN(new_n273_));
  AND3_X1   g072(.A1(new_n271_), .A2(new_n273_), .A3(KEYINPUT87), .ZN(new_n274_));
  AOI21_X1  g073(.A(KEYINPUT87), .B1(new_n271_), .B2(new_n273_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n269_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT21), .ZN(new_n277_));
  AND2_X1   g076(.A1(G197gat), .A2(G204gat), .ZN(new_n278_));
  NOR2_X1   g077(.A1(G197gat), .A2(G204gat), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n277_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n280_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n281_));
  NOR3_X1   g080(.A1(new_n278_), .A2(new_n279_), .A3(new_n277_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n276_), .A2(new_n281_), .A3(new_n283_), .ZN(new_n284_));
  OAI221_X1 g083(.A(new_n280_), .B1(new_n282_), .B2(new_n269_), .C1(new_n274_), .C2(new_n275_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n286_), .B1(G228gat), .B2(G233gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n230_), .A2(new_n239_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT29), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n287_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n289_), .B1(new_n235_), .B2(new_n238_), .ZN(new_n291_));
  OAI211_X1 g090(.A(G228gat), .B(G233gat), .C1(new_n291_), .C2(new_n286_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  XOR2_X1   g092(.A(G78gat), .B(G106gat), .Z(new_n294_));
  OR2_X1    g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n293_), .A2(new_n294_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G22gat), .B(G50gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n288_), .A2(new_n289_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT28), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n299_), .A2(KEYINPUT28), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n298_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n302_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n298_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n304_), .A2(new_n300_), .A3(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n303_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n297_), .A2(new_n307_), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n306_), .A2(new_n303_), .A3(new_n295_), .A4(new_n296_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n268_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G8gat), .B(G36gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT18), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G64gat), .B(G92gat), .ZN(new_n314_));
  XOR2_X1   g113(.A(new_n313_), .B(new_n314_), .Z(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT90), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT89), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT23), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n319_), .B1(G183gat), .B2(G190gat), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(G183gat), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n322_), .A2(KEYINPUT23), .ZN(new_n323_));
  AOI21_X1  g122(.A(KEYINPUT78), .B1(new_n323_), .B2(G190gat), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n319_), .A2(KEYINPUT78), .A3(G183gat), .A4(G190gat), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n321_), .B1(new_n324_), .B2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT88), .ZN(new_n328_));
  NOR2_X1   g127(.A1(G183gat), .A2(G190gat), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n327_), .A2(new_n328_), .A3(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n319_), .A2(G183gat), .A3(G190gat), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT78), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n320_), .B1(new_n334_), .B2(new_n325_), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT88), .B1(new_n335_), .B2(new_n329_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n331_), .A2(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NOR3_X1   g138(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n318_), .B1(new_n337_), .B2(new_n341_), .ZN(new_n342_));
  OR2_X1    g141(.A1(G169gat), .A2(G176gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G169gat), .A2(G176gat), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n343_), .A2(KEYINPUT24), .A3(new_n344_), .ZN(new_n345_));
  OR3_X1    g144(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n322_), .A2(KEYINPUT25), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT25), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(G183gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n347_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(G190gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT26), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT26), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(G190gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n345_), .B(new_n346_), .C1(new_n350_), .C2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G183gat), .A2(G190gat), .ZN(new_n357_));
  AOI22_X1  g156(.A1(new_n323_), .A2(G190gat), .B1(KEYINPUT23), .B2(new_n357_), .ZN(new_n358_));
  OR2_X1    g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n286_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n341_), .ZN(new_n361_));
  AOI211_X1 g160(.A(KEYINPUT89), .B(new_n361_), .C1(new_n331_), .C2(new_n336_), .ZN(new_n362_));
  NOR3_X1   g161(.A1(new_n342_), .A2(new_n360_), .A3(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n341_), .B1(new_n358_), .B2(new_n329_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n364_), .B1(new_n356_), .B2(new_n335_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT79), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  OAI211_X1 g166(.A(new_n364_), .B(KEYINPUT79), .C1(new_n356_), .C2(new_n335_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n286_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G226gat), .A2(G233gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT19), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n371_), .A2(KEYINPUT20), .A3(new_n374_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n317_), .B1(new_n363_), .B2(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n328_), .B1(new_n327_), .B2(new_n330_), .ZN(new_n377_));
  NOR3_X1   g176(.A1(new_n335_), .A2(KEYINPUT88), .A3(new_n329_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n341_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT89), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n337_), .A2(new_n318_), .A3(new_n341_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n380_), .A2(new_n286_), .A3(new_n381_), .A4(new_n359_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT20), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n383_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n384_));
  NAND4_X1  g183(.A1(new_n382_), .A2(KEYINPUT90), .A3(new_n374_), .A4(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n376_), .A2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n380_), .A2(new_n381_), .A3(new_n359_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(new_n370_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n286_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT20), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n374_), .B1(new_n388_), .B2(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n316_), .B1(new_n386_), .B2(new_n392_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n342_), .A2(new_n362_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n286_), .B1(new_n394_), .B2(new_n359_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n373_), .B1(new_n395_), .B2(new_n390_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n396_), .A2(new_n315_), .A3(new_n376_), .A4(new_n385_), .ZN(new_n397_));
  AOI21_X1  g196(.A(KEYINPUT27), .B1(new_n393_), .B2(new_n397_), .ZN(new_n398_));
  AOI211_X1 g197(.A(new_n373_), .B(new_n390_), .C1(new_n370_), .C2(new_n387_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n379_), .A2(new_n286_), .A3(new_n359_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n374_), .B1(new_n384_), .B2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n316_), .B1(new_n399_), .B2(new_n401_), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n397_), .A2(KEYINPUT27), .A3(new_n402_), .ZN(new_n403_));
  NOR3_X1   g202(.A1(new_n311_), .A2(new_n398_), .A3(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT33), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n266_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(KEYINPUT95), .ZN(new_n407_));
  OR2_X1    g206(.A1(new_n266_), .A2(new_n405_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT95), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n266_), .A2(new_n409_), .A3(new_n405_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n252_), .A2(new_n255_), .A3(new_n247_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n243_), .A2(new_n244_), .A3(new_n249_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n411_), .A2(new_n263_), .A3(new_n412_), .ZN(new_n413_));
  AND3_X1   g212(.A1(new_n393_), .A2(new_n397_), .A3(new_n413_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n407_), .A2(new_n408_), .A3(new_n410_), .A4(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(KEYINPUT96), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n266_), .A2(new_n405_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n393_), .A2(new_n397_), .A3(new_n413_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT96), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n419_), .A2(new_n420_), .A3(new_n410_), .A4(new_n407_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n386_), .A2(new_n392_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n315_), .A2(KEYINPUT32), .ZN(new_n423_));
  XOR2_X1   g222(.A(new_n423_), .B(KEYINPUT97), .Z(new_n424_));
  OR2_X1    g223(.A1(new_n399_), .A2(new_n401_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n423_), .ZN(new_n426_));
  AOI22_X1  g225(.A1(new_n422_), .A2(new_n424_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n267_), .A2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n416_), .A2(new_n421_), .A3(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n310_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n404_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n369_), .B(KEYINPUT30), .ZN(new_n432_));
  INV_X1    g231(.A(G99gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n432_), .B(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(KEYINPUT31), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G15gat), .B(G43gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(KEYINPUT80), .B(KEYINPUT81), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n436_), .B(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G227gat), .A2(G233gat), .ZN(new_n439_));
  INV_X1    g238(.A(G71gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n439_), .B(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n438_), .B(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(new_n242_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n435_), .B(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n202_), .B1(new_n431_), .B2(new_n445_), .ZN(new_n446_));
  AOI22_X1  g245(.A1(new_n415_), .A2(KEYINPUT96), .B1(new_n267_), .B2(new_n427_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n310_), .B1(new_n447_), .B2(new_n421_), .ZN(new_n448_));
  OAI211_X1 g247(.A(KEYINPUT98), .B(new_n444_), .C1(new_n448_), .C2(new_n404_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n446_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n393_), .A2(new_n397_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT27), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n397_), .A2(new_n402_), .A3(KEYINPUT27), .ZN(new_n454_));
  AOI21_X1  g253(.A(KEYINPUT99), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT99), .ZN(new_n456_));
  NOR3_X1   g255(.A1(new_n398_), .A2(new_n403_), .A3(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n430_), .B1(new_n455_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT100), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n430_), .B(KEYINPUT100), .C1(new_n455_), .C2(new_n457_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n460_), .A2(new_n268_), .A3(new_n445_), .A4(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT101), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n444_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n465_), .A2(KEYINPUT101), .A3(new_n268_), .A4(new_n461_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n450_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT12), .ZN(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT65), .B(KEYINPUT6), .ZN(new_n470_));
  INV_X1    g269(.A(G106gat), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n433_), .A2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n470_), .B(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT66), .ZN(new_n474_));
  NOR2_X1   g273(.A1(G99gat), .A2(G106gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT7), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(G85gat), .A2(G92gat), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G85gat), .A2(G92gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  OR2_X1    g281(.A1(KEYINPUT67), .A2(KEYINPUT8), .ZN(new_n483_));
  NAND2_X1  g282(.A1(KEYINPUT67), .A2(KEYINPUT8), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n477_), .A2(new_n482_), .A3(new_n483_), .A4(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT8), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n481_), .B1(new_n473_), .B2(new_n476_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n486_), .B1(new_n487_), .B2(KEYINPUT68), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n488_), .B1(KEYINPUT68), .B2(new_n487_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n485_), .A2(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(KEYINPUT10), .B(G99gat), .Z(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(new_n471_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT64), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT9), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n493_), .B1(new_n480_), .B2(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n480_), .A2(new_n493_), .A3(new_n494_), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n496_), .B(new_n479_), .C1(new_n494_), .C2(new_n480_), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n474_), .B(new_n492_), .C1(new_n495_), .C2(new_n497_), .ZN(new_n498_));
  AND2_X1   g297(.A1(new_n490_), .A2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G57gat), .B(G64gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT11), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT69), .ZN(new_n502_));
  XOR2_X1   g301(.A(G71gat), .B(G78gat), .Z(new_n503_));
  OAI21_X1  g302(.A(new_n503_), .B1(KEYINPUT11), .B2(new_n500_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n502_), .B(new_n504_), .ZN(new_n505_));
  OAI211_X1 g304(.A(KEYINPUT70), .B(new_n469_), .C1(new_n499_), .C2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n499_), .A2(new_n505_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n505_), .B1(new_n490_), .B2(new_n498_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT70), .ZN(new_n509_));
  OAI21_X1  g308(.A(KEYINPUT12), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n506_), .A2(new_n507_), .A3(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G230gat), .A2(G233gat), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n507_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n513_), .B1(new_n516_), .B2(new_n508_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  XOR2_X1   g317(.A(G120gat), .B(G148gat), .Z(new_n519_));
  XNOR2_X1  g318(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G176gat), .B(G204gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n518_), .A2(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n515_), .A2(new_n517_), .A3(new_n523_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  OR2_X1    g326(.A1(new_n527_), .A2(KEYINPUT13), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(KEYINPUT13), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  XOR2_X1   g330(.A(KEYINPUT75), .B(G8gat), .Z(new_n532_));
  INV_X1    g331(.A(G1gat), .ZN(new_n533_));
  OAI21_X1  g332(.A(KEYINPUT14), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G15gat), .B(G22gat), .ZN(new_n535_));
  AND2_X1   g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G1gat), .B(G8gat), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n537_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  XOR2_X1   g339(.A(G29gat), .B(G36gat), .Z(new_n541_));
  XOR2_X1   g340(.A(G43gat), .B(G50gat), .Z(new_n542_));
  XOR2_X1   g341(.A(new_n541_), .B(new_n542_), .Z(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n540_), .B(new_n544_), .ZN(new_n545_));
  XOR2_X1   g344(.A(new_n543_), .B(KEYINPUT15), .Z(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n547_), .A2(new_n540_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n548_), .B1(new_n544_), .B2(new_n540_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G229gat), .A2(G233gat), .ZN(new_n550_));
  MUX2_X1   g349(.A(new_n545_), .B(new_n549_), .S(new_n550_), .Z(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(KEYINPUT77), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G113gat), .B(G141gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G169gat), .B(G197gat), .ZN(new_n554_));
  XOR2_X1   g353(.A(new_n553_), .B(new_n554_), .Z(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n552_), .B(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n531_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n468_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G231gat), .A2(G233gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n540_), .B(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(new_n505_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT17), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G127gat), .B(G155gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT16), .ZN(new_n565_));
  XOR2_X1   g364(.A(G183gat), .B(G211gat), .Z(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n562_), .B1(new_n563_), .B2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(KEYINPUT17), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n568_), .B1(new_n569_), .B2(new_n562_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT76), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  OR2_X1    g371(.A1(new_n499_), .A2(new_n547_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(G232gat), .A2(G233gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT34), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n575_), .A2(KEYINPUT35), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n576_), .B1(new_n499_), .B2(new_n544_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n573_), .A2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n578_), .A2(KEYINPUT35), .A3(new_n575_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G190gat), .B(G218gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT72), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G134gat), .B(G162gat), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n581_), .B(new_n582_), .Z(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n584_), .A2(KEYINPUT36), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n575_), .A2(KEYINPUT35), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n573_), .A2(new_n577_), .A3(new_n586_), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n579_), .A2(new_n585_), .A3(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n583_), .B(KEYINPUT36), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n590_), .B1(new_n579_), .B2(new_n587_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n588_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT37), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT74), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n592_), .A2(KEYINPUT74), .A3(new_n593_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n588_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n579_), .A2(new_n587_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n589_), .B(KEYINPUT73), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n598_), .A2(new_n601_), .ZN(new_n602_));
  AOI22_X1  g401(.A1(new_n596_), .A2(new_n597_), .B1(KEYINPUT37), .B2(new_n602_), .ZN(new_n603_));
  NOR3_X1   g402(.A1(new_n559_), .A2(new_n572_), .A3(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n604_), .A2(new_n533_), .A3(new_n267_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT38), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n592_), .B(KEYINPUT102), .ZN(new_n607_));
  NOR3_X1   g406(.A1(new_n559_), .A2(new_n572_), .A3(new_n607_), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n608_), .A2(new_n267_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n606_), .B1(new_n533_), .B2(new_n609_), .ZN(G1324gat));
  NOR2_X1   g409(.A1(new_n455_), .A2(new_n457_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n604_), .A2(new_n532_), .A3(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n608_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n611_), .ZN(new_n614_));
  OAI21_X1  g413(.A(G8gat), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n615_), .A2(KEYINPUT39), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n615_), .A2(KEYINPUT39), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n612_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT40), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  OAI211_X1 g419(.A(KEYINPUT40), .B(new_n612_), .C1(new_n616_), .C2(new_n617_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(G1325gat));
  INV_X1    g421(.A(G15gat), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n604_), .A2(new_n623_), .A3(new_n445_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n608_), .A2(new_n445_), .ZN(new_n625_));
  AND3_X1   g424(.A1(new_n625_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n626_));
  AOI21_X1  g425(.A(KEYINPUT41), .B1(new_n625_), .B2(G15gat), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n624_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n628_), .B(KEYINPUT103), .Z(G1326gat));
  INV_X1    g428(.A(G22gat), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n630_), .B1(new_n608_), .B2(new_n310_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT42), .Z(new_n632_));
  NAND3_X1  g431(.A1(new_n604_), .A2(new_n630_), .A3(new_n310_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(G1327gat));
  NAND2_X1  g433(.A1(new_n607_), .A2(new_n572_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n559_), .A2(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(G29gat), .B1(new_n636_), .B2(new_n267_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(KEYINPUT104), .A2(KEYINPUT44), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT43), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n468_), .A2(new_n639_), .A3(new_n603_), .ZN(new_n640_));
  AOI22_X1  g439(.A1(new_n446_), .A2(new_n449_), .B1(new_n464_), .B2(new_n466_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n602_), .A2(KEYINPUT37), .ZN(new_n642_));
  AOI21_X1  g441(.A(KEYINPUT74), .B1(new_n592_), .B2(new_n593_), .ZN(new_n643_));
  NOR4_X1   g442(.A1(new_n588_), .A2(new_n591_), .A3(new_n595_), .A4(KEYINPUT37), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n642_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(KEYINPUT43), .B1(new_n641_), .B2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n640_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n558_), .A2(new_n572_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n638_), .B1(new_n647_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n647_), .A2(new_n649_), .A3(new_n638_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n267_), .A2(G29gat), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n637_), .B1(new_n653_), .B2(new_n654_), .ZN(G1328gat));
  INV_X1    g454(.A(KEYINPUT46), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(KEYINPUT107), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n614_), .A2(G36gat), .ZN(new_n658_));
  XNOR2_X1  g457(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n659_));
  AND3_X1   g458(.A1(new_n636_), .A2(new_n658_), .A3(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n659_), .B1(new_n636_), .B2(new_n658_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n657_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n652_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n611_), .B1(new_n663_), .B2(new_n650_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n662_), .B1(new_n664_), .B2(G36gat), .ZN(new_n665_));
  AOI21_X1  g464(.A(KEYINPUT107), .B1(new_n656_), .B2(KEYINPUT106), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n665_), .B(new_n666_), .ZN(G1329gat));
  NAND2_X1  g466(.A1(new_n445_), .A2(G43gat), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n668_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n669_));
  AOI21_X1  g468(.A(G43gat), .B1(new_n636_), .B2(new_n445_), .ZN(new_n670_));
  OR3_X1    g469(.A1(new_n669_), .A2(KEYINPUT47), .A3(new_n670_), .ZN(new_n671_));
  OAI21_X1  g470(.A(KEYINPUT47), .B1(new_n669_), .B2(new_n670_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1330gat));
  AOI21_X1  g472(.A(G50gat), .B1(new_n636_), .B2(new_n310_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n310_), .A2(G50gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n674_), .B1(new_n653_), .B2(new_n675_), .ZN(G1331gat));
  INV_X1    g475(.A(new_n557_), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n641_), .A2(new_n530_), .A3(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n607_), .ZN(new_n679_));
  AND3_X1   g478(.A1(new_n678_), .A2(new_n571_), .A3(new_n679_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n680_), .A2(G57gat), .A3(new_n267_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT108), .ZN(new_n682_));
  INV_X1    g481(.A(G57gat), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n603_), .A2(new_n572_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n678_), .A2(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n683_), .B1(new_n685_), .B2(new_n268_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n682_), .A2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(KEYINPUT109), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT109), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n682_), .A2(new_n689_), .A3(new_n686_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(G1332gat));
  INV_X1    g490(.A(G64gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n692_), .B1(new_n680_), .B2(new_n611_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT48), .Z(new_n694_));
  INV_X1    g493(.A(new_n685_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n695_), .A2(new_n692_), .A3(new_n611_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n696_), .ZN(G1333gat));
  AOI21_X1  g496(.A(new_n440_), .B1(new_n680_), .B2(new_n445_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT49), .Z(new_n699_));
  NAND3_X1  g498(.A1(new_n695_), .A2(new_n440_), .A3(new_n445_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1334gat));
  INV_X1    g500(.A(G78gat), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n702_), .B1(new_n680_), .B2(new_n310_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n703_), .B(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n695_), .A2(new_n702_), .A3(new_n310_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(G1335gat));
  NOR3_X1   g506(.A1(new_n530_), .A2(new_n677_), .A3(new_n571_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n647_), .A2(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(G85gat), .B1(new_n709_), .B2(new_n268_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n635_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n678_), .A2(new_n711_), .ZN(new_n712_));
  OR3_X1    g511(.A1(new_n712_), .A2(G85gat), .A3(new_n268_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n710_), .A2(new_n713_), .ZN(G1336gat));
  OAI21_X1  g513(.A(G92gat), .B1(new_n709_), .B2(new_n614_), .ZN(new_n715_));
  OR3_X1    g514(.A1(new_n712_), .A2(G92gat), .A3(new_n614_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1337gat));
  OAI21_X1  g516(.A(G99gat), .B1(new_n709_), .B2(new_n444_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n445_), .A2(new_n491_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n718_), .B1(new_n712_), .B2(new_n719_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g520(.A1(new_n678_), .A2(new_n471_), .A3(new_n310_), .A4(new_n711_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT52), .ZN(new_n723_));
  INV_X1    g522(.A(new_n708_), .ZN(new_n724_));
  AOI211_X1 g523(.A(new_n430_), .B(new_n724_), .C1(new_n640_), .C2(new_n646_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n471_), .B1(new_n725_), .B2(KEYINPUT111), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n724_), .B1(new_n640_), .B2(new_n646_), .ZN(new_n727_));
  AOI21_X1  g526(.A(KEYINPUT111), .B1(new_n727_), .B2(new_n310_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n723_), .B1(new_n726_), .B2(new_n729_), .ZN(new_n730_));
  NAND4_X1  g529(.A1(new_n647_), .A2(KEYINPUT111), .A3(new_n310_), .A4(new_n708_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(G106gat), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n732_), .A2(new_n728_), .A3(KEYINPUT52), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n722_), .B1(new_n730_), .B2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(KEYINPUT53), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT53), .ZN(new_n736_));
  OAI211_X1 g535(.A(new_n736_), .B(new_n722_), .C1(new_n730_), .C2(new_n733_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(G1339gat));
  NAND2_X1  g537(.A1(new_n571_), .A2(new_n557_), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT112), .Z(new_n740_));
  NAND3_X1  g539(.A1(new_n740_), .A2(new_n530_), .A3(new_n645_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT54), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n741_), .B(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT57), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT55), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n511_), .B2(new_n513_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n746_), .A2(new_n514_), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n511_), .A2(new_n745_), .A3(new_n513_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n524_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT56), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n749_), .A2(KEYINPUT113), .A3(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(KEYINPUT113), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n752_), .A2(KEYINPUT114), .ZN(new_n753_));
  OAI211_X1 g552(.A(new_n524_), .B(new_n753_), .C1(new_n747_), .C2(new_n748_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n749_), .A2(new_n750_), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n751_), .B(new_n754_), .C1(new_n755_), .C2(KEYINPUT114), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n677_), .A2(new_n526_), .ZN(new_n757_));
  MUX2_X1   g556(.A(new_n549_), .B(new_n545_), .S(new_n550_), .Z(new_n758_));
  MUX2_X1   g557(.A(new_n551_), .B(new_n758_), .S(new_n556_), .Z(new_n759_));
  AOI22_X1  g558(.A1(new_n756_), .A2(new_n757_), .B1(new_n527_), .B2(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n744_), .B1(new_n760_), .B2(new_n607_), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n506_), .A2(new_n507_), .A3(new_n510_), .ZN(new_n762_));
  OAI21_X1  g561(.A(KEYINPUT55), .B1(new_n762_), .B2(new_n512_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(new_n515_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n748_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n523_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n754_), .B1(new_n766_), .B2(new_n752_), .ZN(new_n767_));
  AOI21_X1  g566(.A(KEYINPUT114), .B1(new_n766_), .B2(KEYINPUT56), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n757_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n527_), .A2(new_n759_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n771_), .A2(KEYINPUT57), .A3(new_n679_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT115), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n526_), .A2(new_n759_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n766_), .A2(KEYINPUT56), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n749_), .A2(new_n750_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n774_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n603_), .B(new_n773_), .C1(new_n777_), .C2(KEYINPUT58), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(KEYINPUT58), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n774_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n766_), .A2(KEYINPUT56), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n781_), .B1(new_n782_), .B2(new_n755_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT58), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n645_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n785_), .A2(new_n773_), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n761_), .B(new_n772_), .C1(new_n780_), .C2(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n743_), .B1(new_n787_), .B2(new_n572_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n465_), .A2(new_n461_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(new_n267_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n788_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(G113gat), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(new_n792_), .A3(new_n677_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT59), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n794_), .B1(new_n788_), .B2(new_n790_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n790_), .ZN(new_n796_));
  AOI21_X1  g595(.A(KEYINPUT57), .B1(new_n771_), .B2(new_n679_), .ZN(new_n797_));
  AOI211_X1 g596(.A(new_n744_), .B(new_n607_), .C1(new_n769_), .C2(new_n770_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n777_), .A2(KEYINPUT58), .ZN(new_n800_));
  OAI21_X1  g599(.A(KEYINPUT115), .B1(new_n800_), .B2(new_n645_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n801_), .A2(new_n778_), .A3(new_n779_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n571_), .B1(new_n799_), .B2(new_n802_), .ZN(new_n803_));
  OAI211_X1 g602(.A(KEYINPUT59), .B(new_n796_), .C1(new_n803_), .C2(new_n743_), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n795_), .A2(KEYINPUT116), .A3(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(KEYINPUT116), .B1(new_n795_), .B2(new_n804_), .ZN(new_n806_));
  NOR3_X1   g605(.A1(new_n805_), .A2(new_n806_), .A3(new_n557_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n793_), .B1(new_n807_), .B2(new_n792_), .ZN(G1340gat));
  INV_X1    g607(.A(G120gat), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n809_), .B1(new_n530_), .B2(KEYINPUT60), .ZN(new_n810_));
  OAI21_X1  g609(.A(KEYINPUT117), .B1(new_n809_), .B2(KEYINPUT60), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT117), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n791_), .B(new_n812_), .C1(new_n813_), .C2(new_n810_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n530_), .B1(new_n795_), .B2(new_n804_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n814_), .B1(new_n815_), .B2(new_n809_), .ZN(G1341gat));
  AOI21_X1  g615(.A(G127gat), .B1(new_n791_), .B2(new_n571_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n805_), .A2(new_n806_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT118), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n819_), .A2(G127gat), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n571_), .A2(KEYINPUT118), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n820_), .B1(new_n821_), .B2(G127gat), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n817_), .B1(new_n818_), .B2(new_n822_), .ZN(G1342gat));
  INV_X1    g622(.A(G134gat), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n791_), .A2(new_n824_), .A3(new_n607_), .ZN(new_n825_));
  NOR3_X1   g624(.A1(new_n805_), .A2(new_n806_), .A3(new_n645_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n825_), .B1(new_n826_), .B2(new_n824_), .ZN(G1343gat));
  NAND3_X1  g626(.A1(new_n614_), .A2(new_n267_), .A3(new_n310_), .ZN(new_n828_));
  NOR3_X1   g627(.A1(new_n788_), .A2(new_n445_), .A3(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n677_), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n830_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g630(.A1(new_n829_), .A2(new_n531_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(KEYINPUT119), .B(G148gat), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n832_), .B(new_n833_), .ZN(G1345gat));
  XNOR2_X1  g633(.A(KEYINPUT120), .B(KEYINPUT121), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  XOR2_X1   g635(.A(KEYINPUT61), .B(G155gat), .Z(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n829_), .A2(new_n571_), .A3(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n838_), .B1(new_n829_), .B2(new_n571_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n836_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n841_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n843_), .A2(new_n835_), .A3(new_n839_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n842_), .A2(new_n844_), .ZN(G1346gat));
  AND3_X1   g644(.A1(new_n829_), .A2(G162gat), .A3(new_n603_), .ZN(new_n846_));
  AOI21_X1  g645(.A(G162gat), .B1(new_n829_), .B2(new_n607_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT122), .ZN(new_n848_));
  OR2_X1    g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n847_), .A2(new_n848_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n846_), .B1(new_n849_), .B2(new_n850_), .ZN(G1347gat));
  NOR2_X1   g650(.A1(new_n788_), .A2(new_n310_), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n614_), .A2(new_n267_), .A3(new_n444_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(KEYINPUT22), .B(G169gat), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n852_), .A2(new_n677_), .A3(new_n853_), .A4(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n853_), .A2(new_n677_), .ZN(new_n856_));
  XOR2_X1   g655(.A(new_n856_), .B(KEYINPUT123), .Z(new_n857_));
  NAND2_X1  g656(.A1(new_n852_), .A2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(G169gat), .ZN(new_n859_));
  AND2_X1   g658(.A1(new_n859_), .A2(KEYINPUT62), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n859_), .A2(KEYINPUT62), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n855_), .B1(new_n860_), .B2(new_n861_), .ZN(G1348gat));
  NAND3_X1  g661(.A1(new_n852_), .A2(new_n531_), .A3(new_n853_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g663(.A1(new_n852_), .A2(new_n853_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n865_), .A2(new_n572_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n866_), .A2(G183gat), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n867_), .B1(new_n350_), .B2(new_n866_), .ZN(G1350gat));
  OAI21_X1  g667(.A(G190gat), .B1(new_n865_), .B2(new_n645_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n607_), .A2(new_n352_), .A3(new_n354_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n869_), .B1(new_n865_), .B2(new_n870_), .ZN(G1351gat));
  NOR2_X1   g670(.A1(new_n788_), .A2(new_n445_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n614_), .A2(new_n311_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(new_n677_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(G197gat), .ZN(G1352gat));
  AND3_X1   g676(.A1(new_n872_), .A2(new_n531_), .A3(new_n873_), .ZN(new_n878_));
  INV_X1    g677(.A(G204gat), .ZN(new_n879_));
  OAI21_X1  g678(.A(KEYINPUT124), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT124), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n881_), .B(G204gat), .C1(new_n874_), .C2(new_n530_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n882_), .ZN(new_n883_));
  NAND4_X1  g682(.A1(new_n872_), .A2(new_n879_), .A3(new_n531_), .A4(new_n873_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(KEYINPUT125), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n885_), .ZN(G1353gat));
  INV_X1    g685(.A(KEYINPUT63), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n887_), .A2(new_n272_), .A3(KEYINPUT126), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n888_), .B1(new_n887_), .B2(new_n272_), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n874_), .A2(new_n572_), .A3(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT126), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n891_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n890_), .B(new_n892_), .ZN(G1354gat));
  AOI21_X1  g692(.A(G218gat), .B1(new_n875_), .B2(new_n607_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n603_), .A2(G218gat), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(KEYINPUT127), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n894_), .B1(new_n875_), .B2(new_n896_), .ZN(G1355gat));
endmodule


