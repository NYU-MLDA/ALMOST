//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 1 1 1 0 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1 1 1 1 1 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n722_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n771_, new_n772_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_, new_n890_, new_n891_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n930_, new_n932_, new_n934_, new_n935_, new_n937_,
    new_n939_, new_n941_, new_n942_, new_n943_, new_n944_, new_n946_,
    new_n947_, new_n948_, new_n949_;
  INV_X1    g000(.A(KEYINPUT38), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT69), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT12), .ZN(new_n204_));
  AND3_X1   g003(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n205_));
  AOI21_X1  g004(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  AND2_X1   g007(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n209_));
  NOR2_X1   g008(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n208_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  OAI22_X1  g010(.A1(KEYINPUT66), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n207_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  AND2_X1   g012(.A1(G85gat), .A2(G92gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G85gat), .A2(G92gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n213_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT8), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT8), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n216_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT65), .ZN(new_n222_));
  NOR3_X1   g021(.A1(new_n205_), .A2(new_n206_), .A3(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G99gat), .A2(G106gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT6), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n227_));
  AOI21_X1  g026(.A(KEYINPUT65), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n223_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n211_), .A2(new_n212_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n221_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(G85gat), .ZN(new_n232_));
  INV_X1    g031(.A(G92gat), .ZN(new_n233_));
  NOR3_X1   g032(.A1(new_n232_), .A2(new_n233_), .A3(KEYINPUT9), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n222_), .B1(new_n205_), .B2(new_n206_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n226_), .A2(KEYINPUT65), .A3(new_n227_), .ZN(new_n236_));
  AOI221_X4 g035(.A(new_n234_), .B1(new_n216_), .B2(KEYINPUT9), .C1(new_n235_), .C2(new_n236_), .ZN(new_n237_));
  XOR2_X1   g036(.A(KEYINPUT10), .B(G99gat), .Z(new_n238_));
  INV_X1    g037(.A(KEYINPUT64), .ZN(new_n239_));
  INV_X1    g038(.A(G106gat), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n238_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT10), .B(G99gat), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT64), .B1(new_n242_), .B2(G106gat), .ZN(new_n243_));
  AND2_X1   g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  AOI22_X1  g043(.A1(new_n218_), .A2(new_n231_), .B1(new_n237_), .B2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G57gat), .A2(G64gat), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(G57gat), .A2(G64gat), .ZN(new_n248_));
  OAI21_X1  g047(.A(KEYINPUT11), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G71gat), .B(G78gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n248_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT11), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n253_), .A2(new_n254_), .A3(new_n246_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n250_), .B1(new_n255_), .B2(new_n249_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n252_), .A2(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n204_), .B1(new_n245_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G230gat), .A2(G233gat), .ZN(new_n259_));
  AOI22_X1  g058(.A1(new_n235_), .A2(new_n236_), .B1(KEYINPUT9), .B2(new_n216_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n234_), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n260_), .A2(new_n261_), .A3(new_n243_), .A4(new_n241_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n219_), .B1(new_n213_), .B2(new_n216_), .ZN(new_n263_));
  AND2_X1   g062(.A1(new_n211_), .A2(new_n212_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n235_), .A2(new_n236_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n220_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n262_), .B(new_n257_), .C1(new_n263_), .C2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n216_), .A2(KEYINPUT9), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n265_), .A2(new_n261_), .A3(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n241_), .A2(new_n243_), .ZN(new_n270_));
  OAI22_X1  g069(.A1(new_n266_), .A2(new_n263_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  AND2_X1   g070(.A1(new_n255_), .A2(new_n249_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n251_), .B1(new_n272_), .B2(new_n250_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT67), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT67), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n257_), .A2(new_n275_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n271_), .A2(new_n274_), .A3(new_n276_), .A4(KEYINPUT12), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n258_), .A2(new_n259_), .A3(new_n267_), .A4(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n259_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n245_), .A2(new_n257_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n267_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n279_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(KEYINPUT68), .B(KEYINPUT5), .Z(new_n283_));
  XNOR2_X1  g082(.A(G120gat), .B(G148gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G176gat), .B(G204gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n278_), .A2(new_n282_), .A3(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n288_), .B1(new_n278_), .B2(new_n282_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n203_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n291_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n293_), .A2(KEYINPUT69), .A3(new_n289_), .ZN(new_n294_));
  AND2_X1   g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  OR2_X1    g094(.A1(new_n295_), .A2(KEYINPUT13), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(KEYINPUT13), .ZN(new_n297_));
  AND2_X1   g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT70), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G127gat), .B(G134gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G113gat), .B(G120gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G155gat), .A2(G162gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT94), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT94), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n306_), .A2(G155gat), .A3(G162gat), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT1), .ZN(new_n308_));
  AND3_X1   g107(.A1(new_n305_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n308_), .B1(new_n305_), .B2(new_n307_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(G155gat), .A2(G162gat), .ZN(new_n311_));
  NOR3_X1   g110(.A1(new_n309_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(G141gat), .A2(G148gat), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G141gat), .A2(G148gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n312_), .A2(new_n316_), .ZN(new_n317_));
  AND2_X1   g116(.A1(new_n305_), .A2(new_n307_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n315_), .B(KEYINPUT2), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n313_), .B(KEYINPUT3), .ZN(new_n320_));
  AOI211_X1 g119(.A(new_n311_), .B(new_n318_), .C1(new_n319_), .C2(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n303_), .B1(new_n317_), .B2(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n311_), .B1(new_n320_), .B2(new_n319_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n318_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n325_), .B(new_n302_), .C1(new_n316_), .C2(new_n312_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n322_), .A2(KEYINPUT4), .A3(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G225gat), .A2(G233gat), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n325_), .B1(new_n316_), .B2(new_n312_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT4), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n330_), .A2(new_n331_), .A3(new_n303_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n327_), .A2(new_n329_), .A3(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT99), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n322_), .A2(new_n328_), .A3(new_n326_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT99), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n327_), .A2(new_n336_), .A3(new_n329_), .A4(new_n332_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n334_), .A2(new_n335_), .A3(new_n337_), .ZN(new_n338_));
  XOR2_X1   g137(.A(G1gat), .B(G29gat), .Z(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT101), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G57gat), .B(G85gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT100), .B(KEYINPUT0), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n338_), .A2(new_n345_), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n334_), .A2(new_n344_), .A3(new_n335_), .A4(new_n337_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  XOR2_X1   g147(.A(G64gat), .B(G92gat), .Z(new_n349_));
  XNOR2_X1  g148(.A(G8gat), .B(G36gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  AND2_X1   g152(.A1(new_n353_), .A2(KEYINPUT32), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT20), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G197gat), .B(G204gat), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT21), .ZN(new_n357_));
  OR2_X1    g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G211gat), .B(G218gat), .ZN(new_n359_));
  OR2_X1    g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n356_), .A2(new_n357_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n358_), .A2(new_n361_), .A3(new_n359_), .ZN(new_n362_));
  AND2_X1   g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(KEYINPUT96), .B(KEYINPUT24), .ZN(new_n364_));
  OR2_X1    g163(.A1(G169gat), .A2(G176gat), .ZN(new_n365_));
  OR2_X1    g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G183gat), .A2(G190gat), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT23), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n370_));
  AND2_X1   g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G169gat), .A2(G176gat), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n364_), .A2(new_n372_), .A3(new_n365_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(KEYINPUT25), .B(G183gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT26), .B(G190gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n366_), .A2(new_n371_), .A3(new_n373_), .A4(new_n376_), .ZN(new_n377_));
  XOR2_X1   g176(.A(KEYINPUT88), .B(G176gat), .Z(new_n378_));
  XNOR2_X1  g177(.A(KEYINPUT22), .B(G169gat), .ZN(new_n379_));
  AOI22_X1  g178(.A1(new_n378_), .A2(new_n379_), .B1(G169gat), .B2(G176gat), .ZN(new_n380_));
  OAI211_X1 g179(.A(new_n369_), .B(new_n370_), .C1(G183gat), .C2(G190gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  AND2_X1   g181(.A1(new_n377_), .A2(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n355_), .B1(new_n363_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(KEYINPUT103), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n365_), .A2(KEYINPUT24), .A3(new_n372_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT85), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT26), .ZN(new_n388_));
  OR3_X1    g187(.A1(new_n387_), .A2(new_n388_), .A3(G190gat), .ZN(new_n389_));
  AND2_X1   g188(.A1(KEYINPUT86), .A2(KEYINPUT26), .ZN(new_n390_));
  NOR2_X1   g189(.A1(KEYINPUT86), .A2(KEYINPUT26), .ZN(new_n391_));
  OAI21_X1  g190(.A(G190gat), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n387_), .B1(new_n388_), .B2(G190gat), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n389_), .A2(new_n392_), .A3(new_n374_), .A4(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT87), .ZN(new_n395_));
  OR3_X1    g194(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n395_), .B1(new_n371_), .B2(new_n396_), .ZN(new_n397_));
  AND4_X1   g196(.A1(new_n395_), .A2(new_n396_), .A3(new_n369_), .A4(new_n370_), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n386_), .B(new_n394_), .C1(new_n397_), .C2(new_n398_), .ZN(new_n399_));
  OR2_X1    g198(.A1(new_n381_), .A2(KEYINPUT89), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n381_), .A2(KEYINPUT89), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n400_), .A2(new_n380_), .A3(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n399_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n360_), .A2(new_n362_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n377_), .A2(new_n382_), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT20), .B1(new_n404_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT103), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n385_), .A2(new_n405_), .A3(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G226gat), .A2(G233gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  AND3_X1   g212(.A1(new_n410_), .A2(KEYINPUT104), .A3(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n363_), .A2(new_n402_), .A3(new_n399_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n413_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n404_), .A2(new_n406_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n415_), .A2(KEYINPUT20), .A3(new_n416_), .A4(new_n417_), .ZN(new_n418_));
  AOI22_X1  g217(.A1(new_n410_), .A2(new_n413_), .B1(KEYINPUT104), .B2(new_n418_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n354_), .B1(new_n414_), .B2(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n354_), .B(KEYINPUT102), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n415_), .A2(KEYINPUT20), .A3(new_n417_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(new_n413_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n384_), .A2(new_n405_), .A3(new_n416_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  OR2_X1    g224(.A1(new_n421_), .A2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n348_), .A2(new_n420_), .A3(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT105), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n353_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n425_), .A2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n423_), .A2(new_n353_), .A3(new_n424_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n431_), .A2(KEYINPUT98), .A3(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT98), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n425_), .A2(new_n434_), .A3(new_n430_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n327_), .A2(new_n328_), .A3(new_n332_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n322_), .A2(new_n329_), .A3(new_n326_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n345_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n347_), .A2(KEYINPUT33), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n347_), .A2(KEYINPUT33), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n436_), .B(new_n439_), .C1(new_n440_), .C2(new_n441_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n348_), .A2(new_n420_), .A3(KEYINPUT105), .A4(new_n426_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n429_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(KEYINPUT93), .B(KEYINPUT31), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G71gat), .B(G99gat), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  OR2_X1    g247(.A1(G15gat), .A2(G43gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G15gat), .A2(G43gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT90), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n449_), .A2(KEYINPUT90), .A3(new_n450_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G227gat), .A2(G233gat), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n453_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n455_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n448_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n458_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n460_), .A2(new_n447_), .A3(new_n456_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n459_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT30), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n399_), .A2(new_n402_), .A3(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n463_), .B1(new_n399_), .B2(new_n402_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n462_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT92), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n403_), .A2(KEYINPUT30), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(new_n464_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT92), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n470_), .A2(new_n471_), .A3(new_n462_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n468_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT91), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n474_), .B1(new_n470_), .B2(new_n462_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n462_), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n476_), .A2(new_n469_), .A3(KEYINPUT91), .A4(new_n464_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n475_), .A2(new_n477_), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n473_), .A2(new_n478_), .A3(new_n303_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n303_), .B1(new_n473_), .B2(new_n478_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n446_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n473_), .A2(new_n478_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(new_n302_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n473_), .A2(new_n478_), .A3(new_n303_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n483_), .A2(new_n445_), .A3(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n481_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT28), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n317_), .A2(new_n321_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT29), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n487_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  NOR3_X1   g289(.A1(new_n330_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G228gat), .A2(G233gat), .ZN(new_n492_));
  INV_X1    g291(.A(G22gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  OR3_X1    g293(.A1(new_n490_), .A2(new_n491_), .A3(new_n494_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n494_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n404_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(G50gat), .ZN(new_n499_));
  XOR2_X1   g298(.A(G78gat), .B(G106gat), .Z(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(G50gat), .ZN(new_n502_));
  OAI211_X1 g301(.A(new_n502_), .B(new_n404_), .C1(new_n488_), .C2(new_n489_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n499_), .A2(new_n501_), .A3(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n501_), .B1(new_n499_), .B2(new_n503_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n497_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n506_), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n508_), .A2(new_n495_), .A3(new_n496_), .A4(new_n504_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n507_), .A2(new_n509_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n486_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n444_), .A2(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n353_), .B(KEYINPUT106), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n513_), .B1(new_n414_), .B2(new_n419_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n514_), .A2(KEYINPUT27), .A3(new_n432_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT27), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n433_), .A2(new_n516_), .A3(new_n435_), .ZN(new_n517_));
  AND2_X1   g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n348_), .ZN(new_n519_));
  AND3_X1   g318(.A1(new_n481_), .A2(new_n485_), .A3(new_n510_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n510_), .B1(new_n481_), .B2(new_n485_), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n518_), .B(new_n519_), .C1(new_n520_), .C2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n512_), .A2(new_n522_), .ZN(new_n523_));
  AND2_X1   g322(.A1(new_n299_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT83), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G1gat), .B(G8gat), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G1gat), .A2(G8gat), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT14), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G15gat), .B(G22gat), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n527_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n529_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(new_n526_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n531_), .A2(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(G29gat), .B(G36gat), .Z(new_n535_));
  XNOR2_X1  g334(.A(G43gat), .B(G50gat), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  XOR2_X1   g336(.A(G43gat), .B(G50gat), .Z(new_n538_));
  XNOR2_X1  g337(.A(G29gat), .B(G36gat), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n537_), .A2(new_n540_), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n534_), .A2(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n534_), .A2(new_n541_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n525_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n534_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n541_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n534_), .A2(new_n541_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n547_), .A2(KEYINPUT83), .A3(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G229gat), .A2(G233gat), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n544_), .A2(new_n549_), .A3(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT15), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n541_), .A2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n537_), .A2(new_n540_), .A3(KEYINPUT15), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n550_), .B(new_n547_), .C1(new_n556_), .C2(new_n545_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n552_), .A2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G113gat), .B(G141gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G169gat), .B(G197gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  AND3_X1   g361(.A1(new_n558_), .A2(KEYINPUT84), .A3(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n562_), .B1(new_n558_), .B2(KEYINPUT84), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  XOR2_X1   g364(.A(G190gat), .B(G218gat), .Z(new_n566_));
  XNOR2_X1  g365(.A(G134gat), .B(G162gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT36), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n262_), .B(new_n546_), .C1(new_n263_), .C2(new_n266_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G232gat), .A2(G233gat), .ZN(new_n571_));
  XOR2_X1   g370(.A(new_n571_), .B(KEYINPUT34), .Z(new_n572_));
  INV_X1    g371(.A(KEYINPUT35), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  XOR2_X1   g373(.A(new_n574_), .B(KEYINPUT72), .Z(new_n575_));
  NAND2_X1  g374(.A1(new_n554_), .A2(new_n555_), .ZN(new_n576_));
  AND3_X1   g375(.A1(new_n271_), .A2(KEYINPUT71), .A3(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(KEYINPUT71), .B1(new_n271_), .B2(new_n576_), .ZN(new_n578_));
  OAI211_X1 g377(.A(new_n570_), .B(new_n575_), .C1(new_n577_), .C2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT73), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n580_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n572_), .A2(new_n573_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n579_), .A2(new_n581_), .A3(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n579_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n569_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT37), .ZN(new_n587_));
  INV_X1    g386(.A(new_n570_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT71), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n589_), .B1(new_n245_), .B2(new_n556_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n271_), .A2(KEYINPUT71), .A3(new_n576_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n588_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(KEYINPUT73), .B1(new_n590_), .B2(new_n591_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n582_), .ZN(new_n594_));
  OAI211_X1 g393(.A(new_n592_), .B(new_n575_), .C1(new_n593_), .C2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT36), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n568_), .A2(new_n596_), .ZN(new_n597_));
  XOR2_X1   g396(.A(new_n597_), .B(KEYINPUT74), .Z(new_n598_));
  NAND3_X1  g397(.A1(new_n595_), .A2(new_n583_), .A3(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n586_), .A2(new_n587_), .A3(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(KEYINPUT76), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n586_), .A2(KEYINPUT75), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT75), .ZN(new_n603_));
  OAI211_X1 g402(.A(new_n603_), .B(new_n569_), .C1(new_n584_), .C2(new_n585_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n602_), .A2(new_n599_), .A3(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n601_), .B1(KEYINPUT37), .B2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT76), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n604_), .A2(new_n599_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n569_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n609_), .B1(new_n595_), .B2(new_n583_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n610_), .A2(new_n603_), .ZN(new_n611_));
  OAI211_X1 g410(.A(new_n607_), .B(KEYINPUT37), .C1(new_n608_), .C2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(KEYINPUT77), .B1(new_n606_), .B2(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(KEYINPUT37), .B1(new_n608_), .B2(new_n611_), .ZN(new_n615_));
  AND3_X1   g414(.A1(new_n595_), .A2(new_n583_), .A3(new_n598_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n616_), .A2(new_n610_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n607_), .B1(new_n617_), .B2(new_n587_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n615_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT77), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n619_), .A2(new_n620_), .A3(new_n612_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n614_), .A2(new_n621_), .ZN(new_n622_));
  XOR2_X1   g421(.A(G183gat), .B(G211gat), .Z(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT80), .ZN(new_n624_));
  XOR2_X1   g423(.A(G127gat), .B(G155gat), .Z(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT79), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n624_), .B(new_n626_), .ZN(new_n627_));
  XOR2_X1   g426(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(KEYINPUT17), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n630_), .A2(KEYINPUT81), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(KEYINPUT81), .ZN(new_n632_));
  NAND2_X1  g431(.A1(G231gat), .A2(G233gat), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n534_), .B(new_n633_), .Z(new_n634_));
  NAND2_X1  g433(.A1(new_n274_), .A2(new_n276_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n631_), .A2(new_n632_), .A3(new_n636_), .ZN(new_n637_));
  XOR2_X1   g436(.A(new_n637_), .B(KEYINPUT82), .Z(new_n638_));
  OR2_X1    g437(.A1(new_n629_), .A2(KEYINPUT17), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n634_), .B(new_n273_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n639_), .A2(new_n630_), .A3(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n638_), .A2(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n622_), .A2(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n524_), .A2(new_n565_), .A3(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n644_), .A2(G1gat), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT107), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n645_), .A2(new_n646_), .A3(new_n348_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n646_), .B1(new_n645_), .B2(new_n348_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n202_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n649_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n651_), .A2(KEYINPUT38), .A3(new_n647_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n565_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n298_), .A2(new_n653_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n654_), .A2(new_n523_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n642_), .A2(new_n617_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  OAI21_X1  g456(.A(G1gat), .B1(new_n657_), .B2(new_n519_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT108), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n650_), .A2(new_n652_), .A3(new_n659_), .ZN(G1324gat));
  NOR3_X1   g459(.A1(new_n644_), .A2(G8gat), .A3(new_n518_), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n657_), .A2(new_n518_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(G8gat), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(KEYINPUT39), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT39), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n662_), .A2(new_n665_), .A3(G8gat), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n661_), .B1(new_n664_), .B2(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT40), .ZN(G1325gat));
  INV_X1    g467(.A(new_n486_), .ZN(new_n669_));
  OAI21_X1  g468(.A(G15gat), .B1(new_n657_), .B2(new_n669_), .ZN(new_n670_));
  XOR2_X1   g469(.A(KEYINPUT109), .B(KEYINPUT41), .Z(new_n671_));
  XOR2_X1   g470(.A(new_n670_), .B(new_n671_), .Z(new_n672_));
  NOR3_X1   g471(.A1(new_n644_), .A2(G15gat), .A3(new_n669_), .ZN(new_n673_));
  OR2_X1    g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1326gat));
  INV_X1    g473(.A(new_n510_), .ZN(new_n675_));
  OAI21_X1  g474(.A(G22gat), .B1(new_n657_), .B2(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT42), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n510_), .A2(new_n493_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n677_), .B1(new_n644_), .B2(new_n678_), .ZN(G1327gat));
  AND3_X1   g478(.A1(new_n619_), .A2(new_n620_), .A3(new_n612_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n620_), .B1(new_n619_), .B2(new_n612_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n523_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT43), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  OAI211_X1 g483(.A(new_n523_), .B(KEYINPUT43), .C1(new_n680_), .C2(new_n681_), .ZN(new_n685_));
  AND3_X1   g484(.A1(new_n684_), .A2(new_n642_), .A3(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n686_), .A2(KEYINPUT44), .A3(new_n654_), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n684_), .A2(new_n642_), .A3(new_n654_), .A4(new_n685_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT44), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n687_), .A2(new_n348_), .A3(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(G29gat), .ZN(new_n692_));
  INV_X1    g491(.A(new_n642_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n617_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n655_), .A2(new_n695_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n519_), .A2(G29gat), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT110), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n692_), .A2(new_n699_), .ZN(G1328gat));
  AND2_X1   g499(.A1(new_n688_), .A2(new_n689_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n701_), .A2(new_n518_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(new_n687_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(G36gat), .ZN(new_n704_));
  INV_X1    g503(.A(G36gat), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n518_), .B(KEYINPUT111), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n696_), .A2(new_n705_), .A3(new_n707_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(KEYINPUT112), .B(KEYINPUT45), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n708_), .B(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n704_), .A2(KEYINPUT46), .A3(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT46), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n705_), .B1(new_n702_), .B2(new_n687_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n713_), .B1(new_n714_), .B2(new_n710_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n712_), .A2(new_n715_), .ZN(G1329gat));
  NAND2_X1  g515(.A1(new_n687_), .A2(G43gat), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n690_), .A2(new_n486_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n696_), .A2(new_n486_), .ZN(new_n719_));
  OAI22_X1  g518(.A1(new_n717_), .A2(new_n718_), .B1(G43gat), .B2(new_n719_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g520(.A(G50gat), .B1(new_n696_), .B2(new_n510_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n687_), .A2(G50gat), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n701_), .A2(new_n675_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n722_), .B1(new_n723_), .B2(new_n724_), .ZN(G1331gat));
  NAND2_X1  g524(.A1(new_n643_), .A2(new_n298_), .ZN(new_n726_));
  OR2_X1    g525(.A1(new_n726_), .A2(KEYINPUT113), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n565_), .B1(new_n512_), .B2(new_n522_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(KEYINPUT113), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n727_), .A2(new_n728_), .A3(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(G57gat), .B1(new_n730_), .B2(new_n348_), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n298_), .B(KEYINPUT70), .Z(new_n732_));
  AND2_X1   g531(.A1(new_n732_), .A2(new_n728_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(new_n656_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n734_), .A2(new_n519_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n731_), .B1(G57gat), .B2(new_n735_), .ZN(G1332gat));
  OAI21_X1  g535(.A(G64gat), .B1(new_n734_), .B2(new_n706_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT48), .ZN(new_n738_));
  INV_X1    g537(.A(G64gat), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n730_), .A2(new_n739_), .A3(new_n707_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n740_), .ZN(G1333gat));
  INV_X1    g540(.A(G71gat), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n730_), .A2(new_n742_), .A3(new_n486_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n733_), .A2(new_n656_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n742_), .B1(new_n744_), .B2(new_n486_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(KEYINPUT114), .B(KEYINPUT49), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n745_), .A2(new_n746_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n743_), .B1(new_n747_), .B2(new_n748_), .ZN(G1334gat));
  NAND2_X1  g548(.A1(new_n744_), .A2(new_n510_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(G78gat), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT115), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT115), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n750_), .A2(new_n753_), .A3(G78gat), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n752_), .A2(KEYINPUT50), .A3(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT50), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n753_), .B1(new_n750_), .B2(G78gat), .ZN(new_n757_));
  INV_X1    g556(.A(G78gat), .ZN(new_n758_));
  AOI211_X1 g557(.A(KEYINPUT115), .B(new_n758_), .C1(new_n744_), .C2(new_n510_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n756_), .B1(new_n757_), .B2(new_n759_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n730_), .A2(new_n758_), .A3(new_n510_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n755_), .A2(new_n760_), .A3(new_n761_), .ZN(G1335gat));
  NAND4_X1  g561(.A1(new_n686_), .A2(KEYINPUT116), .A3(new_n653_), .A4(new_n298_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT116), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n684_), .A2(new_n642_), .A3(new_n298_), .A4(new_n685_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n764_), .B1(new_n765_), .B2(new_n565_), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n763_), .A2(G85gat), .A3(new_n766_), .A4(new_n348_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n733_), .A2(new_n695_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n232_), .B1(new_n768_), .B2(new_n519_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n767_), .A2(new_n769_), .ZN(G1336gat));
  NAND4_X1  g569(.A1(new_n763_), .A2(G92gat), .A3(new_n766_), .A4(new_n707_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n233_), .B1(new_n768_), .B2(new_n518_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n771_), .A2(new_n772_), .ZN(G1337gat));
  NAND3_X1  g572(.A1(new_n763_), .A2(new_n486_), .A3(new_n766_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(G99gat), .ZN(new_n775_));
  INV_X1    g574(.A(new_n768_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n776_), .A2(new_n238_), .A3(new_n486_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(KEYINPUT117), .B(KEYINPUT51), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n775_), .A2(new_n777_), .A3(new_n779_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(G1338gat));
  NAND3_X1  g582(.A1(new_n776_), .A2(new_n240_), .A3(new_n510_), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n765_), .A2(new_n565_), .A3(new_n675_), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n785_), .A2(KEYINPUT52), .A3(new_n240_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n686_), .A2(new_n653_), .A3(new_n298_), .A4(new_n510_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n787_), .B1(new_n788_), .B2(G106gat), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n784_), .B1(new_n786_), .B2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT53), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n792_), .B(new_n784_), .C1(new_n786_), .C2(new_n789_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n791_), .A2(new_n793_), .ZN(G1339gat));
  INV_X1    g593(.A(G113gat), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n518_), .A2(new_n348_), .A3(new_n521_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n565_), .A2(KEYINPUT118), .A3(new_n289_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n558_), .A2(KEYINPUT84), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(new_n561_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n558_), .A2(KEYINPUT84), .A3(new_n562_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n799_), .A2(new_n800_), .A3(new_n289_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT118), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n797_), .A2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n258_), .A2(new_n267_), .A3(new_n277_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT119), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT119), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n258_), .A2(new_n807_), .A3(new_n267_), .A4(new_n277_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n806_), .A2(new_n279_), .A3(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n805_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n810_), .A2(KEYINPUT120), .A3(KEYINPUT55), .A4(new_n259_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n278_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT120), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n814_), .B1(new_n278_), .B2(new_n812_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n809_), .A2(new_n811_), .A3(new_n813_), .A4(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n287_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT56), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n816_), .A2(KEYINPUT56), .A3(new_n287_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n804_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n558_), .A2(new_n561_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n544_), .A2(new_n549_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n550_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n547_), .B1(new_n556_), .B2(new_n545_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n551_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n562_), .B1(new_n824_), .B2(new_n826_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n822_), .A2(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n292_), .A2(new_n294_), .A3(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT121), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT121), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n292_), .A2(new_n294_), .A3(new_n831_), .A4(new_n828_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n694_), .B1(new_n821_), .B2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(KEYINPUT57), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT57), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n836_), .B(new_n694_), .C1(new_n821_), .C2(new_n833_), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n835_), .A2(new_n837_), .ZN(new_n838_));
  AND3_X1   g637(.A1(new_n816_), .A2(KEYINPUT56), .A3(new_n287_), .ZN(new_n839_));
  AOI21_X1  g638(.A(KEYINPUT56), .B1(new_n816_), .B2(new_n287_), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n289_), .B(new_n828_), .C1(new_n839_), .C2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT58), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n819_), .A2(new_n820_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n844_), .A2(KEYINPUT58), .A3(new_n289_), .A4(new_n828_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n846_), .B1(new_n614_), .B2(new_n621_), .ZN(new_n847_));
  OAI21_X1  g646(.A(KEYINPUT122), .B1(new_n838_), .B2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n835_), .A2(new_n837_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT122), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n680_), .A2(new_n681_), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n849_), .B(new_n850_), .C1(new_n851_), .C2(new_n846_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n848_), .A2(new_n642_), .A3(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT54), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n565_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n851_), .A2(new_n854_), .A3(new_n693_), .A4(new_n855_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n614_), .A2(new_n693_), .A3(new_n621_), .A4(new_n855_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(KEYINPUT54), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n856_), .A2(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n796_), .B1(new_n853_), .B2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT123), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  AOI211_X1 g661(.A(KEYINPUT123), .B(new_n796_), .C1(new_n853_), .C2(new_n859_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n565_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n642_), .B1(new_n838_), .B2(new_n847_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n859_), .A2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n867_));
  INV_X1    g666(.A(new_n796_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n866_), .A2(new_n867_), .A3(new_n868_), .ZN(new_n869_));
  OAI211_X1 g668(.A(G113gat), .B(new_n869_), .C1(new_n860_), .C2(new_n867_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  AOI22_X1  g670(.A1(new_n795_), .A2(new_n864_), .B1(new_n871_), .B2(new_n565_), .ZN(G1340gat));
  INV_X1    g671(.A(G120gat), .ZN(new_n873_));
  INV_X1    g672(.A(new_n298_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n873_), .B1(new_n874_), .B2(KEYINPUT60), .ZN(new_n875_));
  OAI221_X1 g674(.A(new_n875_), .B1(KEYINPUT60), .B2(new_n873_), .C1(new_n862_), .C2(new_n863_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n869_), .B1(new_n860_), .B2(new_n867_), .ZN(new_n877_));
  OAI21_X1  g676(.A(G120gat), .B1(new_n877_), .B2(new_n299_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n878_), .ZN(G1341gat));
  INV_X1    g678(.A(G127gat), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n693_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(KEYINPUT124), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n869_), .B(new_n882_), .C1(new_n860_), .C2(new_n867_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT124), .ZN(new_n885_));
  OAI21_X1  g684(.A(G127gat), .B1(new_n642_), .B2(new_n885_), .ZN(new_n886_));
  AOI22_X1  g685(.A1(new_n880_), .A2(new_n881_), .B1(new_n884_), .B2(new_n886_), .ZN(G1342gat));
  OAI211_X1 g686(.A(new_n622_), .B(new_n869_), .C1(new_n860_), .C2(new_n867_), .ZN(new_n888_));
  INV_X1    g687(.A(G134gat), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n617_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n890_), .B1(new_n889_), .B2(new_n891_), .ZN(G1343gat));
  XNOR2_X1  g691(.A(KEYINPUT125), .B(G141gat), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n853_), .A2(new_n859_), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n894_), .A2(new_n348_), .A3(new_n520_), .A4(new_n706_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n893_), .B1(new_n896_), .B2(new_n565_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n893_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n895_), .A2(new_n653_), .A3(new_n898_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n897_), .A2(new_n899_), .ZN(G1344gat));
  OR3_X1    g699(.A1(new_n895_), .A2(G148gat), .A3(new_n299_), .ZN(new_n901_));
  OAI21_X1  g700(.A(G148gat), .B1(new_n895_), .B2(new_n299_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1345gat));
  XNOR2_X1  g702(.A(KEYINPUT61), .B(G155gat), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n904_), .B1(new_n896_), .B2(new_n693_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n904_), .ZN(new_n906_));
  NOR3_X1   g705(.A1(new_n895_), .A2(new_n642_), .A3(new_n906_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n905_), .A2(new_n907_), .ZN(G1346gat));
  NAND2_X1  g707(.A1(new_n896_), .A2(new_n617_), .ZN(new_n909_));
  INV_X1    g708(.A(G162gat), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n851_), .A2(new_n910_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(KEYINPUT126), .ZN(new_n912_));
  AOI22_X1  g711(.A1(new_n909_), .A2(new_n910_), .B1(new_n896_), .B2(new_n912_), .ZN(G1347gat));
  NOR2_X1   g712(.A1(new_n706_), .A2(new_n348_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(new_n521_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  NAND4_X1  g715(.A1(new_n866_), .A2(new_n565_), .A3(new_n379_), .A4(new_n916_), .ZN(new_n917_));
  AOI211_X1 g716(.A(new_n653_), .B(new_n915_), .C1(new_n859_), .C2(new_n865_), .ZN(new_n918_));
  INV_X1    g717(.A(G169gat), .ZN(new_n919_));
  OAI211_X1 g718(.A(new_n917_), .B(KEYINPUT62), .C1(new_n918_), .C2(new_n919_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT62), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n866_), .A2(new_n916_), .ZN(new_n922_));
  OAI211_X1 g721(.A(new_n921_), .B(G169gat), .C1(new_n922_), .C2(new_n653_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n920_), .A2(new_n923_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(KEYINPUT127), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT127), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n920_), .A2(new_n926_), .A3(new_n923_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n925_), .A2(new_n927_), .ZN(G1348gat));
  NAND4_X1  g727(.A1(new_n894_), .A2(G176gat), .A3(new_n732_), .A4(new_n916_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n378_), .B1(new_n922_), .B2(new_n874_), .ZN(new_n930_));
  AND2_X1   g729(.A1(new_n929_), .A2(new_n930_), .ZN(G1349gat));
  NOR2_X1   g730(.A1(new_n922_), .A2(new_n642_), .ZN(new_n932_));
  MUX2_X1   g731(.A(G183gat), .B(new_n374_), .S(new_n932_), .Z(G1350gat));
  OAI21_X1  g732(.A(G190gat), .B1(new_n922_), .B2(new_n851_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n617_), .A2(new_n375_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n934_), .B1(new_n922_), .B2(new_n935_), .ZN(G1351gat));
  NAND4_X1  g735(.A1(new_n894_), .A2(new_n565_), .A3(new_n520_), .A4(new_n914_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(G197gat), .ZN(G1352gat));
  NAND4_X1  g737(.A1(new_n894_), .A2(new_n520_), .A3(new_n732_), .A4(new_n914_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n939_), .B(G204gat), .ZN(G1353gat));
  NAND4_X1  g739(.A1(new_n894_), .A2(new_n693_), .A3(new_n520_), .A4(new_n914_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n942_));
  AND2_X1   g741(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n943_));
  NOR3_X1   g742(.A1(new_n941_), .A2(new_n942_), .A3(new_n943_), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n944_), .B1(new_n941_), .B2(new_n942_), .ZN(G1354gat));
  AND3_X1   g744(.A1(new_n894_), .A2(new_n520_), .A3(new_n914_), .ZN(new_n946_));
  AOI21_X1  g745(.A(G218gat), .B1(new_n946_), .B2(new_n617_), .ZN(new_n947_));
  INV_X1    g746(.A(G218gat), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n851_), .A2(new_n948_), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n947_), .B1(new_n946_), .B2(new_n949_), .ZN(G1355gat));
endmodule


