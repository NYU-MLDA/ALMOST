//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 0 1 1 0 1 1 0 1 1 1 0 0 1 1 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 1 0 0 1 1 1 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n675_, new_n676_, new_n677_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n751_, new_n752_,
    new_n753_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n766_,
    new_n767_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n893_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n918_, new_n919_, new_n921_, new_n922_, new_n924_, new_n925_,
    new_n926_, new_n928_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n935_, new_n936_, new_n937_;
  INV_X1    g000(.A(KEYINPUT4), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT89), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G127gat), .B(G134gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(G113gat), .B(G120gat), .Z(new_n206_));
  AOI21_X1  g005(.A(new_n203_), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G113gat), .B(G120gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n204_), .A2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n207_), .B(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(KEYINPUT91), .A2(KEYINPUT3), .ZN(new_n211_));
  INV_X1    g010(.A(G141gat), .ZN(new_n212_));
  INV_X1    g011(.A(G148gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G141gat), .A2(G148gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT2), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  OAI22_X1  g016(.A1(KEYINPUT91), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n214_), .A2(new_n217_), .A3(new_n218_), .A4(new_n219_), .ZN(new_n220_));
  OR2_X1    g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G155gat), .A2(G162gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n220_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n212_), .A2(new_n213_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n222_), .A2(KEYINPUT1), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(new_n221_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n222_), .A2(KEYINPUT1), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n224_), .B(new_n215_), .C1(new_n226_), .C2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n223_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n210_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n205_), .A2(new_n206_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(new_n209_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT101), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n231_), .A2(KEYINPUT101), .A3(new_n209_), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n234_), .A2(new_n223_), .A3(new_n228_), .A4(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n202_), .B1(new_n230_), .B2(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(KEYINPUT4), .B1(new_n210_), .B2(new_n229_), .ZN(new_n238_));
  OAI211_X1 g037(.A(G225gat), .B(G233gat), .C1(new_n237_), .C2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G225gat), .A2(G233gat), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n230_), .A2(new_n240_), .A3(new_n236_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G1gat), .B(G29gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(G85gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT0), .B(G57gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n239_), .A2(new_n241_), .A3(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT102), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n239_), .A2(new_n241_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(new_n245_), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n239_), .A2(new_n241_), .A3(KEYINPUT102), .A4(new_n246_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n249_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT20), .ZN(new_n255_));
  XOR2_X1   g054(.A(G211gat), .B(G218gat), .Z(new_n256_));
  XOR2_X1   g055(.A(G197gat), .B(G204gat), .Z(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT21), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT93), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n256_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G197gat), .B(G204gat), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT21), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n261_), .A2(KEYINPUT94), .A3(new_n262_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n261_), .A2(new_n262_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT93), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT94), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n266_), .B1(new_n257_), .B2(KEYINPUT21), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n260_), .A2(new_n263_), .A3(new_n265_), .A4(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT95), .ZN(new_n269_));
  OR2_X1    g068(.A1(new_n256_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n256_), .A2(new_n269_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n270_), .A2(new_n264_), .A3(new_n271_), .ZN(new_n272_));
  AND2_X1   g071(.A1(new_n268_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT23), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n274_), .B1(G183gat), .B2(G190gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G183gat), .A2(G190gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT87), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n275_), .B1(new_n277_), .B2(new_n274_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(G183gat), .A2(G190gat), .ZN(new_n279_));
  OR2_X1    g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(G169gat), .ZN(new_n281_));
  INV_X1    g080(.A(G176gat), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT22), .B(G169gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT98), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n283_), .B1(new_n285_), .B2(new_n282_), .ZN(new_n286_));
  AOI21_X1  g085(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n287_), .B1(new_n277_), .B2(KEYINPUT23), .ZN(new_n288_));
  NOR3_X1   g087(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n289_));
  INV_X1    g088(.A(new_n283_), .ZN(new_n290_));
  OAI21_X1  g089(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n289_), .B1(new_n290_), .B2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT26), .B(G190gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT25), .B(G183gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  AND2_X1   g095(.A1(new_n293_), .A2(new_n296_), .ZN(new_n297_));
  AOI22_X1  g096(.A1(new_n280_), .A2(new_n286_), .B1(new_n288_), .B2(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n255_), .B1(new_n273_), .B2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G226gat), .A2(G233gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT19), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n268_), .A2(new_n272_), .ZN(new_n303_));
  AOI211_X1 g102(.A(new_n279_), .B(new_n287_), .C1(new_n277_), .C2(KEYINPUT23), .ZN(new_n304_));
  NOR2_X1   g103(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(new_n281_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT86), .ZN(new_n307_));
  INV_X1    g106(.A(G183gat), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT25), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  OR2_X1    g108(.A1(new_n308_), .A2(KEYINPUT25), .ZN(new_n310_));
  OAI211_X1 g109(.A(new_n294_), .B(new_n309_), .C1(new_n310_), .C2(new_n307_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(new_n293_), .ZN(new_n312_));
  OAI22_X1  g111(.A1(new_n304_), .A2(new_n306_), .B1(new_n312_), .B2(new_n278_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n303_), .A2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n299_), .A2(new_n302_), .A3(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(KEYINPUT100), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT100), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n299_), .A2(new_n317_), .A3(new_n302_), .A4(new_n314_), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT20), .B1(new_n303_), .B2(new_n313_), .ZN(new_n319_));
  OAI21_X1  g118(.A(KEYINPUT99), .B1(new_n273_), .B2(new_n298_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT99), .ZN(new_n321_));
  AND2_X1   g120(.A1(new_n280_), .A2(new_n286_), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n297_), .A2(new_n288_), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n321_), .B(new_n303_), .C1(new_n322_), .C2(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n319_), .B1(new_n320_), .B2(new_n324_), .ZN(new_n325_));
  XOR2_X1   g124(.A(new_n301_), .B(KEYINPUT97), .Z(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n316_), .B(new_n318_), .C1(new_n325_), .C2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G8gat), .B(G36gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT18), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G64gat), .B(G92gat), .ZN(new_n331_));
  XOR2_X1   g130(.A(new_n330_), .B(new_n331_), .Z(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n328_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n320_), .A2(new_n324_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n319_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(new_n326_), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n338_), .A2(new_n332_), .A3(new_n316_), .A4(new_n318_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n334_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT27), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  XOR2_X1   g141(.A(G71gat), .B(G99gat), .Z(new_n343_));
  XNOR2_X1  g142(.A(G15gat), .B(G43gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n313_), .B(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(new_n210_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G227gat), .A2(G233gat), .ZN(new_n349_));
  XOR2_X1   g148(.A(new_n349_), .B(KEYINPUT88), .Z(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT30), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT31), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n346_), .A2(new_n210_), .ZN(new_n354_));
  OR3_X1    g153(.A1(new_n348_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n353_), .B1(new_n348_), .B2(new_n354_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G228gat), .A2(G233gat), .ZN(new_n358_));
  INV_X1    g157(.A(G78gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(G106gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n229_), .A2(KEYINPUT29), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n303_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n362_), .B1(new_n303_), .B2(new_n363_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n361_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n366_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n368_), .A2(new_n360_), .A3(new_n364_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT92), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n367_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(KEYINPUT96), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT96), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n367_), .A2(new_n369_), .A3(new_n373_), .ZN(new_n374_));
  OR2_X1    g173(.A1(new_n229_), .A2(KEYINPUT29), .ZN(new_n375_));
  OR2_X1    g174(.A1(new_n375_), .A2(KEYINPUT28), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(KEYINPUT28), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  XOR2_X1   g177(.A(G22gat), .B(G50gat), .Z(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n379_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n376_), .A2(new_n381_), .A3(new_n377_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n372_), .A2(new_n374_), .A3(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n371_), .A2(KEYINPUT96), .A3(new_n383_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n357_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT103), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n388_), .B1(new_n328_), .B2(new_n333_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n273_), .A2(new_n298_), .ZN(new_n390_));
  AND4_X1   g189(.A1(KEYINPUT20), .A2(new_n390_), .A3(new_n302_), .A4(new_n314_), .ZN(new_n391_));
  AOI22_X1  g190(.A1(new_n337_), .A2(new_n326_), .B1(new_n391_), .B2(new_n317_), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n392_), .A2(KEYINPUT103), .A3(new_n332_), .A4(new_n316_), .ZN(new_n393_));
  AND2_X1   g192(.A1(new_n299_), .A2(new_n314_), .ZN(new_n394_));
  OAI22_X1  g193(.A1(new_n337_), .A2(new_n326_), .B1(new_n394_), .B2(new_n302_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n341_), .B1(new_n395_), .B2(new_n333_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n389_), .A2(new_n393_), .A3(new_n396_), .ZN(new_n397_));
  AND4_X1   g196(.A1(new_n254_), .A2(new_n342_), .A3(new_n387_), .A4(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n230_), .A2(new_n236_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n245_), .B1(new_n399_), .B2(new_n240_), .ZN(new_n400_));
  OR2_X1    g199(.A1(new_n237_), .A2(new_n238_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n400_), .B1(new_n401_), .B2(new_n240_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT33), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n247_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  OR2_X1    g203(.A1(new_n247_), .A2(new_n403_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n334_), .A2(new_n339_), .A3(new_n404_), .A4(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n395_), .A2(KEYINPUT32), .A3(new_n332_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n332_), .A2(KEYINPUT32), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n338_), .A2(new_n316_), .A3(new_n318_), .A4(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n253_), .A2(new_n407_), .A3(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n406_), .A2(new_n410_), .ZN(new_n411_));
  AND3_X1   g210(.A1(new_n371_), .A2(KEYINPUT96), .A3(new_n383_), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n384_), .A2(new_n374_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n412_), .B1(new_n413_), .B2(new_n372_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n411_), .A2(new_n415_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n342_), .A2(new_n397_), .A3(new_n254_), .A4(new_n414_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n357_), .B(KEYINPUT90), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n398_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G229gat), .A2(G233gat), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT14), .ZN(new_n422_));
  XOR2_X1   g221(.A(KEYINPUT80), .B(G1gat), .Z(new_n423_));
  XOR2_X1   g222(.A(KEYINPUT81), .B(G8gat), .Z(new_n424_));
  AOI21_X1  g223(.A(new_n422_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  XOR2_X1   g224(.A(G15gat), .B(G22gat), .Z(new_n426_));
  XNOR2_X1  g225(.A(G1gat), .B(G8gat), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  OR3_X1    g227(.A1(new_n425_), .A2(new_n426_), .A3(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n428_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G29gat), .B(G36gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT75), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G43gat), .B(G50gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n431_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n434_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n433_), .B(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(KEYINPUT15), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n421_), .B(new_n436_), .C1(new_n439_), .C2(new_n431_), .ZN(new_n440_));
  AOI21_X1  g239(.A(KEYINPUT84), .B1(new_n431_), .B2(new_n435_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n441_), .B1(new_n435_), .B2(new_n431_), .ZN(new_n442_));
  AND2_X1   g241(.A1(new_n429_), .A2(new_n430_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n443_), .A2(KEYINPUT84), .A3(new_n438_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n421_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n442_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n440_), .A2(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G113gat), .B(G141gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G169gat), .B(G197gat), .ZN(new_n449_));
  XOR2_X1   g248(.A(new_n448_), .B(new_n449_), .Z(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n447_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT85), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n440_), .A2(new_n446_), .A3(new_n450_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n452_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n447_), .A2(KEYINPUT85), .A3(new_n451_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT104), .B1(new_n420_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT104), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n455_), .A2(new_n456_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n419_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n461_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n459_), .B(new_n460_), .C1(new_n462_), .C2(new_n398_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT13), .ZN(new_n464_));
  XNOR2_X1  g263(.A(KEYINPUT69), .B(G71gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(new_n359_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G57gat), .B(G64gat), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n467_), .A2(KEYINPUT11), .ZN(new_n468_));
  OR2_X1    g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n467_), .A2(KEYINPUT11), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n466_), .B1(new_n468_), .B2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT12), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT6), .ZN(new_n476_));
  AND3_X1   g275(.A1(KEYINPUT65), .A2(G99gat), .A3(G106gat), .ZN(new_n477_));
  AOI21_X1  g276(.A(KEYINPUT65), .B1(G99gat), .B2(G106gat), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n476_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G99gat), .A2(G106gat), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT65), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(KEYINPUT65), .A2(G99gat), .A3(G106gat), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n482_), .A2(KEYINPUT6), .A3(new_n483_), .ZN(new_n484_));
  OR2_X1    g283(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n485_), .A2(new_n362_), .A3(new_n486_), .ZN(new_n487_));
  AND3_X1   g286(.A1(new_n479_), .A2(new_n484_), .A3(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G85gat), .A2(G92gat), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(G85gat), .A2(G92gat), .ZN(new_n491_));
  INV_X1    g290(.A(G92gat), .ZN(new_n492_));
  OAI22_X1  g291(.A1(new_n490_), .A2(new_n491_), .B1(KEYINPUT9), .B2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n491_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT9), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n494_), .A2(new_n495_), .A3(new_n489_), .ZN(new_n496_));
  AND3_X1   g295(.A1(new_n493_), .A2(new_n496_), .A3(KEYINPUT64), .ZN(new_n497_));
  AOI21_X1  g296(.A(KEYINPUT64), .B1(new_n493_), .B2(new_n496_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n488_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT67), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n501_), .A2(KEYINPUT6), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n476_), .A2(KEYINPUT67), .ZN(new_n503_));
  OAI22_X1  g302(.A1(new_n502_), .A2(new_n503_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n504_));
  OR2_X1    g303(.A1(G99gat), .A2(G106gat), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT7), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n506_), .A2(KEYINPUT66), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT66), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n508_), .A2(KEYINPUT7), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n505_), .B1(new_n507_), .B2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n476_), .A2(KEYINPUT67), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n501_), .A2(KEYINPUT6), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n482_), .A2(new_n483_), .A3(new_n511_), .A4(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n508_), .A2(KEYINPUT7), .ZN(new_n514_));
  NOR2_X1   g313(.A1(G99gat), .A2(G106gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n504_), .A2(new_n510_), .A3(new_n513_), .A4(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n490_), .A2(new_n491_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT8), .ZN(new_n520_));
  AND2_X1   g319(.A1(new_n479_), .A2(new_n484_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n516_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n506_), .A2(KEYINPUT66), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n515_), .B1(new_n514_), .B2(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n521_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT8), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n518_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n526_), .A2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n520_), .A2(KEYINPUT70), .A3(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT70), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n527_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n528_), .B1(new_n521_), .B2(new_n525_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n532_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n500_), .B1(new_n531_), .B2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT71), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  AOI211_X1 g337(.A(KEYINPUT71), .B(new_n500_), .C1(new_n531_), .C2(new_n535_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n475_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G230gat), .A2(G233gat), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n499_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT68), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  OAI211_X1 g343(.A(new_n499_), .B(KEYINPUT68), .C1(new_n533_), .C2(new_n534_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n472_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n544_), .A2(new_n545_), .A3(new_n472_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n546_), .B1(new_n474_), .B2(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n540_), .A2(new_n541_), .A3(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n544_), .A2(new_n545_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(new_n473_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(new_n547_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n541_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n549_), .A2(new_n554_), .ZN(new_n555_));
  XOR2_X1   g354(.A(G120gat), .B(G148gat), .Z(new_n556_));
  XNOR2_X1  g355(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  XOR2_X1   g357(.A(G176gat), .B(G204gat), .Z(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  AND2_X1   g359(.A1(new_n560_), .A2(KEYINPUT72), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n555_), .A2(new_n561_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n555_), .A2(new_n561_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n464_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n555_), .A2(new_n561_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n555_), .A2(new_n561_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n565_), .A2(KEYINPUT13), .A3(new_n566_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n564_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(KEYINPUT74), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n564_), .A2(new_n567_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT74), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n569_), .A2(new_n572_), .ZN(new_n573_));
  AND3_X1   g372(.A1(new_n458_), .A2(new_n463_), .A3(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G232gat), .A2(G233gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT34), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT35), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(KEYINPUT70), .B1(new_n520_), .B2(new_n530_), .ZN(new_n580_));
  NOR3_X1   g379(.A1(new_n533_), .A2(new_n534_), .A3(new_n532_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n499_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(KEYINPUT71), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n536_), .A2(new_n537_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n439_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  AOI22_X1  g384(.A1(new_n550_), .A2(new_n435_), .B1(new_n578_), .B2(new_n577_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n579_), .B1(new_n585_), .B2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n439_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n589_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n579_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n590_), .A2(new_n591_), .A3(new_n586_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G190gat), .B(G218gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT76), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G134gat), .B(G162gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT36), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  XOR2_X1   g397(.A(KEYINPUT77), .B(KEYINPUT78), .Z(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n588_), .A2(new_n592_), .A3(new_n600_), .ZN(new_n601_));
  AND2_X1   g400(.A1(new_n588_), .A2(new_n592_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n596_), .B(new_n597_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT79), .ZN(new_n604_));
  OAI211_X1 g403(.A(KEYINPUT37), .B(new_n601_), .C1(new_n602_), .C2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT37), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n588_), .A2(new_n592_), .A3(new_n600_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n604_), .B1(new_n588_), .B2(new_n592_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n606_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n605_), .A2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n431_), .A2(G231gat), .A3(G233gat), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n431_), .B1(G231gat), .B2(G233gat), .ZN(new_n613_));
  NOR3_X1   g412(.A1(new_n612_), .A2(new_n613_), .A3(new_n473_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G127gat), .B(G155gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G183gat), .B(G211gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n473_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n615_), .A2(KEYINPUT17), .A3(new_n620_), .A4(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT83), .ZN(new_n623_));
  INV_X1    g422(.A(new_n621_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n624_), .A2(new_n614_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n620_), .B(KEYINPUT17), .ZN(new_n626_));
  OAI211_X1 g425(.A(new_n622_), .B(new_n623_), .C1(new_n625_), .C2(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n626_), .B1(new_n615_), .B2(new_n621_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n620_), .A2(KEYINPUT17), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n624_), .A2(new_n614_), .A3(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(KEYINPUT83), .B1(new_n628_), .B2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n627_), .A2(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n610_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n574_), .A2(new_n633_), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n254_), .A2(KEYINPUT105), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n254_), .A2(KEYINPUT105), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  OR3_X1    g436(.A1(new_n634_), .A2(new_n423_), .A3(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n607_), .A2(new_n608_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n420_), .A2(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n628_), .A2(new_n630_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n457_), .B1(new_n569_), .B2(new_n572_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n642_), .A2(new_n643_), .A3(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(G1gat), .B1(new_n645_), .B2(new_n254_), .ZN(new_n646_));
  AND3_X1   g445(.A1(new_n638_), .A2(KEYINPUT107), .A3(new_n639_), .ZN(new_n647_));
  AOI21_X1  g446(.A(KEYINPUT107), .B1(new_n638_), .B2(new_n639_), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n640_), .B(new_n646_), .C1(new_n647_), .C2(new_n648_), .ZN(G1324gat));
  XNOR2_X1  g448(.A(KEYINPUT109), .B(KEYINPUT40), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n342_), .A2(new_n397_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n642_), .A2(new_n643_), .A3(new_n644_), .A4(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT39), .ZN(new_n654_));
  AND4_X1   g453(.A1(KEYINPUT108), .A2(new_n653_), .A3(new_n654_), .A4(G8gat), .ZN(new_n655_));
  OAI21_X1  g454(.A(G8gat), .B1(new_n654_), .B2(KEYINPUT108), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  AOI22_X1  g456(.A1(new_n653_), .A2(new_n657_), .B1(KEYINPUT108), .B2(new_n654_), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n655_), .A2(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n651_), .A2(new_n424_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n574_), .A2(new_n633_), .A3(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n650_), .B1(new_n659_), .B2(new_n661_), .ZN(new_n662_));
  OAI211_X1 g461(.A(new_n661_), .B(new_n650_), .C1(new_n655_), .C2(new_n658_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n662_), .A2(new_n664_), .ZN(G1325gat));
  OR3_X1    g464(.A1(new_n634_), .A2(G15gat), .A3(new_n419_), .ZN(new_n666_));
  OR2_X1    g465(.A1(new_n645_), .A2(new_n419_), .ZN(new_n667_));
  AND3_X1   g466(.A1(new_n667_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n668_));
  AOI21_X1  g467(.A(KEYINPUT41), .B1(new_n667_), .B2(G15gat), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n666_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT110), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  OAI211_X1 g471(.A(new_n666_), .B(KEYINPUT110), .C1(new_n668_), .C2(new_n669_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1326gat));
  OAI21_X1  g473(.A(G22gat), .B1(new_n645_), .B2(new_n415_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT42), .ZN(new_n676_));
  OR2_X1    g475(.A1(new_n415_), .A2(G22gat), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n676_), .B1(new_n634_), .B2(new_n677_), .ZN(G1327gat));
  NAND2_X1  g477(.A1(new_n641_), .A2(new_n632_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT112), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n458_), .A2(new_n463_), .A3(new_n573_), .A4(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(G29gat), .B1(new_n682_), .B2(new_n253_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n632_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n610_), .B1(new_n462_), .B2(new_n398_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n610_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT111), .ZN(new_n687_));
  OAI21_X1  g486(.A(KEYINPUT43), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n684_), .B1(new_n685_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT43), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n690_), .B1(new_n610_), .B2(KEYINPUT111), .ZN(new_n691_));
  OAI211_X1 g490(.A(new_n610_), .B(new_n691_), .C1(new_n462_), .C2(new_n398_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n689_), .A2(new_n692_), .A3(new_n644_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  NAND4_X1  g494(.A1(new_n689_), .A2(new_n692_), .A3(KEYINPUT44), .A4(new_n644_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n637_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n698_), .A2(G29gat), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n683_), .B1(new_n697_), .B2(new_n699_), .ZN(G1328gat));
  NAND3_X1  g499(.A1(new_n695_), .A2(new_n652_), .A3(new_n696_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(G36gat), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT113), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n651_), .A2(G36gat), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n574_), .A2(new_n703_), .A3(new_n680_), .A4(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT45), .ZN(new_n706_));
  INV_X1    g505(.A(new_n704_), .ZN(new_n707_));
  OAI21_X1  g506(.A(KEYINPUT113), .B1(new_n681_), .B2(new_n707_), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n705_), .A2(new_n706_), .A3(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n706_), .B1(new_n705_), .B2(new_n708_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n702_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT46), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n702_), .B(KEYINPUT46), .C1(new_n709_), .C2(new_n710_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(G1329gat));
  INV_X1    g514(.A(G43gat), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n357_), .A2(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n695_), .A2(new_n696_), .A3(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT114), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n682_), .A2(new_n461_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(new_n720_), .B2(new_n716_), .ZN(new_n721_));
  AOI211_X1 g520(.A(KEYINPUT114), .B(G43gat), .C1(new_n682_), .C2(new_n461_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n718_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(KEYINPUT47), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT47), .ZN(new_n725_));
  OAI211_X1 g524(.A(new_n725_), .B(new_n718_), .C1(new_n721_), .C2(new_n722_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(G1330gat));
  AOI21_X1  g526(.A(G50gat), .B1(new_n682_), .B2(new_n414_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n414_), .A2(G50gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n697_), .B2(new_n729_), .ZN(G1331gat));
  AND2_X1   g529(.A1(new_n569_), .A2(new_n572_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n460_), .A2(new_n632_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n642_), .A2(new_n731_), .A3(new_n732_), .ZN(new_n733_));
  OAI21_X1  g532(.A(G57gat), .B1(new_n733_), .B2(new_n254_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n731_), .A2(KEYINPUT115), .A3(new_n633_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT115), .ZN(new_n736_));
  INV_X1    g535(.A(new_n633_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n736_), .B1(new_n573_), .B2(new_n737_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n420_), .A2(new_n460_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n735_), .A2(new_n738_), .A3(new_n739_), .ZN(new_n740_));
  OR2_X1    g539(.A1(new_n637_), .A2(G57gat), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n734_), .B1(new_n740_), .B2(new_n741_), .ZN(G1332gat));
  OAI21_X1  g541(.A(G64gat), .B1(new_n733_), .B2(new_n651_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT48), .ZN(new_n744_));
  OR2_X1    g543(.A1(new_n651_), .A2(G64gat), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n744_), .B1(new_n740_), .B2(new_n745_), .ZN(G1333gat));
  OAI21_X1  g545(.A(G71gat), .B1(new_n733_), .B2(new_n419_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT49), .ZN(new_n748_));
  OR2_X1    g547(.A1(new_n419_), .A2(G71gat), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n748_), .B1(new_n740_), .B2(new_n749_), .ZN(G1334gat));
  OAI21_X1  g549(.A(G78gat), .B1(new_n733_), .B2(new_n415_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT50), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n414_), .A2(new_n359_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n752_), .B1(new_n740_), .B2(new_n753_), .ZN(G1335gat));
  NOR2_X1   g553(.A1(new_n573_), .A2(new_n460_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n689_), .A2(new_n692_), .A3(new_n755_), .ZN(new_n756_));
  OAI21_X1  g555(.A(G85gat), .B1(new_n756_), .B2(new_n254_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n739_), .A2(new_n731_), .A3(new_n680_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT116), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT116), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n739_), .A2(new_n731_), .A3(new_n760_), .A4(new_n680_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  OR2_X1    g562(.A1(new_n637_), .A2(G85gat), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n757_), .B1(new_n763_), .B2(new_n764_), .ZN(G1336gat));
  OAI21_X1  g564(.A(G92gat), .B1(new_n756_), .B2(new_n651_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n652_), .A2(new_n492_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n766_), .B1(new_n763_), .B2(new_n767_), .ZN(G1337gat));
  OAI21_X1  g567(.A(G99gat), .B1(new_n756_), .B2(new_n419_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT117), .ZN(new_n770_));
  AND4_X1   g569(.A1(new_n485_), .A2(new_n355_), .A3(new_n486_), .A4(new_n356_), .ZN(new_n771_));
  AND3_X1   g570(.A1(new_n762_), .A2(new_n770_), .A3(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n770_), .B1(new_n762_), .B2(new_n771_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n769_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n774_), .A2(KEYINPUT118), .A3(KEYINPUT51), .ZN(new_n775_));
  NAND2_X1  g574(.A1(KEYINPUT118), .A2(KEYINPUT51), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n776_), .B(new_n769_), .C1(new_n772_), .C2(new_n773_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(G1338gat));
  NAND3_X1  g577(.A1(new_n762_), .A2(new_n362_), .A3(new_n414_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n689_), .A2(new_n692_), .A3(new_n414_), .A4(new_n755_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT52), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n780_), .A2(new_n781_), .A3(G106gat), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n781_), .B1(new_n780_), .B2(G106gat), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n779_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT53), .ZN(G1339gat));
  AND4_X1   g584(.A1(new_n609_), .A2(new_n605_), .A3(new_n684_), .A4(new_n457_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT119), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT54), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n786_), .A2(new_n568_), .A3(new_n787_), .A4(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n786_), .A2(new_n788_), .A3(new_n568_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT119), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n732_), .A2(new_n609_), .A3(new_n605_), .ZN(new_n792_));
  OAI21_X1  g591(.A(KEYINPUT54), .B1(new_n792_), .B2(new_n570_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT120), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT120), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n795_), .B(KEYINPUT54), .C1(new_n792_), .C2(new_n570_), .ZN(new_n796_));
  AOI22_X1  g595(.A1(new_n789_), .A2(new_n791_), .B1(new_n794_), .B2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n641_), .ZN(new_n798_));
  OR2_X1    g597(.A1(new_n555_), .A2(new_n560_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n460_), .A2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n475_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n801_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n547_), .A2(new_n474_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n551_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n553_), .B1(new_n802_), .B2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT121), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT55), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n549_), .A2(new_n807_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n540_), .A2(new_n548_), .A3(KEYINPUT55), .A4(new_n541_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT121), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n810_), .B(new_n553_), .C1(new_n802_), .C2(new_n804_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n806_), .A2(new_n808_), .A3(new_n809_), .A4(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n560_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT56), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n812_), .A2(KEYINPUT56), .A3(new_n560_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n800_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n442_), .A2(new_n444_), .A3(new_n421_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n439_), .A2(new_n431_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n436_), .A2(new_n445_), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n818_), .B(new_n451_), .C1(new_n819_), .C2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n454_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n822_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n798_), .B1(new_n817_), .B2(new_n823_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(KEYINPUT122), .A2(KEYINPUT57), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n800_), .ZN(new_n827_));
  AND3_X1   g626(.A1(new_n812_), .A2(KEYINPUT56), .A3(new_n560_), .ZN(new_n828_));
  AOI21_X1  g627(.A(KEYINPUT56), .B1(new_n812_), .B2(new_n560_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n827_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n823_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n641_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n825_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT123), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n835_), .A2(KEYINPUT58), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n815_), .A2(new_n816_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n822_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n799_), .A2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n837_), .B1(new_n838_), .B2(new_n841_), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n837_), .B(new_n841_), .C1(new_n828_), .C2(new_n829_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n610_), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n826_), .B(new_n834_), .C1(new_n842_), .C2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n643_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n797_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n698_), .A2(new_n651_), .A3(new_n387_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(G113gat), .B1(new_n849_), .B2(new_n460_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT59), .ZN(new_n851_));
  OAI22_X1  g650(.A1(new_n832_), .A2(new_n833_), .B1(new_n844_), .B2(new_n842_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n824_), .A2(new_n825_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n846_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n791_), .A2(new_n789_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n794_), .A2(new_n796_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n854_), .A2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n848_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n851_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n851_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n845_), .A2(new_n632_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n861_), .B1(new_n862_), .B2(new_n857_), .ZN(new_n863_));
  OAI21_X1  g662(.A(KEYINPUT124), .B1(new_n860_), .B2(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(KEYINPUT59), .B1(new_n847_), .B2(new_n848_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT124), .ZN(new_n866_));
  INV_X1    g665(.A(new_n844_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n842_), .ZN(new_n868_));
  AOI22_X1  g667(.A1(new_n867_), .A2(new_n868_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n684_), .B1(new_n869_), .B2(new_n834_), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n851_), .B(new_n859_), .C1(new_n870_), .C2(new_n797_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n865_), .A2(new_n866_), .A3(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n864_), .A2(new_n872_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n460_), .A2(G113gat), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n850_), .B1(new_n873_), .B2(new_n874_), .ZN(G1340gat));
  INV_X1    g674(.A(G120gat), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n876_), .B1(new_n573_), .B2(KEYINPUT60), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n849_), .B(new_n877_), .C1(KEYINPUT60), .C2(new_n876_), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n860_), .A2(new_n863_), .A3(new_n573_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n879_), .B2(new_n876_), .ZN(G1341gat));
  AOI21_X1  g679(.A(G127gat), .B1(new_n849_), .B2(new_n684_), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n643_), .A2(G127gat), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n881_), .B1(new_n873_), .B2(new_n882_), .ZN(G1342gat));
  AOI21_X1  g682(.A(G134gat), .B1(new_n849_), .B2(new_n641_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(KEYINPUT125), .B(G134gat), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n686_), .A2(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n884_), .B1(new_n873_), .B2(new_n886_), .ZN(G1343gat));
  NAND4_X1  g686(.A1(new_n698_), .A2(new_n414_), .A3(new_n651_), .A4(new_n419_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(KEYINPUT126), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n847_), .A2(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(new_n460_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g691(.A1(new_n890_), .A2(new_n731_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g693(.A1(new_n890_), .A2(new_n684_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(KEYINPUT61), .B(G155gat), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n895_), .B(new_n896_), .ZN(G1346gat));
  INV_X1    g696(.A(new_n890_), .ZN(new_n898_));
  OR3_X1    g697(.A1(new_n898_), .A2(G162gat), .A3(new_n798_), .ZN(new_n899_));
  OAI21_X1  g698(.A(G162gat), .B1(new_n898_), .B2(new_n686_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(G1347gat));
  XNOR2_X1  g700(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n698_), .A2(new_n419_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n652_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n904_), .A2(new_n414_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n905_), .B1(new_n870_), .B2(new_n797_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n906_), .A2(new_n457_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n902_), .B1(new_n907_), .B2(new_n281_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n902_), .ZN(new_n909_));
  OAI211_X1 g708(.A(G169gat), .B(new_n909_), .C1(new_n906_), .C2(new_n457_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n907_), .A2(new_n285_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n908_), .A2(new_n910_), .A3(new_n911_), .ZN(G1348gat));
  INV_X1    g711(.A(new_n906_), .ZN(new_n913_));
  AOI21_X1  g712(.A(G176gat), .B1(new_n913_), .B2(new_n731_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n847_), .A2(new_n414_), .ZN(new_n915_));
  NOR3_X1   g714(.A1(new_n904_), .A2(new_n573_), .A3(new_n282_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n914_), .B1(new_n915_), .B2(new_n916_), .ZN(G1349gat));
  NOR3_X1   g716(.A1(new_n906_), .A2(new_n846_), .A3(new_n295_), .ZN(new_n918_));
  NAND4_X1  g717(.A1(new_n915_), .A2(new_n684_), .A3(new_n652_), .A4(new_n903_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n918_), .B1(new_n919_), .B2(new_n308_), .ZN(G1350gat));
  OAI21_X1  g719(.A(G190gat), .B1(new_n906_), .B2(new_n686_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n641_), .A2(new_n294_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n921_), .B1(new_n906_), .B2(new_n922_), .ZN(G1351gat));
  NAND4_X1  g722(.A1(new_n652_), .A2(new_n254_), .A3(new_n414_), .A4(new_n419_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n847_), .A2(new_n924_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(new_n460_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g726(.A1(new_n925_), .A2(new_n731_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g728(.A1(new_n925_), .A2(new_n643_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(KEYINPUT63), .B(G211gat), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n930_), .A2(new_n931_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n932_), .B1(new_n930_), .B2(new_n933_), .ZN(G1354gat));
  INV_X1    g733(.A(G218gat), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n925_), .A2(new_n935_), .A3(new_n641_), .ZN(new_n936_));
  NOR3_X1   g735(.A1(new_n847_), .A2(new_n686_), .A3(new_n924_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n936_), .B1(new_n937_), .B2(new_n935_), .ZN(G1355gat));
endmodule


