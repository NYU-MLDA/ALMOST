//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 0 0 1 0 0 1 0 1 1 1 0 0 0 0 1 1 0 1 0 1 0 0 0 0 0 1 1 1 1 0 1 1 0 1 1 1 0 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n810_, new_n811_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n832_, new_n833_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n842_, new_n843_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_,
    new_n859_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n936_, new_n937_, new_n939_, new_n940_, new_n942_,
    new_n944_, new_n945_, new_n946_, new_n948_, new_n949_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n961_, new_n962_, new_n963_, new_n964_,
    new_n966_, new_n968_, new_n969_, new_n970_, new_n971_, new_n972_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n983_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n990_, new_n991_, new_n992_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT81), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT81), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n204_), .A2(G183gat), .A3(G190gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n205_), .A3(KEYINPUT23), .ZN(new_n206_));
  OR2_X1    g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT23), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n202_), .A2(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n206_), .A2(new_n207_), .A3(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT22), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(G169gat), .ZN(new_n213_));
  NOR3_X1   g012(.A1(new_n213_), .A2(KEYINPUT82), .A3(KEYINPUT83), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT82), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n212_), .A2(G169gat), .ZN(new_n216_));
  INV_X1    g015(.A(G169gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n217_), .A2(KEYINPUT22), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n215_), .B1(new_n216_), .B2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT83), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n217_), .A2(KEYINPUT22), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n220_), .B1(new_n221_), .B2(KEYINPUT82), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n214_), .B1(new_n219_), .B2(new_n222_), .ZN(new_n223_));
  XOR2_X1   g022(.A(KEYINPUT84), .B(G176gat), .Z(new_n224_));
  OAI211_X1 g023(.A(new_n210_), .B(new_n211_), .C1(new_n223_), .C2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT30), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT26), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(G190gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT80), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  AND2_X1   g029(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n231_));
  NOR2_X1   g030(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(G190gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT26), .ZN(new_n235_));
  AND2_X1   g034(.A1(new_n228_), .A2(new_n235_), .ZN(new_n236_));
  OAI211_X1 g035(.A(new_n230_), .B(new_n233_), .C1(new_n236_), .C2(new_n229_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n203_), .A2(new_n205_), .A3(new_n208_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n202_), .A2(KEYINPUT23), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(G176gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n217_), .A2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n242_), .A2(KEYINPUT24), .A3(new_n211_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n242_), .A2(KEYINPUT24), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n237_), .A2(new_n240_), .A3(new_n243_), .A4(new_n245_), .ZN(new_n246_));
  AND3_X1   g045(.A1(new_n225_), .A2(new_n226_), .A3(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n226_), .B1(new_n225_), .B2(new_n246_), .ZN(new_n248_));
  OAI21_X1  g047(.A(KEYINPUT87), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n225_), .A2(new_n246_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT30), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT87), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n225_), .A2(new_n226_), .A3(new_n246_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n251_), .A2(new_n252_), .A3(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G227gat), .A2(G233gat), .ZN(new_n255_));
  XOR2_X1   g054(.A(new_n255_), .B(KEYINPUT85), .Z(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT86), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G71gat), .B(G99gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G15gat), .B(G43gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n257_), .B(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n249_), .A2(new_n254_), .A3(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n261_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n247_), .A2(new_n248_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n263_), .A2(new_n264_), .A3(new_n252_), .ZN(new_n265_));
  OR2_X1    g064(.A1(G127gat), .A2(G134gat), .ZN(new_n266_));
  INV_X1    g065(.A(G113gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G127gat), .A2(G134gat), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n266_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n269_));
  AND2_X1   g068(.A1(G127gat), .A2(G134gat), .ZN(new_n270_));
  NOR2_X1   g069(.A1(G127gat), .A2(G134gat), .ZN(new_n271_));
  OAI21_X1  g070(.A(G113gat), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  AND3_X1   g071(.A1(new_n269_), .A2(new_n272_), .A3(G120gat), .ZN(new_n273_));
  AOI21_X1  g072(.A(G120gat), .B1(new_n269_), .B2(new_n272_), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT31), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n273_), .A2(new_n274_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT31), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT88), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  AND3_X1   g081(.A1(new_n262_), .A2(new_n265_), .A3(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n280_), .B1(new_n262_), .B2(new_n265_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G22gat), .B(G50gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(G78gat), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT29), .ZN(new_n289_));
  INV_X1    g088(.A(G141gat), .ZN(new_n290_));
  INV_X1    g089(.A(G148gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  AND2_X1   g091(.A1(KEYINPUT91), .A2(KEYINPUT3), .ZN(new_n293_));
  NOR2_X1   g092(.A1(KEYINPUT91), .A2(KEYINPUT3), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n292_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G141gat), .A2(G148gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(KEYINPUT2), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT2), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n298_), .A2(G141gat), .A3(G148gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(KEYINPUT91), .A2(KEYINPUT3), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n301_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n295_), .A2(new_n300_), .A3(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT92), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  OR2_X1    g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G155gat), .A2(G162gat), .ZN(new_n307_));
  AND2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n295_), .A2(new_n300_), .A3(KEYINPUT92), .A4(new_n302_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n305_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT1), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n306_), .A2(new_n311_), .A3(new_n307_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n313_));
  AND2_X1   g112(.A1(new_n313_), .A2(new_n296_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n312_), .A2(new_n314_), .A3(new_n292_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT90), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n312_), .A2(new_n314_), .A3(KEYINPUT90), .A4(new_n292_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n289_), .B1(new_n310_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G228gat), .A2(G233gat), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT21), .ZN(new_n323_));
  INV_X1    g122(.A(G204gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(G197gat), .ZN(new_n325_));
  INV_X1    g124(.A(G197gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(G204gat), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n323_), .B1(new_n325_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT95), .ZN(new_n329_));
  AND2_X1   g128(.A1(G211gat), .A2(G218gat), .ZN(new_n330_));
  NOR2_X1   g129(.A1(G211gat), .A2(G218gat), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n329_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  OR2_X1    g131(.A1(G211gat), .A2(G218gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G211gat), .A2(G218gat), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n333_), .A2(KEYINPUT95), .A3(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n328_), .A2(new_n332_), .A3(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT96), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n328_), .A2(new_n335_), .A3(new_n332_), .A4(KEYINPUT96), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n325_), .A2(new_n327_), .ZN(new_n341_));
  AOI22_X1  g140(.A1(new_n335_), .A2(new_n332_), .B1(new_n341_), .B2(KEYINPUT21), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n323_), .A2(KEYINPUT93), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT93), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT21), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G197gat), .B(G204gat), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n346_), .A2(new_n347_), .A3(KEYINPUT94), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(KEYINPUT94), .B1(new_n346_), .B2(new_n347_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n342_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  AND3_X1   g150(.A1(new_n340_), .A2(KEYINPUT97), .A3(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(KEYINPUT97), .B1(new_n340_), .B2(new_n351_), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n321_), .B(new_n322_), .C1(new_n352_), .C2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n350_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(new_n348_), .ZN(new_n356_));
  AOI22_X1  g155(.A1(new_n356_), .A2(new_n342_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n357_));
  OAI211_X1 g156(.A(G228gat), .B(G233gat), .C1(new_n320_), .C2(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n288_), .B1(new_n354_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n310_), .A2(new_n319_), .A3(new_n289_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT28), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT28), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n310_), .A2(new_n319_), .A3(new_n363_), .A4(new_n289_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(G106gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n354_), .A2(new_n358_), .A3(new_n288_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n360_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n365_), .B(G106gat), .ZN(new_n370_));
  INV_X1    g169(.A(new_n368_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n370_), .B1(new_n371_), .B2(new_n359_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n285_), .B1(new_n369_), .B2(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT89), .B1(new_n283_), .B2(new_n284_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n262_), .A2(new_n265_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n280_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT89), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n262_), .A2(new_n265_), .A3(new_n282_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n377_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n374_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n372_), .A2(new_n369_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n373_), .B1(new_n381_), .B2(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT18), .B(G64gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(G92gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G8gat), .B(G36gat), .ZN(new_n387_));
  XOR2_X1   g186(.A(new_n386_), .B(new_n387_), .Z(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n250_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G226gat), .A2(G233gat), .ZN(new_n391_));
  XOR2_X1   g190(.A(new_n391_), .B(KEYINPUT98), .Z(new_n392_));
  XOR2_X1   g191(.A(new_n392_), .B(KEYINPUT19), .Z(new_n393_));
  INV_X1    g192(.A(KEYINPUT20), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT101), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n221_), .A2(new_n213_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT100), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT22), .B(G169gat), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT100), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n398_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n224_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n240_), .A2(new_n207_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n404_), .A2(new_n211_), .A3(new_n405_), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n228_), .B(new_n235_), .C1(new_n231_), .C2(new_n232_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(new_n243_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(KEYINPUT99), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n206_), .A2(new_n209_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT99), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n407_), .A2(new_n412_), .A3(new_n243_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n409_), .A2(new_n411_), .A3(new_n245_), .A4(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n406_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n340_), .A2(new_n351_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n396_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n357_), .A2(KEYINPUT101), .A3(new_n414_), .A4(new_n406_), .ZN(new_n418_));
  AND4_X1   g217(.A1(new_n390_), .A2(new_n395_), .A3(new_n417_), .A4(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n393_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n357_), .A2(KEYINPUT97), .ZN(new_n421_));
  INV_X1    g220(.A(new_n250_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT97), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n416_), .A2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n421_), .A2(new_n422_), .A3(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n394_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n420_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n389_), .B1(new_n419_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT102), .ZN(new_n429_));
  NOR3_X1   g228(.A1(new_n352_), .A2(new_n353_), .A3(new_n250_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n412_), .B1(new_n407_), .B2(new_n243_), .ZN(new_n431_));
  NOR3_X1   g230(.A1(new_n431_), .A2(new_n410_), .A3(new_n244_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n211_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n433_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n434_));
  AOI22_X1  g233(.A1(new_n432_), .A2(new_n413_), .B1(new_n434_), .B2(new_n405_), .ZN(new_n435_));
  OAI21_X1  g234(.A(KEYINPUT20), .B1(new_n435_), .B2(new_n357_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n393_), .B1(new_n430_), .B2(new_n436_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n390_), .A2(new_n395_), .A3(new_n417_), .A4(new_n418_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n437_), .A2(new_n438_), .A3(new_n388_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n428_), .A2(new_n429_), .A3(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT27), .ZN(new_n441_));
  OAI211_X1 g240(.A(KEYINPUT102), .B(new_n389_), .C1(new_n419_), .C2(new_n427_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n440_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G225gat), .A2(G233gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n310_), .A2(new_n319_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT4), .ZN(new_n446_));
  AND4_X1   g245(.A1(KEYINPUT103), .A2(new_n445_), .A3(new_n446_), .A4(new_n275_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n278_), .B1(new_n310_), .B2(new_n319_), .ZN(new_n448_));
  AOI21_X1  g247(.A(KEYINPUT103), .B1(new_n448_), .B2(new_n446_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n445_), .A2(new_n275_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n310_), .A2(new_n319_), .A3(new_n278_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n451_), .A2(KEYINPUT4), .A3(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n444_), .B1(new_n450_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n444_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n455_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G1gat), .B(G29gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G57gat), .B(G85gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n457_), .B(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(KEYINPUT104), .B(KEYINPUT0), .ZN(new_n460_));
  XOR2_X1   g259(.A(new_n459_), .B(new_n460_), .Z(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NOR3_X1   g261(.A1(new_n454_), .A2(new_n456_), .A3(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n445_), .A2(new_n446_), .A3(new_n275_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT103), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n448_), .A2(KEYINPUT103), .A3(new_n446_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n453_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n456_), .B1(new_n468_), .B2(new_n455_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n469_), .A2(new_n461_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n463_), .A2(new_n470_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n420_), .B1(new_n430_), .B2(new_n436_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n394_), .B1(new_n435_), .B2(new_n357_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n390_), .A2(new_n473_), .A3(new_n393_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  OAI211_X1 g274(.A(new_n439_), .B(KEYINPUT27), .C1(new_n475_), .C2(new_n388_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n443_), .A2(new_n471_), .A3(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n450_), .A2(new_n444_), .A3(new_n453_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n451_), .A2(new_n455_), .A3(new_n452_), .ZN(new_n479_));
  AND3_X1   g278(.A1(new_n478_), .A2(new_n461_), .A3(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n480_), .B1(new_n440_), .B2(new_n442_), .ZN(new_n481_));
  OAI211_X1 g280(.A(KEYINPUT33), .B(new_n462_), .C1(new_n454_), .C2(new_n456_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT33), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n483_), .B1(new_n469_), .B2(new_n461_), .ZN(new_n484_));
  AND2_X1   g283(.A1(new_n482_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n388_), .A2(KEYINPUT32), .ZN(new_n486_));
  AND3_X1   g285(.A1(new_n437_), .A2(new_n438_), .A3(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n462_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n469_), .A2(new_n461_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n487_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  OR2_X1    g289(.A1(new_n475_), .A2(new_n486_), .ZN(new_n491_));
  AOI22_X1  g290(.A1(new_n481_), .A2(new_n485_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n382_), .A2(new_n374_), .A3(new_n380_), .ZN(new_n493_));
  OAI22_X1  g292(.A1(new_n384_), .A2(new_n477_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT13), .ZN(new_n495_));
  XOR2_X1   g294(.A(G57gat), .B(G64gat), .Z(new_n496_));
  INV_X1    g295(.A(KEYINPUT11), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G57gat), .B(G64gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT11), .ZN(new_n500_));
  XOR2_X1   g299(.A(G71gat), .B(G78gat), .Z(new_n501_));
  NAND3_X1  g300(.A1(new_n498_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  OR2_X1    g301(.A1(new_n500_), .A2(new_n501_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT12), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT66), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT7), .ZN(new_n508_));
  INV_X1    g307(.A(G99gat), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n508_), .A2(new_n509_), .A3(new_n366_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G99gat), .A2(G106gat), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT6), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n514_));
  OAI21_X1  g313(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n510_), .A2(new_n513_), .A3(new_n514_), .A4(new_n515_), .ZN(new_n516_));
  OR2_X1    g315(.A1(G85gat), .A2(G92gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G85gat), .A2(G92gat), .ZN(new_n518_));
  AND2_X1   g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  AND3_X1   g318(.A1(new_n516_), .A2(KEYINPUT8), .A3(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(KEYINPUT8), .B1(new_n516_), .B2(new_n519_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  XOR2_X1   g321(.A(KEYINPUT10), .B(G99gat), .Z(new_n523_));
  XOR2_X1   g322(.A(KEYINPUT64), .B(G106gat), .Z(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  OR2_X1    g324(.A1(new_n518_), .A2(KEYINPUT9), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n517_), .A2(KEYINPUT9), .A3(new_n518_), .ZN(new_n527_));
  AND2_X1   g326(.A1(new_n513_), .A2(new_n514_), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n525_), .A2(new_n526_), .A3(new_n527_), .A4(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n507_), .B1(new_n522_), .B2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n516_), .A2(new_n519_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT8), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n516_), .A2(KEYINPUT8), .A3(new_n519_), .ZN(new_n534_));
  AND4_X1   g333(.A1(new_n507_), .A2(new_n529_), .A3(new_n533_), .A4(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n506_), .B1(new_n530_), .B2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(KEYINPUT67), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n529_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT66), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n522_), .A2(new_n507_), .A3(new_n529_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT67), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n541_), .A2(new_n542_), .A3(new_n506_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n537_), .A2(new_n543_), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n502_), .A2(new_n503_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n538_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n538_), .A2(new_n545_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(new_n505_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT68), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT68), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n547_), .A2(new_n550_), .A3(new_n505_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n546_), .B1(new_n549_), .B2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G230gat), .A2(G233gat), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n544_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(KEYINPUT65), .B1(new_n538_), .B2(new_n545_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(new_n546_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n556_), .A2(G230gat), .A3(G233gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G120gat), .B(G148gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(new_n324_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT5), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(new_n241_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n554_), .A2(new_n557_), .A3(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(KEYINPUT69), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT69), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n554_), .A2(new_n564_), .A3(new_n557_), .A4(new_n561_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n561_), .B1(new_n554_), .B2(new_n557_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n495_), .B1(new_n566_), .B2(new_n568_), .ZN(new_n569_));
  AOI211_X1 g368(.A(KEYINPUT13), .B(new_n567_), .C1(new_n563_), .C2(new_n565_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  XOR2_X1   g370(.A(new_n571_), .B(KEYINPUT70), .Z(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT15), .ZN(new_n574_));
  XOR2_X1   g373(.A(G29gat), .B(G36gat), .Z(new_n575_));
  INV_X1    g374(.A(G43gat), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G29gat), .B(G36gat), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(G43gat), .ZN(new_n579_));
  AND3_X1   g378(.A1(new_n577_), .A2(G50gat), .A3(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(G50gat), .B1(new_n577_), .B2(new_n579_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n574_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n577_), .A2(new_n579_), .ZN(new_n583_));
  INV_X1    g382(.A(G50gat), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n577_), .A2(G50gat), .A3(new_n579_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n585_), .A2(KEYINPUT15), .A3(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n582_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(G1gat), .ZN(new_n590_));
  INV_X1    g389(.A(G8gat), .ZN(new_n591_));
  OAI21_X1  g390(.A(KEYINPUT14), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT76), .ZN(new_n593_));
  INV_X1    g392(.A(G15gat), .ZN(new_n594_));
  INV_X1    g393(.A(G22gat), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(G15gat), .A2(G22gat), .ZN(new_n597_));
  AOI22_X1  g396(.A1(new_n592_), .A2(new_n593_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n598_), .B1(new_n593_), .B2(new_n592_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G1gat), .B(G8gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT77), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n599_), .B(new_n601_), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n589_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G229gat), .A2(G233gat), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n580_), .A2(new_n581_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n602_), .A2(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n603_), .A2(new_n604_), .A3(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n602_), .B(new_n605_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n608_), .A2(G229gat), .A3(G233gat), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n607_), .A2(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G113gat), .B(G141gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(new_n217_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(new_n326_), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n610_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n610_), .A2(new_n613_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n602_), .B(new_n504_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(G231gat), .A2(G233gat), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n618_), .B(KEYINPUT78), .Z(new_n619_));
  OR2_X1    g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(KEYINPUT16), .B(G183gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(G211gat), .ZN(new_n622_));
  XOR2_X1   g421(.A(G127gat), .B(G155gat), .Z(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT17), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n617_), .A2(new_n619_), .ZN(new_n626_));
  AND3_X1   g425(.A1(new_n620_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT79), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n620_), .A2(new_n626_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT17), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n624_), .A2(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(KEYINPUT79), .B1(new_n630_), .B2(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n629_), .B1(new_n633_), .B2(new_n627_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n541_), .A2(new_n588_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(G232gat), .A2(G233gat), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT34), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(KEYINPUT35), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n637_), .A2(KEYINPUT35), .ZN(new_n639_));
  NOR3_X1   g438(.A1(new_n538_), .A2(new_n580_), .A3(new_n581_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n635_), .A2(new_n638_), .A3(new_n639_), .A4(new_n641_), .ZN(new_n642_));
  AOI22_X1  g441(.A1(new_n539_), .A2(new_n540_), .B1(new_n587_), .B2(new_n582_), .ZN(new_n643_));
  OAI211_X1 g442(.A(KEYINPUT35), .B(new_n637_), .C1(new_n643_), .C2(new_n640_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(KEYINPUT71), .B(G190gat), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(G218gat), .ZN(new_n646_));
  XOR2_X1   g445(.A(G134gat), .B(G162gat), .Z(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(G218gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n645_), .B(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n647_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n648_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT36), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n653_), .B(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(KEYINPUT74), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n653_), .A2(new_n654_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT74), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n648_), .A2(new_n652_), .A3(KEYINPUT36), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n657_), .A2(new_n658_), .A3(new_n659_), .ZN(new_n660_));
  AOI22_X1  g459(.A1(new_n642_), .A2(new_n644_), .B1(new_n656_), .B2(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(KEYINPUT37), .B1(new_n661_), .B2(KEYINPUT73), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n657_), .B(KEYINPUT72), .Z(new_n663_));
  AND3_X1   g462(.A1(new_n642_), .A2(new_n663_), .A3(new_n644_), .ZN(new_n664_));
  NOR3_X1   g463(.A1(new_n664_), .A2(new_n661_), .A3(KEYINPUT75), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT75), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n642_), .A2(new_n644_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n656_), .A2(new_n660_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n642_), .A2(new_n663_), .A3(new_n644_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n666_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n662_), .B1(new_n665_), .B2(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(KEYINPUT75), .B1(new_n664_), .B2(new_n661_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n669_), .A2(new_n666_), .A3(new_n670_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT73), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n669_), .A2(new_n675_), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n673_), .A2(new_n674_), .A3(KEYINPUT37), .A4(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n634_), .B1(new_n672_), .B2(new_n677_), .ZN(new_n678_));
  AND4_X1   g477(.A1(new_n494_), .A2(new_n573_), .A3(new_n616_), .A4(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n471_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n679_), .A2(new_n590_), .A3(new_n680_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT38), .ZN(new_n682_));
  INV_X1    g481(.A(new_n616_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n571_), .A2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(new_n494_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n664_), .A2(new_n661_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n634_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n685_), .A2(new_n471_), .A3(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n682_), .B1(new_n590_), .B2(new_n689_), .ZN(G1324gat));
  NOR2_X1   g489(.A1(new_n685_), .A2(new_n688_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n443_), .A2(new_n476_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n591_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT39), .Z(new_n694_));
  NAND3_X1  g493(.A1(new_n679_), .A2(new_n591_), .A3(new_n692_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  XOR2_X1   g495(.A(new_n696_), .B(KEYINPUT40), .Z(G1325gat));
  NAND2_X1  g496(.A1(new_n374_), .A2(new_n380_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n594_), .B1(new_n691_), .B2(new_n698_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT41), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n679_), .A2(new_n594_), .A3(new_n698_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(G1326gat));
  AOI21_X1  g501(.A(new_n595_), .B1(new_n691_), .B2(new_n383_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT105), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT42), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n383_), .A2(new_n595_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT106), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n679_), .A2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n705_), .A2(new_n708_), .ZN(G1327gat));
  NAND2_X1  g508(.A1(new_n634_), .A2(new_n686_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT110), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n685_), .A2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(G29gat), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n712_), .A2(new_n713_), .A3(new_n680_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n672_), .A2(new_n677_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT43), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n716_), .A2(KEYINPUT107), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n490_), .A2(new_n491_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n480_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n439_), .A2(new_n429_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n388_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n442_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n720_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n482_), .A2(new_n484_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n719_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n493_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n443_), .A2(new_n471_), .A3(new_n476_), .ZN(new_n730_));
  NOR3_X1   g529(.A1(new_n371_), .A2(new_n370_), .A3(new_n359_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n367_), .B1(new_n360_), .B2(new_n368_), .ZN(new_n732_));
  OAI22_X1  g531(.A1(new_n731_), .A2(new_n732_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n733_), .B1(new_n698_), .B2(new_n382_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n730_), .A2(new_n734_), .ZN(new_n735_));
  AOI211_X1 g534(.A(new_n715_), .B(new_n718_), .C1(new_n729_), .C2(new_n735_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n715_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n494_), .B2(new_n739_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n736_), .A2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n742_), .A2(KEYINPUT108), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT108), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n745_), .A2(KEYINPUT44), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  OAI211_X1 g546(.A(new_n634_), .B(new_n616_), .C1(new_n569_), .C2(new_n570_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n741_), .A2(new_n744_), .A3(new_n747_), .A4(new_n749_), .ZN(new_n750_));
  AOI22_X1  g549(.A1(new_n727_), .A2(new_n728_), .B1(new_n730_), .B2(new_n734_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n737_), .B1(new_n751_), .B2(new_n715_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n381_), .A2(new_n383_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n477_), .B1(new_n753_), .B2(new_n733_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n481_), .A2(new_n485_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n493_), .B1(new_n755_), .B2(new_n719_), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n739_), .B(new_n717_), .C1(new_n754_), .C2(new_n756_), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n752_), .A2(new_n747_), .A3(new_n757_), .A4(new_n749_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(new_n743_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n750_), .A2(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n713_), .B1(new_n760_), .B2(new_n680_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT109), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n761_), .A2(new_n762_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n714_), .B1(new_n763_), .B2(new_n764_), .ZN(G1328gat));
  INV_X1    g564(.A(G36gat), .ZN(new_n766_));
  XNOR2_X1  g565(.A(KEYINPUT111), .B(KEYINPUT112), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT45), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n712_), .A2(new_n766_), .A3(new_n692_), .A4(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n768_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n711_), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n771_), .A2(new_n684_), .A3(new_n766_), .A4(new_n494_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n692_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n770_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n769_), .A2(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n773_), .B1(new_n750_), .B2(new_n759_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n775_), .B1(new_n776_), .B2(new_n766_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT113), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n715_), .B1(new_n729_), .B2(new_n735_), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n757_), .B(new_n749_), .C1(new_n779_), .C2(new_n738_), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n780_), .A2(new_n745_), .A3(KEYINPUT44), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n758_), .A2(new_n743_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n692_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(G36gat), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT113), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n784_), .A2(new_n785_), .A3(new_n775_), .ZN(new_n786_));
  XOR2_X1   g585(.A(KEYINPUT114), .B(KEYINPUT46), .Z(new_n787_));
  NAND3_X1  g586(.A1(new_n778_), .A2(new_n786_), .A3(new_n787_), .ZN(new_n788_));
  OAI211_X1 g587(.A(KEYINPUT46), .B(new_n775_), .C1(new_n776_), .C2(new_n766_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT115), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT115), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n784_), .A2(new_n791_), .A3(KEYINPUT46), .A4(new_n775_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n788_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT116), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n788_), .A2(new_n793_), .A3(KEYINPUT116), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(G1329gat));
  INV_X1    g597(.A(new_n285_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n760_), .A2(new_n799_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n381_), .A2(G43gat), .ZN(new_n801_));
  AOI22_X1  g600(.A1(new_n800_), .A2(G43gat), .B1(new_n712_), .B2(new_n801_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(KEYINPUT117), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(KEYINPUT47), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT117), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n802_), .B(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT47), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n804_), .A2(new_n808_), .ZN(G1330gat));
  AOI21_X1  g608(.A(G50gat), .B1(new_n712_), .B2(new_n383_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n584_), .B1(new_n750_), .B2(new_n759_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n810_), .B1(new_n811_), .B2(new_n383_), .ZN(G1331gat));
  INV_X1    g611(.A(new_n571_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n813_), .A2(new_n616_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n814_), .A2(new_n494_), .A3(new_n678_), .ZN(new_n815_));
  XOR2_X1   g614(.A(new_n815_), .B(KEYINPUT118), .Z(new_n816_));
  AOI21_X1  g615(.A(G57gat), .B1(new_n816_), .B2(new_n680_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n572_), .A2(new_n494_), .A3(new_n683_), .ZN(new_n818_));
  NOR3_X1   g617(.A1(new_n818_), .A2(new_n471_), .A3(new_n688_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n817_), .B1(G57gat), .B2(new_n819_), .ZN(G1332gat));
  INV_X1    g619(.A(G64gat), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n818_), .A2(new_n688_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n821_), .B1(new_n822_), .B2(new_n692_), .ZN(new_n823_));
  XOR2_X1   g622(.A(new_n823_), .B(KEYINPUT48), .Z(new_n824_));
  NAND3_X1  g623(.A1(new_n816_), .A2(new_n821_), .A3(new_n692_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(G1333gat));
  INV_X1    g625(.A(G71gat), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n827_), .B1(new_n822_), .B2(new_n698_), .ZN(new_n828_));
  XOR2_X1   g627(.A(new_n828_), .B(KEYINPUT49), .Z(new_n829_));
  NAND3_X1  g628(.A1(new_n816_), .A2(new_n827_), .A3(new_n698_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(G1334gat));
  INV_X1    g630(.A(G78gat), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n832_), .B1(new_n822_), .B2(new_n383_), .ZN(new_n833_));
  XOR2_X1   g632(.A(new_n833_), .B(KEYINPUT50), .Z(new_n834_));
  NAND3_X1  g633(.A1(new_n816_), .A2(new_n832_), .A3(new_n383_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(G1335gat));
  NOR2_X1   g635(.A1(new_n818_), .A2(new_n711_), .ZN(new_n837_));
  AOI21_X1  g636(.A(G85gat), .B1(new_n837_), .B2(new_n680_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n741_), .A2(new_n634_), .A3(new_n814_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n839_), .A2(new_n471_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n838_), .B1(G85gat), .B2(new_n840_), .ZN(G1336gat));
  AOI21_X1  g640(.A(G92gat), .B1(new_n837_), .B2(new_n692_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n839_), .A2(new_n773_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n842_), .B1(G92gat), .B2(new_n843_), .ZN(G1337gat));
  NAND3_X1  g643(.A1(new_n837_), .A2(new_n523_), .A3(new_n799_), .ZN(new_n845_));
  OAI21_X1  g644(.A(G99gat), .B1(new_n839_), .B2(new_n381_), .ZN(new_n846_));
  XOR2_X1   g645(.A(KEYINPUT119), .B(KEYINPUT51), .Z(new_n847_));
  NAND3_X1  g646(.A1(new_n845_), .A2(new_n846_), .A3(new_n847_), .ZN(new_n848_));
  OR2_X1    g647(.A1(new_n848_), .A2(KEYINPUT120), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n845_), .A2(new_n846_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(KEYINPUT51), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n848_), .A2(KEYINPUT120), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n849_), .A2(new_n851_), .A3(new_n852_), .ZN(G1338gat));
  NAND3_X1  g652(.A1(new_n837_), .A2(new_n524_), .A3(new_n383_), .ZN(new_n854_));
  OAI21_X1  g653(.A(G106gat), .B1(new_n839_), .B2(new_n382_), .ZN(new_n855_));
  OR2_X1    g654(.A1(new_n855_), .A2(KEYINPUT52), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n855_), .A2(KEYINPUT52), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n854_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g659(.A1(new_n692_), .A2(new_n471_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT56), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n553_), .B1(new_n544_), .B2(new_n552_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT55), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n554_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n544_), .A2(new_n552_), .A3(KEYINPUT55), .A4(new_n553_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n561_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n864_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  AOI211_X1 g670(.A(KEYINPUT56), .B(new_n561_), .C1(new_n867_), .C2(new_n868_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n566_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n871_), .A2(new_n872_), .A3(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n566_), .A2(new_n568_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n608_), .A2(new_n604_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n603_), .A2(new_n606_), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n613_), .B(new_n876_), .C1(new_n877_), .C2(new_n604_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n614_), .A2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  AOI22_X1  g679(.A1(new_n874_), .A2(new_n616_), .B1(new_n875_), .B2(new_n880_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n863_), .B1(new_n881_), .B2(new_n686_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n875_), .A2(new_n880_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n871_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n872_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n884_), .A2(new_n885_), .A3(new_n566_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n883_), .B1(new_n886_), .B2(new_n683_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n686_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n887_), .A2(KEYINPUT57), .A3(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT58), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n890_), .B1(new_n886_), .B2(new_n879_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n874_), .A2(KEYINPUT58), .A3(new_n880_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n891_), .A2(new_n892_), .A3(new_n739_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n882_), .A2(new_n889_), .A3(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n634_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n569_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n570_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n616_), .B1(new_n896_), .B2(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT121), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT54), .ZN(new_n900_));
  NAND4_X1  g699(.A1(new_n898_), .A2(new_n899_), .A3(new_n900_), .A4(new_n678_), .ZN(new_n901_));
  OAI211_X1 g700(.A(new_n678_), .B(new_n683_), .C1(new_n569_), .C2(new_n570_), .ZN(new_n902_));
  OAI21_X1  g701(.A(KEYINPUT121), .B1(new_n902_), .B2(KEYINPUT54), .ZN(new_n903_));
  AND2_X1   g702(.A1(new_n901_), .A2(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT122), .ZN(new_n905_));
  AND3_X1   g704(.A1(new_n902_), .A2(new_n905_), .A3(KEYINPUT54), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n905_), .B1(new_n902_), .B2(KEYINPUT54), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n904_), .A2(new_n908_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n862_), .B1(new_n895_), .B2(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(new_n373_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  AOI21_X1  g711(.A(G113gat), .B1(new_n912_), .B2(new_n616_), .ZN(new_n913_));
  AOI21_X1  g712(.A(KEYINPUT59), .B1(new_n910_), .B2(new_n373_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n914_), .ZN(new_n915_));
  AOI22_X1  g714(.A1(new_n894_), .A2(new_n634_), .B1(new_n904_), .B2(new_n908_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT59), .ZN(new_n917_));
  NOR4_X1   g716(.A1(new_n916_), .A2(new_n917_), .A3(new_n733_), .A4(new_n862_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n683_), .B1(new_n915_), .B2(new_n919_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n913_), .B1(new_n920_), .B2(G113gat), .ZN(G1340gat));
  OAI21_X1  g720(.A(new_n572_), .B1(new_n914_), .B2(new_n918_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(KEYINPUT123), .ZN(new_n923_));
  INV_X1    g722(.A(KEYINPUT123), .ZN(new_n924_));
  OAI211_X1 g723(.A(new_n924_), .B(new_n572_), .C1(new_n914_), .C2(new_n918_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n923_), .A2(G120gat), .A3(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(G120gat), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n927_), .B1(new_n813_), .B2(KEYINPUT60), .ZN(new_n928_));
  OAI211_X1 g727(.A(new_n912_), .B(new_n928_), .C1(KEYINPUT60), .C2(new_n927_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n926_), .A2(new_n929_), .ZN(G1341gat));
  INV_X1    g729(.A(G127gat), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n931_), .B1(new_n911_), .B2(new_n634_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(KEYINPUT124), .ZN(new_n933_));
  AOI211_X1 g732(.A(new_n931_), .B(new_n634_), .C1(new_n915_), .C2(new_n919_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n933_), .A2(new_n934_), .ZN(G1342gat));
  AOI21_X1  g734(.A(G134gat), .B1(new_n912_), .B2(new_n686_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n715_), .B1(new_n915_), .B2(new_n919_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n936_), .B1(new_n937_), .B2(G134gat), .ZN(G1343gat));
  NOR3_X1   g737(.A1(new_n916_), .A2(new_n753_), .A3(new_n862_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n939_), .A2(new_n616_), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n940_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g740(.A1(new_n939_), .A2(new_n572_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n942_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g742(.A(new_n634_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n939_), .A2(new_n944_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(KEYINPUT61), .B(G155gat), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n945_), .B(new_n946_), .ZN(G1346gat));
  AOI21_X1  g746(.A(G162gat), .B1(new_n939_), .B2(new_n686_), .ZN(new_n948_));
  AND2_X1   g747(.A1(new_n739_), .A2(G162gat), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n948_), .B1(new_n939_), .B2(new_n949_), .ZN(G1347gat));
  NOR3_X1   g749(.A1(new_n916_), .A2(new_n680_), .A3(new_n773_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n381_), .A2(new_n383_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n951_), .A2(new_n952_), .ZN(new_n953_));
  OAI21_X1  g752(.A(G169gat), .B1(new_n953_), .B2(new_n683_), .ZN(new_n954_));
  INV_X1    g753(.A(KEYINPUT62), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n954_), .A2(new_n955_), .ZN(new_n956_));
  INV_X1    g755(.A(new_n953_), .ZN(new_n957_));
  NAND3_X1  g756(.A1(new_n957_), .A2(new_n402_), .A3(new_n616_), .ZN(new_n958_));
  OAI211_X1 g757(.A(KEYINPUT62), .B(G169gat), .C1(new_n953_), .C2(new_n683_), .ZN(new_n959_));
  NAND3_X1  g758(.A1(new_n956_), .A2(new_n958_), .A3(new_n959_), .ZN(G1348gat));
  AOI21_X1  g759(.A(new_n224_), .B1(new_n957_), .B2(new_n571_), .ZN(new_n961_));
  NAND3_X1  g760(.A1(new_n951_), .A2(G176gat), .A3(new_n952_), .ZN(new_n962_));
  OR3_X1    g761(.A1(new_n962_), .A2(KEYINPUT125), .A3(new_n573_), .ZN(new_n963_));
  OAI21_X1  g762(.A(KEYINPUT125), .B1(new_n962_), .B2(new_n573_), .ZN(new_n964_));
  AOI21_X1  g763(.A(new_n961_), .B1(new_n963_), .B2(new_n964_), .ZN(G1349gat));
  NOR2_X1   g764(.A1(new_n953_), .A2(new_n634_), .ZN(new_n966_));
  MUX2_X1   g765(.A(G183gat), .B(new_n233_), .S(new_n966_), .Z(G1350gat));
  NAND3_X1  g766(.A1(new_n957_), .A2(new_n686_), .A3(new_n236_), .ZN(new_n968_));
  NAND3_X1  g767(.A1(new_n951_), .A2(new_n739_), .A3(new_n952_), .ZN(new_n969_));
  INV_X1    g768(.A(KEYINPUT126), .ZN(new_n970_));
  AND3_X1   g769(.A1(new_n969_), .A2(new_n970_), .A3(G190gat), .ZN(new_n971_));
  AOI21_X1  g770(.A(new_n970_), .B1(new_n969_), .B2(G190gat), .ZN(new_n972_));
  OAI21_X1  g771(.A(new_n968_), .B1(new_n971_), .B2(new_n972_), .ZN(G1351gat));
  INV_X1    g772(.A(KEYINPUT127), .ZN(new_n974_));
  INV_X1    g773(.A(new_n753_), .ZN(new_n975_));
  NAND3_X1  g774(.A1(new_n951_), .A2(new_n974_), .A3(new_n975_), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n895_), .A2(new_n909_), .ZN(new_n977_));
  NOR2_X1   g776(.A1(new_n773_), .A2(new_n680_), .ZN(new_n978_));
  NAND3_X1  g777(.A1(new_n977_), .A2(new_n975_), .A3(new_n978_), .ZN(new_n979_));
  NAND2_X1  g778(.A1(new_n979_), .A2(KEYINPUT127), .ZN(new_n980_));
  AOI21_X1  g779(.A(new_n683_), .B1(new_n976_), .B2(new_n980_), .ZN(new_n981_));
  XNOR2_X1  g780(.A(new_n981_), .B(new_n326_), .ZN(G1352gat));
  AOI21_X1  g781(.A(new_n573_), .B1(new_n976_), .B2(new_n980_), .ZN(new_n983_));
  XNOR2_X1  g782(.A(new_n983_), .B(new_n324_), .ZN(G1353gat));
  AOI21_X1  g783(.A(new_n634_), .B1(new_n976_), .B2(new_n980_), .ZN(new_n985_));
  NOR2_X1   g784(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n986_));
  AND2_X1   g785(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n987_));
  OAI21_X1  g786(.A(new_n985_), .B1(new_n986_), .B2(new_n987_), .ZN(new_n988_));
  OAI21_X1  g787(.A(new_n988_), .B1(new_n985_), .B2(new_n986_), .ZN(G1354gat));
  NAND2_X1  g788(.A1(new_n976_), .A2(new_n980_), .ZN(new_n990_));
  AOI21_X1  g789(.A(G218gat), .B1(new_n990_), .B2(new_n686_), .ZN(new_n991_));
  AOI21_X1  g790(.A(new_n715_), .B1(new_n976_), .B2(new_n980_), .ZN(new_n992_));
  AOI21_X1  g791(.A(new_n991_), .B1(G218gat), .B2(new_n992_), .ZN(G1355gat));
endmodule


