//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 0 1 0 0 1 0 1 1 0 0 1 1 1 1 0 1 0 1 0 1 0 0 1 0 0 1 1 0 1 0 0 0 0 0 1 0 0 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n832_, new_n833_, new_n834_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n858_,
    new_n860_, new_n861_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n889_, new_n891_, new_n892_, new_n893_,
    new_n895_, new_n896_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_;
  XNOR2_X1  g000(.A(KEYINPUT25), .B(G183gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT26), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT80), .B(G190gat), .ZN(new_n204_));
  INV_X1    g003(.A(G190gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(KEYINPUT81), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT81), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT26), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n205_), .B1(new_n206_), .B2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT82), .ZN(new_n210_));
  AND2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n209_), .A2(new_n210_), .ZN(new_n212_));
  OAI221_X1 g011(.A(new_n202_), .B1(new_n203_), .B2(new_n204_), .C1(new_n211_), .C2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G169gat), .ZN(new_n214_));
  INV_X1    g013(.A(G176gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n216_), .A2(KEYINPUT24), .A3(new_n217_), .ZN(new_n218_));
  OR2_X1    g017(.A1(new_n216_), .A2(KEYINPUT24), .ZN(new_n219_));
  INV_X1    g018(.A(G183gat), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT23), .B1(new_n220_), .B2(new_n205_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n221_), .B(KEYINPUT83), .ZN(new_n222_));
  OR3_X1    g021(.A1(new_n220_), .A2(new_n205_), .A3(KEYINPUT23), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n213_), .A2(new_n218_), .A3(new_n219_), .A4(new_n224_), .ZN(new_n225_));
  NOR3_X1   g024(.A1(KEYINPUT84), .A2(KEYINPUT85), .A3(KEYINPUT22), .ZN(new_n226_));
  OAI21_X1  g025(.A(G169gat), .B1(new_n226_), .B2(G176gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n214_), .A2(KEYINPUT22), .ZN(new_n228_));
  AOI21_X1  g027(.A(G176gat), .B1(new_n228_), .B2(KEYINPUT84), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT22), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(G169gat), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n229_), .B(new_n231_), .C1(KEYINPUT84), .C2(new_n228_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT85), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n227_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT86), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n223_), .A2(new_n221_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n237_), .B1(G183gat), .B2(new_n204_), .ZN(new_n238_));
  OAI211_X1 g037(.A(KEYINPUT86), .B(new_n227_), .C1(new_n232_), .C2(new_n233_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n236_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n225_), .A2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G127gat), .B(G134gat), .ZN(new_n242_));
  INV_X1    g041(.A(G113gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(G120gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n241_), .B(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT30), .B(G71gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT87), .B(G99gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT31), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G15gat), .B(G43gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n252_), .B(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G227gat), .A2(G233gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n250_), .B(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(G141gat), .A2(G148gat), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G141gat), .A2(G148gat), .ZN(new_n261_));
  NOR2_X1   g060(.A1(G155gat), .A2(G162gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT88), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G155gat), .A2(G162gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT1), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n264_), .A2(KEYINPUT1), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT89), .ZN(new_n268_));
  OAI211_X1 g067(.A(new_n260_), .B(new_n261_), .C1(new_n266_), .C2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n259_), .B(KEYINPUT3), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT90), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT2), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n261_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n273_), .B1(KEYINPUT90), .B2(KEYINPUT2), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n261_), .A2(new_n271_), .A3(new_n272_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n270_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT91), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n270_), .A2(new_n274_), .A3(KEYINPUT91), .A4(new_n275_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n263_), .A2(new_n264_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT92), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n263_), .A2(KEYINPUT92), .A3(new_n264_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  AND3_X1   g084(.A1(new_n280_), .A2(KEYINPUT93), .A3(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(KEYINPUT93), .B1(new_n280_), .B2(new_n285_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n269_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  OAI21_X1  g087(.A(KEYINPUT28), .B1(new_n288_), .B2(KEYINPUT29), .ZN(new_n289_));
  INV_X1    g088(.A(new_n269_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n280_), .A2(new_n285_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT93), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n280_), .A2(KEYINPUT93), .A3(new_n285_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n290_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT28), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT29), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n295_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n289_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(G50gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G78gat), .B(G106gat), .ZN(new_n303_));
  INV_X1    g102(.A(G22gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n288_), .A2(KEYINPUT29), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G228gat), .A2(G233gat), .ZN(new_n308_));
  INV_X1    g107(.A(G197gat), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n309_), .A2(G204gat), .ZN(new_n310_));
  INV_X1    g109(.A(G204gat), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n311_), .A2(G197gat), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT21), .B1(new_n310_), .B2(new_n312_), .ZN(new_n313_));
  XOR2_X1   g112(.A(G211gat), .B(G218gat), .Z(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  OR3_X1    g114(.A1(new_n309_), .A2(KEYINPUT94), .A3(G204gat), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n312_), .A2(KEYINPUT94), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n316_), .B1(new_n317_), .B2(new_n310_), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n313_), .B(new_n315_), .C1(new_n318_), .C2(KEYINPUT21), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n318_), .A2(KEYINPUT21), .A3(new_n314_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n307_), .A2(new_n308_), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(KEYINPUT95), .ZN(new_n323_));
  AOI22_X1  g122(.A1(new_n288_), .A2(KEYINPUT29), .B1(G228gat), .B2(G233gat), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT95), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n324_), .A2(new_n325_), .A3(new_n321_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n323_), .A2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n321_), .B(KEYINPUT96), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n308_), .B1(new_n307_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n306_), .B1(new_n327_), .B2(new_n330_), .ZN(new_n331_));
  AOI211_X1 g130(.A(new_n329_), .B(new_n305_), .C1(new_n323_), .C2(new_n326_), .ZN(new_n332_));
  NOR3_X1   g131(.A1(new_n302_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n322_), .A2(KEYINPUT95), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n325_), .B1(new_n324_), .B2(new_n321_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n330_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(new_n305_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n327_), .A2(new_n330_), .A3(new_n306_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n301_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n258_), .B1(new_n333_), .B2(new_n339_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n302_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n337_), .A2(new_n301_), .A3(new_n338_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n341_), .A2(new_n342_), .A3(new_n257_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n340_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n321_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n225_), .A2(new_n240_), .A3(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n346_), .A2(KEYINPUT97), .A3(KEYINPUT20), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(KEYINPUT97), .B1(new_n346_), .B2(KEYINPUT20), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT103), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G226gat), .A2(G233gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT19), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n224_), .B1(G183gat), .B2(G190gat), .ZN(new_n355_));
  AND2_X1   g154(.A1(new_n231_), .A2(new_n228_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(new_n215_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n355_), .A2(new_n217_), .A3(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT98), .B(KEYINPUT24), .ZN(new_n359_));
  OR2_X1    g158(.A1(new_n359_), .A2(new_n216_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT26), .B(G190gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n202_), .A2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n359_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n360_), .A2(new_n237_), .A3(new_n362_), .A4(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n358_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(new_n321_), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n350_), .A2(new_n351_), .A3(new_n354_), .A4(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n346_), .A2(KEYINPUT20), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT97), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n370_), .A2(new_n354_), .A3(new_n366_), .A4(new_n347_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(KEYINPUT103), .ZN(new_n372_));
  OR2_X1    g171(.A1(new_n328_), .A2(new_n365_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n345_), .B1(new_n225_), .B2(new_n240_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(KEYINPUT102), .A2(KEYINPUT20), .ZN(new_n376_));
  OR2_X1    g175(.A1(KEYINPUT102), .A2(KEYINPUT20), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n373_), .A2(new_n375_), .A3(new_n376_), .A4(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(new_n353_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n367_), .A2(new_n372_), .A3(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G8gat), .B(G36gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G64gat), .B(G92gat), .ZN(new_n384_));
  XOR2_X1   g183(.A(new_n383_), .B(new_n384_), .Z(new_n385_));
  NAND2_X1  g184(.A1(new_n380_), .A2(new_n385_), .ZN(new_n386_));
  OAI211_X1 g185(.A(KEYINPUT20), .B(new_n354_), .C1(new_n365_), .C2(new_n321_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n387_), .A2(new_n374_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n370_), .A2(new_n366_), .A3(new_n347_), .ZN(new_n389_));
  AOI211_X1 g188(.A(new_n385_), .B(new_n388_), .C1(new_n389_), .C2(new_n353_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n386_), .A2(new_n391_), .A3(KEYINPUT27), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G1gat), .B(G29gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(G85gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(KEYINPUT0), .ZN(new_n395_));
  INV_X1    g194(.A(G57gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT100), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n295_), .A2(new_n399_), .A3(new_n246_), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n399_), .B(new_n269_), .C1(new_n286_), .C2(new_n287_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(new_n247_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n400_), .A2(new_n402_), .A3(KEYINPUT4), .ZN(new_n403_));
  OR3_X1    g202(.A1(new_n295_), .A2(KEYINPUT4), .A3(new_n246_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G225gat), .A2(G233gat), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n405_), .A2(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n407_), .B1(new_n400_), .B2(new_n402_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n398_), .B1(new_n408_), .B2(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n406_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n412_));
  NOR3_X1   g211(.A1(new_n412_), .A2(new_n409_), .A3(new_n397_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n411_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT27), .ZN(new_n415_));
  INV_X1    g214(.A(new_n385_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n389_), .A2(new_n353_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n388_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n416_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n415_), .B1(new_n419_), .B2(new_n390_), .ZN(new_n420_));
  AND3_X1   g219(.A1(new_n392_), .A2(new_n414_), .A3(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n397_), .B1(new_n412_), .B2(new_n409_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT33), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n400_), .A2(new_n402_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n398_), .B1(new_n425_), .B2(new_n406_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT101), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  OAI211_X1 g227(.A(KEYINPUT101), .B(new_n398_), .C1(new_n425_), .C2(new_n406_), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n428_), .B(new_n429_), .C1(new_n407_), .C2(new_n405_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n419_), .A2(new_n390_), .ZN(new_n431_));
  OAI211_X1 g230(.A(KEYINPUT33), .B(new_n397_), .C1(new_n412_), .C2(new_n409_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n424_), .A2(new_n430_), .A3(new_n431_), .A4(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n416_), .A2(KEYINPUT32), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n380_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n417_), .A2(new_n418_), .A3(new_n434_), .ZN(new_n437_));
  OAI211_X1 g236(.A(new_n436_), .B(new_n437_), .C1(new_n411_), .C2(new_n413_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n257_), .B1(new_n433_), .B2(new_n438_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n333_), .A2(new_n339_), .ZN(new_n440_));
  AOI22_X1  g239(.A1(new_n344_), .A2(new_n421_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(KEYINPUT10), .B(G99gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(KEYINPUT65), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT66), .ZN(new_n444_));
  INV_X1    g243(.A(G106gat), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n443_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n442_), .A2(KEYINPUT65), .ZN(new_n447_));
  INV_X1    g246(.A(G99gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT10), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT10), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(G99gat), .ZN(new_n451_));
  AND3_X1   g250(.A1(new_n449_), .A2(new_n451_), .A3(KEYINPUT65), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n445_), .B1(new_n447_), .B2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT66), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n446_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G85gat), .A2(G92gat), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(G85gat), .A2(G92gat), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  OR2_X1    g258(.A1(KEYINPUT67), .A2(KEYINPUT9), .ZN(new_n460_));
  NAND2_X1  g259(.A1(KEYINPUT67), .A2(KEYINPUT9), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n459_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G99gat), .A2(G106gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT6), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT6), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n465_), .A2(G99gat), .A3(G106gat), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT9), .ZN(new_n467_));
  AOI22_X1  g266(.A1(new_n464_), .A2(new_n466_), .B1(new_n457_), .B2(new_n467_), .ZN(new_n468_));
  AND3_X1   g267(.A1(new_n455_), .A2(new_n462_), .A3(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT8), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n448_), .A2(new_n445_), .A3(KEYINPUT7), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT7), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n472_), .B1(G99gat), .B2(G106gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n464_), .A2(new_n466_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n470_), .B1(new_n476_), .B2(new_n459_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT69), .ZN(new_n478_));
  AOI22_X1  g277(.A1(new_n473_), .A2(new_n471_), .B1(new_n464_), .B2(new_n466_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT68), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n470_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n474_), .A2(new_n475_), .A3(new_n480_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(new_n459_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n478_), .B1(new_n481_), .B2(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(KEYINPUT8), .B1(new_n476_), .B2(KEYINPUT68), .ZN(new_n485_));
  INV_X1    g284(.A(new_n459_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n486_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n485_), .A2(new_n487_), .A3(KEYINPUT69), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n477_), .B1(new_n484_), .B2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G57gat), .B(G64gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(KEYINPUT11), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G71gat), .B(G78gat), .ZN(new_n492_));
  XOR2_X1   g291(.A(new_n491_), .B(new_n492_), .Z(new_n493_));
  OAI21_X1  g292(.A(new_n493_), .B1(KEYINPUT11), .B2(new_n490_), .ZN(new_n494_));
  NOR3_X1   g293(.A1(new_n469_), .A2(new_n489_), .A3(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT12), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n496_), .A2(KEYINPUT72), .ZN(new_n497_));
  INV_X1    g296(.A(new_n477_), .ZN(new_n498_));
  NOR3_X1   g297(.A1(new_n481_), .A2(new_n483_), .A3(new_n478_), .ZN(new_n499_));
  AOI21_X1  g298(.A(KEYINPUT69), .B1(new_n485_), .B2(new_n487_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n498_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n455_), .A2(new_n462_), .A3(new_n468_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n497_), .B1(new_n503_), .B2(new_n494_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n496_), .A2(KEYINPUT72), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n495_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT71), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT70), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n501_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n489_), .A2(KEYINPUT70), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n469_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n494_), .A2(KEYINPUT12), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n507_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n489_), .A2(KEYINPUT70), .ZN(new_n514_));
  AOI211_X1 g313(.A(new_n508_), .B(new_n477_), .C1(new_n484_), .C2(new_n488_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n502_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n516_), .A2(KEYINPUT71), .A3(KEYINPUT12), .A4(new_n494_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G230gat), .A2(G233gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT64), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n506_), .A2(new_n513_), .A3(new_n517_), .A4(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n519_), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n503_), .A2(new_n494_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n521_), .B1(new_n522_), .B2(new_n495_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n520_), .A2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G120gat), .B(G148gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT5), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(G176gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(new_n311_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n529_), .A2(KEYINPUT73), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n524_), .A2(new_n530_), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n520_), .B(new_n523_), .C1(KEYINPUT73), .C2(new_n529_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT13), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n531_), .A2(KEYINPUT13), .A3(new_n532_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(KEYINPUT77), .B(G15gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(G22gat), .ZN(new_n539_));
  INV_X1    g338(.A(G1gat), .ZN(new_n540_));
  INV_X1    g339(.A(G8gat), .ZN(new_n541_));
  OAI21_X1  g340(.A(KEYINPUT14), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n539_), .A2(new_n542_), .ZN(new_n543_));
  XOR2_X1   g342(.A(G1gat), .B(G8gat), .Z(new_n544_));
  XOR2_X1   g343(.A(new_n543_), .B(new_n544_), .Z(new_n545_));
  XNOR2_X1  g344(.A(G29gat), .B(G36gat), .ZN(new_n546_));
  INV_X1    g345(.A(G43gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(new_n300_), .ZN(new_n549_));
  AND2_X1   g348(.A1(new_n549_), .A2(KEYINPUT15), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n549_), .A2(KEYINPUT15), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n545_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT78), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n549_), .B(KEYINPUT15), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT78), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n554_), .A2(new_n555_), .A3(new_n545_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G229gat), .A2(G233gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n548_), .B(G50gat), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n545_), .A2(new_n558_), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n553_), .A2(new_n556_), .A3(new_n557_), .A4(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n545_), .B(new_n558_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n557_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G113gat), .B(G141gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(new_n214_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(new_n309_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n560_), .A2(new_n563_), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT79), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n560_), .A2(new_n563_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(new_n566_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n570_), .B(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n537_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G231gat), .A2(G233gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n545_), .B(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(new_n494_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G127gat), .B(G155gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT16), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(new_n220_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(G211gat), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT17), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n583_), .A2(new_n584_), .ZN(new_n586_));
  OR3_X1    g385(.A1(new_n579_), .A2(new_n585_), .A3(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n579_), .A2(new_n585_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n501_), .A2(new_n502_), .A3(new_n549_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G232gat), .A2(G233gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT74), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT34), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT35), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n554_), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n590_), .B(new_n596_), .C1(new_n511_), .C2(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n594_), .A2(new_n595_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n516_), .A2(new_n554_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n599_), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n601_), .A2(new_n602_), .A3(new_n596_), .A4(new_n590_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT36), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G190gat), .B(G218gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(G134gat), .ZN(new_n606_));
  INV_X1    g405(.A(G162gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  AOI22_X1  g407(.A1(new_n600_), .A2(new_n603_), .B1(new_n604_), .B2(new_n608_), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n608_), .A2(new_n604_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(KEYINPUT75), .B(KEYINPUT36), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n600_), .A2(new_n612_), .A3(new_n603_), .A4(new_n608_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT37), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT76), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n615_), .B1(new_n613_), .B2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n614_), .A2(new_n617_), .ZN(new_n618_));
  OAI211_X1 g417(.A(new_n611_), .B(new_n613_), .C1(new_n616_), .C2(new_n615_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n589_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n441_), .A2(new_n576_), .A3(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n414_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n622_), .A2(new_n540_), .A3(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT38), .ZN(new_n625_));
  INV_X1    g424(.A(new_n614_), .ZN(new_n626_));
  NOR4_X1   g425(.A1(new_n441_), .A2(new_n576_), .A3(new_n589_), .A4(new_n626_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n627_), .A2(new_n623_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n625_), .B1(new_n540_), .B2(new_n628_), .ZN(G1324gat));
  INV_X1    g428(.A(KEYINPUT40), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n392_), .A2(new_n420_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n627_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(G8gat), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n634_), .A2(KEYINPUT39), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n634_), .A2(KEYINPUT39), .ZN(new_n636_));
  OR2_X1    g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT104), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n622_), .A2(new_n541_), .A3(new_n632_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n637_), .A2(new_n638_), .A3(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n638_), .B1(new_n637_), .B2(new_n639_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n630_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n642_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n644_), .A2(KEYINPUT40), .A3(new_n640_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n643_), .A2(new_n645_), .ZN(G1325gat));
  INV_X1    g445(.A(G15gat), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n647_), .B1(new_n627_), .B2(new_n257_), .ZN(new_n648_));
  XOR2_X1   g447(.A(KEYINPUT105), .B(KEYINPUT41), .Z(new_n649_));
  XNOR2_X1  g448(.A(new_n648_), .B(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n622_), .A2(new_n647_), .A3(new_n257_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(G1326gat));
  INV_X1    g451(.A(new_n440_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n304_), .B1(new_n627_), .B2(new_n653_), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT42), .Z(new_n655_));
  NAND3_X1  g454(.A1(new_n622_), .A2(new_n304_), .A3(new_n653_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(G1327gat));
  NOR2_X1   g456(.A1(new_n441_), .A2(new_n576_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n626_), .A2(new_n589_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT107), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(G29gat), .B1(new_n662_), .B2(new_n623_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n618_), .A2(new_n619_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT106), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n664_), .B(new_n665_), .ZN(new_n666_));
  OAI21_X1  g465(.A(KEYINPUT43), .B1(new_n666_), .B2(new_n441_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n343_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n257_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n421_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n439_), .A2(new_n440_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT43), .ZN(new_n673_));
  INV_X1    g472(.A(new_n664_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n672_), .A2(new_n673_), .A3(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n667_), .A2(new_n675_), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n676_), .A2(KEYINPUT44), .A3(new_n575_), .A4(new_n589_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n677_), .A2(G29gat), .A3(new_n623_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n664_), .B(KEYINPUT106), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n673_), .B1(new_n680_), .B2(new_n672_), .ZN(new_n681_));
  AOI211_X1 g480(.A(KEYINPUT43), .B(new_n664_), .C1(new_n670_), .C2(new_n671_), .ZN(new_n682_));
  OAI211_X1 g481(.A(new_n575_), .B(new_n589_), .C1(new_n681_), .C2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n663_), .B1(new_n679_), .B2(new_n685_), .ZN(G1328gat));
  INV_X1    g485(.A(G36gat), .ZN(new_n687_));
  INV_X1    g486(.A(new_n685_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n688_), .A2(new_n631_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n687_), .B1(new_n689_), .B2(new_n677_), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n661_), .A2(G36gat), .A3(new_n631_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT45), .ZN(new_n692_));
  OAI21_X1  g491(.A(KEYINPUT108), .B1(new_n690_), .B2(new_n692_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT46), .ZN(G1329gat));
  INV_X1    g493(.A(KEYINPUT47), .ZN(new_n695_));
  NAND4_X1  g494(.A1(new_n685_), .A2(new_n677_), .A3(G43gat), .A4(new_n257_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT110), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n547_), .B1(new_n661_), .B2(new_n258_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n696_), .A2(new_n697_), .A3(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n697_), .B1(new_n696_), .B2(new_n698_), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n700_), .A2(new_n701_), .A3(KEYINPUT109), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT109), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n696_), .A2(new_n698_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(KEYINPUT110), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n703_), .B1(new_n705_), .B2(new_n699_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n695_), .B1(new_n702_), .B2(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(KEYINPUT109), .B1(new_n700_), .B2(new_n701_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n705_), .A2(new_n703_), .A3(new_n699_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n708_), .A2(new_n709_), .A3(KEYINPUT47), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n707_), .A2(new_n710_), .ZN(G1330gat));
  AOI21_X1  g510(.A(G50gat), .B1(new_n662_), .B2(new_n653_), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n688_), .A2(new_n300_), .A3(new_n440_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n713_), .B2(new_n677_), .ZN(G1331gat));
  AND2_X1   g513(.A1(new_n535_), .A2(new_n536_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n715_), .A2(new_n573_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n672_), .A2(new_n716_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n717_), .A2(new_n621_), .ZN(new_n718_));
  AOI21_X1  g517(.A(G57gat), .B1(new_n718_), .B2(new_n623_), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT111), .Z(new_n720_));
  NOR3_X1   g519(.A1(new_n717_), .A2(new_n589_), .A3(new_n626_), .ZN(new_n721_));
  XOR2_X1   g520(.A(KEYINPUT112), .B(G57gat), .Z(new_n722_));
  NOR2_X1   g521(.A1(new_n414_), .A2(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n720_), .B1(new_n721_), .B2(new_n723_), .ZN(G1332gat));
  INV_X1    g523(.A(G64gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n725_), .B1(new_n721_), .B2(new_n632_), .ZN(new_n726_));
  XOR2_X1   g525(.A(KEYINPUT113), .B(KEYINPUT48), .Z(new_n727_));
  XNOR2_X1  g526(.A(new_n726_), .B(new_n727_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n718_), .A2(new_n725_), .A3(new_n632_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(G1333gat));
  INV_X1    g529(.A(G71gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n731_), .B1(new_n721_), .B2(new_n257_), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT49), .Z(new_n733_));
  NAND2_X1  g532(.A1(new_n257_), .A2(new_n731_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT114), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n718_), .A2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n733_), .A2(new_n736_), .ZN(G1334gat));
  INV_X1    g536(.A(G78gat), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n738_), .B1(new_n721_), .B2(new_n653_), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT50), .Z(new_n740_));
  NAND3_X1  g539(.A1(new_n718_), .A2(new_n738_), .A3(new_n653_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(G1335gat));
  AND3_X1   g541(.A1(new_n672_), .A2(new_n660_), .A3(new_n716_), .ZN(new_n743_));
  AOI21_X1  g542(.A(G85gat), .B1(new_n743_), .B2(new_n623_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n716_), .A2(new_n589_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT115), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n746_), .B1(new_n667_), .B2(new_n675_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n623_), .A2(G85gat), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n744_), .B1(new_n747_), .B2(new_n748_), .ZN(G1336gat));
  AOI21_X1  g548(.A(G92gat), .B1(new_n743_), .B2(new_n632_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n632_), .A2(G92gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(new_n747_), .B2(new_n751_), .ZN(G1337gat));
  AOI21_X1  g551(.A(new_n448_), .B1(new_n747_), .B2(new_n257_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n257_), .A2(new_n443_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n743_), .B2(new_n754_), .ZN(new_n755_));
  XOR2_X1   g554(.A(new_n755_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g555(.A1(new_n743_), .A2(new_n445_), .A3(new_n653_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n747_), .A2(new_n653_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(G106gat), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n759_), .A2(KEYINPUT52), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n759_), .A2(KEYINPUT52), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n757_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g562(.A1(new_n513_), .A2(new_n506_), .A3(new_n517_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(new_n521_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n765_), .A2(KEYINPUT55), .A3(new_n520_), .ZN(new_n766_));
  OR2_X1    g565(.A1(new_n520_), .A2(KEYINPUT55), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n766_), .A2(new_n528_), .A3(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(KEYINPUT56), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n520_), .A2(new_n523_), .A3(new_n529_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT56), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n766_), .A2(new_n767_), .A3(new_n771_), .A4(new_n528_), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n769_), .A2(new_n573_), .A3(new_n770_), .A4(new_n772_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n553_), .A2(new_n556_), .A3(new_n562_), .A4(new_n559_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n561_), .A2(new_n557_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n774_), .A2(new_n566_), .A3(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n568_), .ZN(new_n777_));
  XOR2_X1   g576(.A(new_n777_), .B(KEYINPUT117), .Z(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(new_n533_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n773_), .A2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(new_n614_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT57), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n781_), .A2(KEYINPUT118), .A3(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT118), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n626_), .B1(new_n773_), .B2(new_n779_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n784_), .B1(new_n785_), .B2(KEYINPUT57), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(KEYINPUT57), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n769_), .A2(new_n772_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n788_), .A2(KEYINPUT58), .A3(new_n778_), .A4(new_n770_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n778_), .A2(new_n769_), .A3(new_n770_), .A4(new_n772_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT58), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n789_), .A2(new_n674_), .A3(new_n792_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n783_), .A2(new_n786_), .A3(new_n787_), .A4(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(new_n589_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT116), .ZN(new_n796_));
  AND4_X1   g595(.A1(new_n796_), .A2(new_n620_), .A3(new_n715_), .A4(new_n574_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  AOI211_X1 g597(.A(new_n589_), .B(new_n573_), .C1(new_n618_), .C2(new_n619_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n715_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT116), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n798_), .A2(new_n801_), .A3(KEYINPUT54), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n796_), .B1(new_n799_), .B2(new_n715_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n803_), .B1(new_n804_), .B2(new_n797_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n802_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n795_), .A2(new_n806_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n632_), .A2(new_n414_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n809_), .A2(new_n343_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n807_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT119), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n807_), .A2(KEYINPUT119), .A3(new_n810_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(G113gat), .B1(new_n815_), .B2(new_n573_), .ZN(new_n816_));
  AND2_X1   g615(.A1(new_n793_), .A2(new_n787_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n817_), .B1(KEYINPUT57), .B2(new_n785_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n589_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n806_), .ZN(new_n820_));
  NOR3_X1   g619(.A1(new_n809_), .A2(KEYINPUT59), .A3(new_n343_), .ZN(new_n821_));
  AOI22_X1  g620(.A1(new_n820_), .A2(new_n821_), .B1(new_n811_), .B2(KEYINPUT59), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n574_), .A2(new_n243_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n816_), .B1(new_n822_), .B2(new_n823_), .ZN(G1340gat));
  AND2_X1   g623(.A1(new_n813_), .A2(new_n814_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT60), .B1(new_n537_), .B2(new_n245_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n822_), .A2(new_n537_), .ZN(new_n828_));
  OAI21_X1  g627(.A(G120gat), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  OR3_X1    g628(.A1(new_n825_), .A2(KEYINPUT60), .A3(new_n826_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(G1341gat));
  INV_X1    g630(.A(new_n589_), .ZN(new_n832_));
  AOI21_X1  g631(.A(G127gat), .B1(new_n815_), .B2(new_n832_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n832_), .A2(G127gat), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n833_), .B1(new_n822_), .B2(new_n834_), .ZN(G1342gat));
  INV_X1    g634(.A(G134gat), .ZN(new_n836_));
  OAI211_X1 g635(.A(KEYINPUT120), .B(new_n836_), .C1(new_n825_), .C2(new_n614_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT120), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n614_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n838_), .B1(new_n839_), .B2(G134gat), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n836_), .A2(KEYINPUT121), .ZN(new_n841_));
  OR2_X1    g640(.A1(new_n836_), .A2(KEYINPUT121), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n664_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  AOI22_X1  g642(.A1(new_n837_), .A2(new_n840_), .B1(new_n822_), .B2(new_n843_), .ZN(G1343gat));
  AOI21_X1  g643(.A(KEYINPUT118), .B1(new_n781_), .B2(new_n782_), .ZN(new_n845_));
  NOR3_X1   g644(.A1(new_n785_), .A2(new_n784_), .A3(KEYINPUT57), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n832_), .B1(new_n847_), .B2(new_n817_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n802_), .A2(new_n805_), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n669_), .B(new_n808_), .C1(new_n848_), .C2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT122), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n340_), .B1(new_n795_), .B2(new_n806_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n853_), .A2(KEYINPUT122), .A3(new_n808_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n852_), .A2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n573_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n537_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g658(.A1(new_n855_), .A2(new_n832_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(KEYINPUT61), .B(G155gat), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n860_), .B(new_n861_), .ZN(G1346gat));
  INV_X1    g661(.A(KEYINPUT123), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n614_), .A2(G162gat), .ZN(new_n864_));
  AOI21_X1  g663(.A(KEYINPUT122), .B1(new_n853_), .B2(new_n808_), .ZN(new_n865_));
  AOI22_X1  g664(.A1(new_n794_), .A2(new_n589_), .B1(new_n802_), .B2(new_n805_), .ZN(new_n866_));
  NOR4_X1   g665(.A1(new_n866_), .A2(new_n851_), .A3(new_n340_), .A4(new_n809_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n864_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n666_), .B1(new_n852_), .B2(new_n854_), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n863_), .B(new_n868_), .C1(new_n869_), .C2(new_n607_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n680_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(G162gat), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n863_), .B1(new_n873_), .B2(new_n868_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n871_), .A2(new_n874_), .ZN(G1347gat));
  XNOR2_X1  g674(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n631_), .A2(new_n623_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n879_), .A2(new_n343_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n820_), .A2(new_n880_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n881_), .A2(new_n574_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n877_), .B1(new_n882_), .B2(new_n214_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n356_), .ZN(new_n884_));
  OAI211_X1 g683(.A(G169gat), .B(new_n876_), .C1(new_n881_), .C2(new_n574_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n883_), .A2(new_n884_), .A3(new_n885_), .ZN(G1348gat));
  INV_X1    g685(.A(new_n881_), .ZN(new_n887_));
  AOI21_X1  g686(.A(G176gat), .B1(new_n887_), .B2(new_n537_), .ZN(new_n888_));
  NOR3_X1   g687(.A1(new_n866_), .A2(new_n215_), .A3(new_n715_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n888_), .B1(new_n880_), .B2(new_n889_), .ZN(G1349gat));
  NOR3_X1   g689(.A1(new_n881_), .A2(new_n202_), .A3(new_n589_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n807_), .A2(new_n832_), .A3(new_n880_), .ZN(new_n892_));
  XOR2_X1   g691(.A(new_n892_), .B(KEYINPUT125), .Z(new_n893_));
  AOI21_X1  g692(.A(new_n891_), .B1(new_n893_), .B2(new_n220_), .ZN(G1350gat));
  OAI21_X1  g693(.A(G190gat), .B1(new_n881_), .B2(new_n664_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n626_), .A2(new_n361_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n881_), .B2(new_n896_), .ZN(G1351gat));
  NOR3_X1   g696(.A1(new_n866_), .A2(new_n340_), .A3(new_n879_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(new_n573_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g699(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n901_));
  XNOR2_X1  g700(.A(KEYINPUT126), .B(G204gat), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n898_), .A2(new_n537_), .ZN(new_n903_));
  MUX2_X1   g702(.A(new_n901_), .B(new_n902_), .S(new_n903_), .Z(G1353gat));
  NAND2_X1  g703(.A1(new_n898_), .A2(new_n832_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n906_));
  AND2_X1   g705(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n905_), .A2(new_n906_), .A3(new_n907_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n908_), .B1(new_n906_), .B2(new_n905_), .ZN(G1354gat));
  NAND2_X1  g708(.A1(new_n898_), .A2(new_n626_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(KEYINPUT127), .B(G218gat), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n664_), .A2(new_n911_), .ZN(new_n912_));
  AOI22_X1  g711(.A1(new_n910_), .A2(new_n911_), .B1(new_n898_), .B2(new_n912_), .ZN(G1355gat));
endmodule


