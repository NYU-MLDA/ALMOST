//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 0 1 0 0 1 0 1 0 0 1 0 0 1 1 0 0 0 1 0 1 0 1 1 0 1 0 0 1 1 1 1 1 1 1 0 1 0 1 0 0 0 0 1 0 0 1 1 0 0 0 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n798_, new_n799_, new_n800_, new_n802_, new_n803_,
    new_n804_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n909_, new_n910_, new_n912_,
    new_n914_, new_n915_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n949_, new_n950_, new_n952_, new_n953_, new_n955_,
    new_n956_, new_n958_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n973_, new_n974_;
  NAND2_X1  g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT94), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT1), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT95), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n202_), .B(KEYINPUT94), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT95), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n208_), .A2(new_n209_), .A3(KEYINPUT1), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n206_), .A2(new_n207_), .A3(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT96), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n204_), .A2(new_n205_), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n206_), .A2(new_n210_), .A3(KEYINPUT96), .A4(new_n207_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n213_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  XOR2_X1   g015(.A(G141gat), .B(G148gat), .Z(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT106), .ZN(new_n219_));
  INV_X1    g018(.A(G141gat), .ZN(new_n220_));
  INV_X1    g019(.A(G148gat), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT98), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  OR2_X1    g021(.A1(new_n222_), .A2(KEYINPUT2), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n220_), .A2(new_n221_), .A3(KEYINPUT97), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT3), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n224_), .A2(KEYINPUT3), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n222_), .A2(KEYINPUT2), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n223_), .A2(new_n225_), .A3(new_n226_), .A4(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n228_), .A2(new_n208_), .A3(new_n207_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n218_), .A2(new_n219_), .A3(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G127gat), .B(G134gat), .ZN(new_n231_));
  INV_X1    g030(.A(G113gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n231_), .B(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(new_n233_), .B(G120gat), .Z(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n230_), .A2(KEYINPUT105), .A3(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT105), .ZN(new_n237_));
  INV_X1    g036(.A(new_n229_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n238_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n237_), .B1(new_n239_), .B2(new_n219_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n234_), .B1(new_n239_), .B2(new_n237_), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n236_), .B(KEYINPUT4), .C1(new_n240_), .C2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G225gat), .A2(G233gat), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  OR3_X1    g043(.A1(new_n239_), .A2(KEYINPUT4), .A3(new_n234_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n242_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  OAI211_X1 g045(.A(new_n236_), .B(new_n243_), .C1(new_n240_), .C2(new_n241_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT0), .B(G57gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(G85gat), .ZN(new_n249_));
  XOR2_X1   g048(.A(G1gat), .B(G29gat), .Z(new_n250_));
  XOR2_X1   g049(.A(new_n249_), .B(new_n250_), .Z(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n246_), .A2(new_n247_), .A3(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT107), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT33), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n242_), .A2(new_n243_), .A3(new_n245_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n236_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n256_), .B(new_n251_), .C1(new_n257_), .C2(new_n243_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT104), .ZN(new_n259_));
  OR2_X1    g058(.A1(G211gat), .A2(G218gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G211gat), .A2(G218gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT21), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G197gat), .B(G204gat), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT21), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n260_), .A2(new_n266_), .A3(new_n261_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n263_), .A2(new_n265_), .A3(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n262_), .A2(new_n264_), .A3(KEYINPUT21), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(G183gat), .ZN(new_n272_));
  INV_X1    g071(.A(G190gat), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT23), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT23), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n275_), .A2(G183gat), .A3(G190gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n274_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n272_), .A2(new_n273_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT89), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(G169gat), .ZN(new_n282_));
  INV_X1    g081(.A(G176gat), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  OR2_X1    g083(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n284_), .B1(new_n287_), .B2(new_n283_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n277_), .A2(KEYINPUT89), .A3(new_n278_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n281_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(G169gat), .A2(G176gat), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT87), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT24), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n294_), .B1(G169gat), .B2(G176gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n291_), .B(KEYINPUT87), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(new_n294_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT25), .B(G183gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT26), .B(G190gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n276_), .A2(KEYINPUT88), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT88), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n303_), .A2(new_n275_), .A3(G183gat), .A4(G190gat), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n302_), .A2(new_n274_), .A3(new_n304_), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n296_), .A2(new_n298_), .A3(new_n301_), .A4(new_n305_), .ZN(new_n306_));
  AND3_X1   g105(.A1(new_n290_), .A2(new_n306_), .A3(KEYINPUT90), .ZN(new_n307_));
  AOI21_X1  g106(.A(KEYINPUT90), .B1(new_n290_), .B2(new_n306_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n271_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G226gat), .A2(G233gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT19), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n309_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT103), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n287_), .A2(KEYINPUT102), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT102), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n316_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n283_), .B1(new_n315_), .B2(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n284_), .B1(new_n305_), .B2(new_n278_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n291_), .A2(new_n294_), .ZN(new_n320_));
  AND3_X1   g119(.A1(new_n301_), .A2(new_n277_), .A3(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(KEYINPUT101), .B1(new_n284_), .B2(new_n294_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT101), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n295_), .A2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n293_), .A2(new_n322_), .A3(new_n324_), .ZN(new_n325_));
  AOI22_X1  g124(.A1(new_n318_), .A2(new_n319_), .B1(new_n321_), .B2(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n314_), .B1(new_n326_), .B2(new_n270_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n319_), .A2(new_n318_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n321_), .A2(new_n325_), .ZN(new_n329_));
  AND4_X1   g128(.A1(new_n314_), .A2(new_n270_), .A3(new_n328_), .A4(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT20), .B1(new_n327_), .B2(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n259_), .B1(new_n313_), .B2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT20), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n270_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(KEYINPUT103), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n326_), .A2(new_n314_), .A3(new_n270_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n333_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n337_), .A2(KEYINPUT104), .A3(new_n312_), .A4(new_n309_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n332_), .A2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT18), .B(G64gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(G92gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G8gat), .B(G36gat), .ZN(new_n342_));
  XOR2_X1   g141(.A(new_n341_), .B(new_n342_), .Z(new_n343_));
  OR2_X1    g142(.A1(new_n326_), .A2(new_n270_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n290_), .A2(new_n306_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT90), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n290_), .A2(new_n306_), .A3(KEYINPUT90), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  OAI211_X1 g148(.A(KEYINPUT20), .B(new_n344_), .C1(new_n349_), .C2(new_n271_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(new_n311_), .ZN(new_n351_));
  AND3_X1   g150(.A1(new_n339_), .A2(new_n343_), .A3(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n343_), .B1(new_n339_), .B2(new_n351_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  AND2_X1   g153(.A1(new_n258_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT33), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n253_), .A2(KEYINPUT107), .A3(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n255_), .A2(new_n355_), .A3(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n246_), .A2(new_n247_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(new_n251_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(new_n253_), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n309_), .A2(new_n334_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n312_), .B1(new_n362_), .B2(KEYINPUT20), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n350_), .A2(new_n311_), .ZN(new_n364_));
  OAI211_X1 g163(.A(KEYINPUT32), .B(new_n343_), .C1(new_n363_), .C2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n343_), .A2(KEYINPUT32), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n339_), .A2(new_n366_), .A3(new_n351_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n361_), .A2(new_n365_), .A3(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n358_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G228gat), .A2(G233gat), .ZN(new_n370_));
  XOR2_X1   g169(.A(new_n370_), .B(KEYINPUT99), .Z(new_n371_));
  INV_X1    g170(.A(KEYINPUT29), .ZN(new_n372_));
  OAI211_X1 g171(.A(new_n271_), .B(new_n371_), .C1(new_n239_), .C2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n218_), .A2(new_n229_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n270_), .B1(new_n374_), .B2(KEYINPUT29), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n370_), .A2(KEYINPUT99), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n373_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  XOR2_X1   g176(.A(G78gat), .B(G106gat), .Z(new_n378_));
  AOI21_X1  g177(.A(KEYINPUT100), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n374_), .A2(KEYINPUT29), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G22gat), .B(G50gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT28), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n380_), .B(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n271_), .B1(new_n239_), .B2(new_n372_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n384_), .A2(KEYINPUT99), .A3(new_n370_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n378_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(new_n386_), .A3(new_n373_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n386_), .B1(new_n385_), .B2(new_n373_), .ZN(new_n389_));
  OAI22_X1  g188(.A1(new_n379_), .A2(new_n383_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n383_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n377_), .A2(new_n378_), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n391_), .A2(KEYINPUT100), .A3(new_n392_), .A4(new_n387_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n390_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G227gat), .A2(G233gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT91), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G71gat), .B(G99gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  XOR2_X1   g198(.A(G15gat), .B(G43gat), .Z(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT30), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n347_), .A2(new_n403_), .A3(new_n348_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n403_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT92), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n349_), .A2(KEYINPUT30), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT92), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n408_), .A2(new_n409_), .A3(new_n404_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n402_), .B1(new_n407_), .B2(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n409_), .B1(new_n408_), .B2(new_n404_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n412_), .A2(new_n401_), .ZN(new_n413_));
  OAI21_X1  g212(.A(KEYINPUT93), .B1(new_n411_), .B2(new_n413_), .ZN(new_n414_));
  NOR3_X1   g213(.A1(new_n405_), .A2(KEYINPUT92), .A3(new_n406_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n401_), .B1(new_n415_), .B2(new_n412_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT93), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n407_), .A2(new_n402_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n416_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n234_), .B(KEYINPUT31), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n414_), .A2(new_n419_), .A3(new_n421_), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n416_), .A2(new_n417_), .A3(new_n418_), .A4(new_n420_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n395_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n394_), .A2(new_n424_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n390_), .A2(new_n393_), .A3(new_n422_), .A4(new_n423_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n361_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n339_), .A2(new_n343_), .A3(new_n351_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n343_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n431_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n430_), .A2(new_n432_), .A3(KEYINPUT27), .ZN(new_n433_));
  OR2_X1    g232(.A1(new_n433_), .A2(KEYINPUT108), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT27), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n435_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n433_), .A2(KEYINPUT108), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n434_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  AOI22_X1  g238(.A1(new_n369_), .A2(new_n426_), .B1(new_n429_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT15), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G29gat), .B(G36gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G43gat), .B(G50gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n442_), .A2(new_n443_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(KEYINPUT75), .B(KEYINPUT76), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NOR3_X1   g247(.A1(new_n445_), .A2(new_n446_), .A3(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n442_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n443_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n447_), .B1(new_n452_), .B2(new_n444_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n441_), .B1(new_n449_), .B2(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n448_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n452_), .A2(new_n447_), .A3(new_n444_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(KEYINPUT15), .A3(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G1gat), .B(G8gat), .ZN(new_n458_));
  OR2_X1    g257(.A1(new_n458_), .A2(KEYINPUT81), .ZN(new_n459_));
  INV_X1    g258(.A(G15gat), .ZN(new_n460_));
  INV_X1    g259(.A(G22gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G15gat), .A2(G22gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G1gat), .A2(G8gat), .ZN(new_n464_));
  AOI22_X1  g263(.A1(new_n462_), .A2(new_n463_), .B1(KEYINPUT14), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n458_), .A2(KEYINPUT81), .ZN(new_n466_));
  AND3_X1   g265(.A1(new_n459_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n465_), .B1(new_n459_), .B2(new_n466_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n454_), .A2(new_n457_), .A3(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT86), .ZN(new_n471_));
  INV_X1    g270(.A(new_n469_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n455_), .A2(new_n456_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT85), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(KEYINPUT85), .B1(new_n455_), .B2(new_n456_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n472_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT86), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n454_), .A2(new_n469_), .A3(new_n478_), .A4(new_n457_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n471_), .A2(new_n477_), .A3(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G229gat), .A2(G233gat), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  OR2_X1    g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n477_), .ZN(new_n484_));
  NOR3_X1   g283(.A1(new_n475_), .A2(new_n472_), .A3(new_n476_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n482_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G113gat), .B(G141gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(new_n282_), .ZN(new_n488_));
  INV_X1    g287(.A(G197gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n488_), .B(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  AND3_X1   g290(.A1(new_n483_), .A2(new_n486_), .A3(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n491_), .B1(new_n483_), .B2(new_n486_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G99gat), .A2(G106gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(KEYINPUT6), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT6), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n497_), .A2(G99gat), .A3(G106gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(G85gat), .ZN(new_n500_));
  INV_X1    g299(.A(G92gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G85gat), .A2(G92gat), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n502_), .A2(KEYINPUT9), .A3(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n503_), .A2(KEYINPUT9), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n499_), .A2(new_n504_), .A3(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(KEYINPUT10), .B(G99gat), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n508_), .A2(G106gat), .ZN(new_n509_));
  OAI21_X1  g308(.A(KEYINPUT65), .B1(new_n507_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n503_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(G85gat), .A2(G92gat), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n505_), .B1(new_n513_), .B2(KEYINPUT9), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT65), .ZN(new_n515_));
  INV_X1    g314(.A(G106gat), .ZN(new_n516_));
  INV_X1    g315(.A(G99gat), .ZN(new_n517_));
  AND2_X1   g316(.A1(new_n517_), .A2(KEYINPUT10), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n517_), .A2(KEYINPUT10), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n516_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n514_), .A2(new_n515_), .A3(new_n499_), .A4(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n510_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT8), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT67), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n497_), .B1(G99gat), .B2(G106gat), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n495_), .A2(KEYINPUT6), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n524_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n517_), .A2(new_n516_), .A3(KEYINPUT66), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT7), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT7), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n530_), .A2(new_n517_), .A3(new_n516_), .A4(KEYINPUT66), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n496_), .A2(new_n498_), .A3(KEYINPUT67), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n527_), .A2(new_n529_), .A3(new_n531_), .A4(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n523_), .B1(new_n533_), .B2(new_n513_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n529_), .A2(new_n499_), .A3(new_n531_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n535_), .A2(new_n523_), .A3(new_n513_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n522_), .B1(new_n534_), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(G57gat), .ZN(new_n539_));
  INV_X1    g338(.A(G64gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT11), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G57gat), .A2(G64gat), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n541_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G71gat), .A2(G78gat), .ZN(new_n545_));
  INV_X1    g344(.A(G71gat), .ZN(new_n546_));
  INV_X1    g345(.A(G78gat), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n544_), .A2(new_n545_), .A3(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(KEYINPUT68), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n542_), .B1(new_n541_), .B2(new_n543_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT68), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n544_), .A2(new_n552_), .A3(new_n545_), .A4(new_n548_), .ZN(new_n553_));
  AND3_X1   g352(.A1(new_n550_), .A2(new_n551_), .A3(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n551_), .B1(new_n550_), .B2(new_n553_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n538_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT12), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT69), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n560_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n550_), .A2(new_n553_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n551_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n550_), .A2(new_n551_), .A3(new_n553_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n564_), .A2(KEYINPUT69), .A3(new_n565_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n561_), .A2(new_n566_), .A3(new_n538_), .A4(KEYINPUT12), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G230gat), .A2(G233gat), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n568_), .B(KEYINPUT64), .Z(new_n569_));
  NAND2_X1  g368(.A1(new_n564_), .A2(new_n565_), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n570_), .B(new_n522_), .C1(new_n534_), .C2(new_n537_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n559_), .A2(new_n567_), .A3(new_n569_), .A4(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n569_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n557_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n538_), .A2(new_n556_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n573_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  XOR2_X1   g375(.A(G120gat), .B(G148gat), .Z(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT72), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G176gat), .B(G204gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n572_), .A2(new_n576_), .A3(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT73), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n572_), .A2(new_n576_), .A3(KEYINPUT73), .A4(new_n582_), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT70), .ZN(new_n588_));
  AND3_X1   g387(.A1(new_n572_), .A2(new_n588_), .A3(new_n576_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n588_), .B1(new_n572_), .B2(new_n576_), .ZN(new_n590_));
  NOR3_X1   g389(.A1(new_n589_), .A2(new_n590_), .A3(new_n582_), .ZN(new_n591_));
  OAI21_X1  g390(.A(KEYINPUT74), .B1(new_n587_), .B2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n585_), .A2(new_n586_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n572_), .A2(new_n576_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(KEYINPUT70), .ZN(new_n595_));
  INV_X1    g394(.A(new_n582_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n572_), .A2(new_n588_), .A3(new_n576_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n595_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT74), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n593_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n592_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT13), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n592_), .A2(KEYINPUT13), .A3(new_n600_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NOR3_X1   g404(.A1(new_n440_), .A2(new_n494_), .A3(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT80), .ZN(new_n607_));
  INV_X1    g406(.A(new_n473_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(G232gat), .A2(G233gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT34), .ZN(new_n610_));
  OAI22_X1  g409(.A1(new_n538_), .A2(new_n608_), .B1(KEYINPUT35), .B2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n454_), .A2(new_n457_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT77), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n614_), .A2(new_n615_), .A3(new_n538_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n538_), .ZN(new_n617_));
  OAI21_X1  g416(.A(KEYINPUT77), .B1(new_n617_), .B2(new_n613_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n612_), .A2(new_n616_), .A3(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n610_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT35), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n611_), .B1(KEYINPUT78), .B2(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n623_), .A2(KEYINPUT78), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n625_), .B1(new_n614_), .B2(new_n538_), .ZN(new_n626_));
  AOI22_X1  g425(.A1(new_n619_), .A2(new_n622_), .B1(new_n624_), .B2(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G190gat), .B(G218gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(G134gat), .ZN(new_n629_));
  INV_X1    g428(.A(G162gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT36), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(new_n633_));
  OAI211_X1 g432(.A(new_n607_), .B(KEYINPUT37), .C1(new_n627_), .C2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT79), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n627_), .A2(new_n632_), .A3(new_n631_), .ZN(new_n636_));
  OR2_X1    g435(.A1(new_n627_), .A2(new_n633_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  OAI211_X1 g437(.A(new_n635_), .B(new_n636_), .C1(new_n638_), .C2(KEYINPUT79), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT37), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n637_), .A2(new_n636_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n640_), .B1(new_n641_), .B2(KEYINPUT80), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n639_), .A2(new_n642_), .ZN(new_n643_));
  AND2_X1   g442(.A1(G231gat), .A2(G233gat), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n469_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n469_), .A2(new_n644_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(new_n556_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n645_), .A2(new_n570_), .A3(new_n646_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(KEYINPUT16), .B(G183gat), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(G211gat), .ZN(new_n652_));
  XOR2_X1   g451(.A(G127gat), .B(G155gat), .Z(new_n653_));
  XNOR2_X1  g452(.A(new_n652_), .B(new_n653_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT17), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n650_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(KEYINPUT83), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT83), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n650_), .A2(new_n658_), .A3(new_n655_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n657_), .A2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n561_), .A2(new_n566_), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n661_), .A2(KEYINPUT82), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(KEYINPUT82), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n664_), .A2(new_n646_), .A3(new_n645_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT17), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n654_), .A2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n662_), .A2(new_n647_), .A3(new_n663_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n665_), .A2(new_n667_), .A3(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n660_), .A2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(KEYINPUT84), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT84), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n660_), .A2(new_n672_), .A3(new_n669_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n671_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n643_), .A2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n606_), .A2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n361_), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n677_), .A2(G1gat), .A3(new_n678_), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n679_), .B(KEYINPUT38), .Z(new_n680_));
  INV_X1    g479(.A(new_n670_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n606_), .A2(new_n641_), .A3(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(G1gat), .B1(new_n682_), .B2(new_n678_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n680_), .A2(new_n683_), .ZN(G1324gat));
  XNOR2_X1  g483(.A(KEYINPUT109), .B(KEYINPUT40), .ZN(new_n685_));
  OAI21_X1  g484(.A(G8gat), .B1(new_n682_), .B2(new_n439_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(KEYINPUT39), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT39), .ZN(new_n688_));
  OAI211_X1 g487(.A(new_n688_), .B(G8gat), .C1(new_n682_), .C2(new_n439_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n689_), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n677_), .A2(G8gat), .A3(new_n439_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n685_), .B1(new_n690_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n685_), .ZN(new_n694_));
  AOI211_X1 g493(.A(new_n694_), .B(new_n691_), .C1(new_n687_), .C2(new_n689_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n693_), .A2(new_n695_), .ZN(G1325gat));
  INV_X1    g495(.A(KEYINPUT41), .ZN(new_n697_));
  OAI21_X1  g496(.A(G15gat), .B1(new_n682_), .B2(new_n424_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT110), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n698_), .A2(KEYINPUT110), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n697_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n701_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n703_), .A2(KEYINPUT41), .A3(new_n699_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n677_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n424_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n705_), .A2(new_n460_), .A3(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n702_), .A2(new_n704_), .A3(new_n707_), .ZN(G1326gat));
  NAND3_X1  g507(.A1(new_n705_), .A2(new_n461_), .A3(new_n394_), .ZN(new_n709_));
  OAI21_X1  g508(.A(G22gat), .B1(new_n682_), .B2(new_n395_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n710_), .A2(KEYINPUT42), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n710_), .A2(KEYINPUT42), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n709_), .B1(new_n711_), .B2(new_n712_), .ZN(G1327gat));
  NOR3_X1   g512(.A1(new_n605_), .A2(new_n494_), .A3(new_n674_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n715_), .A2(new_n440_), .A3(new_n641_), .ZN(new_n716_));
  AOI21_X1  g515(.A(G29gat), .B1(new_n716_), .B2(new_n361_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n643_), .ZN(new_n718_));
  OAI21_X1  g517(.A(KEYINPUT43), .B1(new_n440_), .B2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT43), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n429_), .A2(new_n439_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n425_), .B1(new_n358_), .B2(new_n368_), .ZN(new_n722_));
  OAI211_X1 g521(.A(new_n720_), .B(new_n643_), .C1(new_n721_), .C2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n719_), .A2(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(KEYINPUT44), .B1(new_n724_), .B2(new_n714_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n726_));
  AOI211_X1 g525(.A(new_n726_), .B(new_n715_), .C1(new_n719_), .C2(new_n723_), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n725_), .A2(new_n727_), .A3(new_n678_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n717_), .B1(new_n728_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g528(.A(KEYINPUT46), .ZN(new_n730_));
  INV_X1    g529(.A(G36gat), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n725_), .A2(new_n727_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n731_), .B1(new_n732_), .B2(new_n438_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n716_), .A2(new_n731_), .A3(new_n438_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT45), .Z(new_n735_));
  OAI21_X1  g534(.A(new_n730_), .B1(new_n733_), .B2(new_n735_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n734_), .B(KEYINPUT45), .ZN(new_n737_));
  NOR3_X1   g536(.A1(new_n725_), .A2(new_n727_), .A3(new_n439_), .ZN(new_n738_));
  OAI211_X1 g537(.A(new_n737_), .B(KEYINPUT46), .C1(new_n738_), .C2(new_n731_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n736_), .A2(new_n739_), .ZN(G1329gat));
  INV_X1    g539(.A(new_n725_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n724_), .A2(KEYINPUT44), .A3(new_n714_), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n741_), .A2(G43gat), .A3(new_n706_), .A4(new_n742_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n716_), .A2(new_n706_), .ZN(new_n744_));
  OR2_X1    g543(.A1(new_n744_), .A2(G43gat), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(KEYINPUT47), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT47), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n743_), .A2(new_n748_), .A3(new_n745_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(G1330gat));
  AOI21_X1  g549(.A(G50gat), .B1(new_n716_), .B2(new_n394_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n394_), .A2(G50gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n732_), .B2(new_n752_), .ZN(G1331gat));
  INV_X1    g552(.A(new_n605_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n494_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n756_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n641_), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n757_), .A2(new_n758_), .A3(new_n675_), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n759_), .A2(G57gat), .A3(new_n361_), .ZN(new_n760_));
  NOR3_X1   g559(.A1(new_n757_), .A2(new_n643_), .A3(new_n675_), .ZN(new_n761_));
  AOI21_X1  g560(.A(G57gat), .B1(new_n761_), .B2(new_n361_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n760_), .A2(new_n762_), .ZN(G1332gat));
  NAND3_X1  g562(.A1(new_n761_), .A2(new_n540_), .A3(new_n438_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT111), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n759_), .A2(new_n438_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n765_), .B1(new_n766_), .B2(G64gat), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  AOI211_X1 g567(.A(KEYINPUT111), .B(new_n540_), .C1(new_n759_), .C2(new_n438_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(KEYINPUT48), .B1(new_n768_), .B2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT48), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n767_), .A2(new_n769_), .A3(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n764_), .B1(new_n771_), .B2(new_n773_), .ZN(G1333gat));
  NAND3_X1  g573(.A1(new_n761_), .A2(new_n546_), .A3(new_n706_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n759_), .ZN(new_n776_));
  OAI21_X1  g575(.A(G71gat), .B1(new_n776_), .B2(new_n424_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n777_), .A2(KEYINPUT49), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n777_), .A2(KEYINPUT49), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n775_), .B1(new_n778_), .B2(new_n779_), .ZN(G1334gat));
  NAND3_X1  g579(.A1(new_n761_), .A2(new_n547_), .A3(new_n394_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT50), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n759_), .A2(new_n394_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n782_), .B1(new_n783_), .B2(G78gat), .ZN(new_n784_));
  AOI211_X1 g583(.A(KEYINPUT50), .B(new_n547_), .C1(new_n759_), .C2(new_n394_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n781_), .B1(new_n784_), .B2(new_n785_), .ZN(G1335gat));
  INV_X1    g585(.A(new_n756_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n787_), .A2(new_n674_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n440_), .A2(new_n641_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n791_), .A2(new_n500_), .A3(new_n361_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n724_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n788_), .ZN(new_n794_));
  NOR3_X1   g593(.A1(new_n793_), .A2(new_n678_), .A3(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n792_), .B1(new_n795_), .B2(new_n500_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT112), .ZN(G1336gat));
  AOI21_X1  g596(.A(G92gat), .B1(new_n791_), .B2(new_n438_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n793_), .A2(new_n794_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n439_), .A2(new_n501_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n798_), .B1(new_n799_), .B2(new_n800_), .ZN(G1337gat));
  OR3_X1    g600(.A1(new_n790_), .A2(new_n508_), .A3(new_n424_), .ZN(new_n802_));
  NOR3_X1   g601(.A1(new_n793_), .A2(new_n424_), .A3(new_n794_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n802_), .B1(new_n803_), .B2(new_n517_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g604(.A1(new_n791_), .A2(new_n516_), .A3(new_n394_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n724_), .A2(new_n394_), .A3(new_n788_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n807_), .A2(new_n808_), .A3(G106gat), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n808_), .B1(new_n807_), .B2(G106gat), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n806_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(KEYINPUT53), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT53), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n813_), .B(new_n806_), .C1(new_n809_), .C2(new_n810_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(new_n814_), .ZN(G1339gat));
  INV_X1    g614(.A(new_n428_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n438_), .A2(new_n678_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT115), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n818_), .A2(KEYINPUT57), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT114), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n480_), .A2(new_n821_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n471_), .A2(new_n477_), .A3(KEYINPUT114), .A4(new_n479_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n822_), .A2(new_n482_), .A3(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n481_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n824_), .A2(new_n490_), .A3(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n483_), .A2(new_n486_), .A3(new_n491_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n559_), .A2(new_n571_), .A3(new_n567_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n573_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n831_), .A2(KEYINPUT55), .A3(new_n572_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n575_), .B1(new_n558_), .B2(new_n557_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT55), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n833_), .A2(new_n834_), .A3(new_n569_), .A4(new_n567_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n832_), .A2(new_n596_), .A3(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT56), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n832_), .A2(KEYINPUT56), .A3(new_n596_), .A4(new_n835_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n494_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n601_), .A2(new_n829_), .B1(new_n840_), .B2(new_n593_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n820_), .B1(new_n841_), .B2(new_n758_), .ZN(new_n842_));
  AND3_X1   g641(.A1(new_n593_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n599_), .B1(new_n593_), .B2(new_n598_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n829_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n838_), .A2(new_n839_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n846_), .A2(new_n755_), .A3(new_n593_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n758_), .B1(new_n845_), .B2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n819_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n842_), .A2(new_n849_), .ZN(new_n850_));
  AOI211_X1 g649(.A(new_n587_), .B(new_n828_), .C1(new_n838_), .C2(new_n839_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT116), .ZN(new_n852_));
  OAI21_X1  g651(.A(KEYINPUT58), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n846_), .A2(new_n593_), .A3(new_n829_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT58), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n854_), .A2(KEYINPUT116), .A3(new_n855_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n853_), .A2(new_n643_), .A3(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n681_), .B1(new_n850_), .B2(new_n857_), .ZN(new_n858_));
  AND4_X1   g657(.A1(new_n494_), .A2(new_n639_), .A3(new_n674_), .A4(new_n642_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT54), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n860_), .A2(KEYINPUT113), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n859_), .A2(new_n604_), .A3(new_n603_), .A4(new_n861_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n639_), .A2(new_n674_), .A3(new_n642_), .A4(new_n494_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n605_), .B2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n862_), .A2(new_n865_), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n816_), .B(new_n817_), .C1(new_n858_), .C2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(KEYINPUT59), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n848_), .A2(new_n819_), .ZN(new_n869_));
  AOI211_X1 g668(.A(new_n758_), .B(new_n820_), .C1(new_n845_), .C2(new_n847_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n857_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n675_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n866_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT59), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n874_), .A2(new_n875_), .A3(new_n816_), .A4(new_n817_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n868_), .A2(new_n876_), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n877_), .A2(new_n232_), .A3(new_n494_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n867_), .A2(KEYINPUT117), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n871_), .A2(new_n670_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n873_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT117), .ZN(new_n882_));
  NAND4_X1  g681(.A1(new_n881_), .A2(new_n882_), .A3(new_n816_), .A4(new_n817_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n879_), .A2(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(G113gat), .B1(new_n884_), .B2(new_n755_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n878_), .A2(new_n885_), .ZN(G1340gat));
  XOR2_X1   g685(.A(KEYINPUT118), .B(G120gat), .Z(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n888_), .B1(new_n754_), .B2(KEYINPUT60), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n884_), .B(new_n889_), .C1(KEYINPUT60), .C2(new_n888_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n887_), .B1(new_n877_), .B2(new_n754_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(G1341gat));
  AOI21_X1  g691(.A(G127gat), .B1(new_n884_), .B2(new_n674_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n877_), .ZN(new_n894_));
  XOR2_X1   g693(.A(KEYINPUT119), .B(G127gat), .Z(new_n895_));
  NAND2_X1  g694(.A1(new_n681_), .A2(new_n895_), .ZN(new_n896_));
  XOR2_X1   g695(.A(new_n896_), .B(KEYINPUT120), .Z(new_n897_));
  AOI21_X1  g696(.A(new_n893_), .B1(new_n894_), .B2(new_n897_), .ZN(G1342gat));
  XNOR2_X1  g697(.A(KEYINPUT121), .B(G134gat), .ZN(new_n899_));
  NAND4_X1  g698(.A1(new_n868_), .A2(new_n876_), .A3(new_n643_), .A4(new_n899_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n641_), .B1(new_n879_), .B2(new_n883_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(G134gat), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT122), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  OAI211_X1 g703(.A(KEYINPUT122), .B(new_n900_), .C1(new_n901_), .C2(G134gat), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(G1343gat));
  AOI21_X1  g705(.A(new_n866_), .B1(new_n670_), .B2(new_n871_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n907_), .A2(new_n427_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(new_n817_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n909_), .A2(new_n494_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(new_n220_), .ZN(G1344gat));
  NOR2_X1   g710(.A1(new_n909_), .A2(new_n754_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(new_n221_), .ZN(G1345gat));
  NOR2_X1   g712(.A1(new_n909_), .A2(new_n675_), .ZN(new_n914_));
  XOR2_X1   g713(.A(KEYINPUT61), .B(G155gat), .Z(new_n915_));
  XNOR2_X1  g714(.A(new_n914_), .B(new_n915_), .ZN(G1346gat));
  NOR3_X1   g715(.A1(new_n909_), .A2(new_n630_), .A3(new_n718_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n630_), .B1(new_n909_), .B2(new_n641_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(KEYINPUT123), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT123), .ZN(new_n920_));
  OAI211_X1 g719(.A(new_n920_), .B(new_n630_), .C1(new_n909_), .C2(new_n641_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n917_), .B1(new_n919_), .B2(new_n921_), .ZN(G1347gat));
  INV_X1    g721(.A(KEYINPUT62), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n428_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n439_), .A2(new_n361_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n924_), .A2(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(new_n755_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n923_), .B1(new_n928_), .B2(G169gat), .ZN(new_n929_));
  AOI211_X1 g728(.A(KEYINPUT62), .B(new_n282_), .C1(new_n927_), .C2(new_n755_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n755_), .B1(new_n317_), .B2(new_n315_), .ZN(new_n931_));
  XOR2_X1   g730(.A(new_n931_), .B(KEYINPUT124), .Z(new_n932_));
  OAI22_X1  g731(.A1(new_n929_), .A2(new_n930_), .B1(new_n926_), .B2(new_n932_), .ZN(G1348gat));
  AOI21_X1  g732(.A(G176gat), .B1(new_n927_), .B2(new_n605_), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT125), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n935_), .B1(new_n907_), .B2(new_n394_), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n881_), .A2(KEYINPUT125), .A3(new_n395_), .ZN(new_n937_));
  AND4_X1   g736(.A1(new_n706_), .A2(new_n936_), .A3(new_n937_), .A4(new_n925_), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT126), .ZN(new_n939_));
  NAND4_X1  g738(.A1(new_n938_), .A2(new_n939_), .A3(G176gat), .A4(new_n605_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n881_), .A2(new_n395_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n424_), .B1(new_n941_), .B2(new_n935_), .ZN(new_n942_));
  INV_X1    g741(.A(new_n925_), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n394_), .B1(new_n880_), .B2(new_n873_), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n943_), .B1(new_n944_), .B2(KEYINPUT125), .ZN(new_n945_));
  NAND4_X1  g744(.A1(new_n942_), .A2(G176gat), .A3(new_n605_), .A4(new_n945_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n946_), .A2(KEYINPUT126), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n934_), .B1(new_n940_), .B2(new_n947_), .ZN(G1349gat));
  NOR3_X1   g747(.A1(new_n926_), .A2(new_n299_), .A3(new_n670_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n938_), .A2(new_n674_), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n949_), .B1(new_n950_), .B2(new_n272_), .ZN(G1350gat));
  OAI21_X1  g750(.A(G190gat), .B1(new_n926_), .B2(new_n718_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n758_), .A2(new_n300_), .ZN(new_n953_));
  OAI21_X1  g752(.A(new_n952_), .B1(new_n926_), .B2(new_n953_), .ZN(G1351gat));
  NOR3_X1   g753(.A1(new_n907_), .A2(new_n427_), .A3(new_n943_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n955_), .A2(new_n755_), .ZN(new_n956_));
  XNOR2_X1  g755(.A(new_n956_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g756(.A1(new_n955_), .A2(new_n605_), .ZN(new_n958_));
  XNOR2_X1  g757(.A(new_n958_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g758(.A1(new_n908_), .A2(new_n925_), .ZN(new_n960_));
  NOR2_X1   g759(.A1(new_n960_), .A2(new_n670_), .ZN(new_n961_));
  INV_X1    g760(.A(KEYINPUT127), .ZN(new_n962_));
  INV_X1    g761(.A(KEYINPUT63), .ZN(new_n963_));
  INV_X1    g762(.A(G211gat), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n963_), .A2(new_n964_), .ZN(new_n965_));
  NOR2_X1   g764(.A1(new_n963_), .A2(new_n964_), .ZN(new_n966_));
  INV_X1    g765(.A(new_n966_), .ZN(new_n967_));
  NAND4_X1  g766(.A1(new_n961_), .A2(new_n962_), .A3(new_n965_), .A4(new_n967_), .ZN(new_n968_));
  OAI211_X1 g767(.A(new_n963_), .B(new_n964_), .C1(new_n960_), .C2(new_n670_), .ZN(new_n969_));
  NAND3_X1  g768(.A1(new_n955_), .A2(new_n681_), .A3(new_n965_), .ZN(new_n970_));
  OAI21_X1  g769(.A(KEYINPUT127), .B1(new_n970_), .B2(new_n966_), .ZN(new_n971_));
  AND3_X1   g770(.A1(new_n968_), .A2(new_n969_), .A3(new_n971_), .ZN(G1354gat));
  AOI21_X1  g771(.A(G218gat), .B1(new_n955_), .B2(new_n758_), .ZN(new_n973_));
  NOR2_X1   g772(.A1(new_n960_), .A2(new_n718_), .ZN(new_n974_));
  AOI21_X1  g773(.A(new_n973_), .B1(new_n974_), .B2(G218gat), .ZN(G1355gat));
endmodule


