//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 1 1 0 1 0 1 0 0 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1 0 1 1 0 0 1 0 1 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n898_, new_n900_,
    new_n901_, new_n903_, new_n904_, new_n905_, new_n907_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_, new_n921_, new_n922_, new_n923_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n948_, new_n949_;
  INV_X1    g000(.A(KEYINPUT82), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G183gat), .A2(G190gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n203_), .A2(KEYINPUT23), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT23), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT81), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT81), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT23), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n204_), .B1(new_n209_), .B2(new_n203_), .ZN(new_n210_));
  OR2_X1    g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n211_), .A2(KEYINPUT24), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n202_), .B1(new_n210_), .B2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n212_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT81), .B(KEYINPUT23), .ZN(new_n215_));
  INV_X1    g014(.A(new_n203_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  OAI211_X1 g016(.A(KEYINPUT82), .B(new_n214_), .C1(new_n217_), .C2(new_n204_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219_));
  AND3_X1   g018(.A1(new_n211_), .A2(KEYINPUT24), .A3(new_n219_), .ZN(new_n220_));
  AND2_X1   g019(.A1(KEYINPUT80), .A2(G183gat), .ZN(new_n221_));
  NOR2_X1   g020(.A1(KEYINPUT80), .A2(G183gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT25), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n223_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(G190gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT26), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT26), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(G190gat), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n220_), .B1(new_n226_), .B2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n213_), .A2(new_n218_), .A3(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n219_), .ZN(new_n234_));
  XOR2_X1   g033(.A(KEYINPUT83), .B(G176gat), .Z(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  XOR2_X1   g035(.A(KEYINPUT22), .B(G169gat), .Z(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n234_), .B1(new_n236_), .B2(new_n238_), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n221_), .A2(new_n222_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n240_), .A2(G190gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n203_), .A2(new_n205_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n242_), .B1(new_n215_), .B2(new_n203_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n239_), .B1(new_n241_), .B2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n233_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G71gat), .B(G99gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(G43gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n245_), .B(new_n247_), .ZN(new_n248_));
  XOR2_X1   g047(.A(G127gat), .B(G134gat), .Z(new_n249_));
  XOR2_X1   g048(.A(G113gat), .B(G120gat), .Z(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n248_), .B(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G227gat), .A2(G233gat), .ZN(new_n254_));
  INV_X1    g053(.A(G15gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT30), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT31), .ZN(new_n258_));
  XOR2_X1   g057(.A(new_n253_), .B(new_n258_), .Z(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G141gat), .A2(G148gat), .ZN(new_n261_));
  INV_X1    g060(.A(G141gat), .ZN(new_n262_));
  INV_X1    g061(.A(G148gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G155gat), .A2(G162gat), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT84), .B1(new_n265_), .B2(KEYINPUT1), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(KEYINPUT1), .ZN(new_n267_));
  NOR2_X1   g066(.A1(G155gat), .A2(G162gat), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n266_), .A2(new_n267_), .A3(new_n269_), .ZN(new_n270_));
  NOR3_X1   g069(.A1(new_n265_), .A2(KEYINPUT84), .A3(KEYINPUT1), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n261_), .B(new_n264_), .C1(new_n270_), .C2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT2), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n261_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT85), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT85), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n276_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT86), .ZN(new_n280_));
  AND3_X1   g079(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n262_), .A2(new_n263_), .A3(KEYINPUT3), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT3), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n283_), .B1(G141gat), .B2(G148gat), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n281_), .B1(new_n282_), .B2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n279_), .A2(new_n280_), .A3(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT87), .ZN(new_n287_));
  AND3_X1   g086(.A1(new_n269_), .A2(new_n287_), .A3(new_n265_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n287_), .B1(new_n269_), .B2(new_n265_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n286_), .A2(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n280_), .B1(new_n279_), .B2(new_n285_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n272_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(new_n252_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n277_), .B(new_n275_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n281_), .ZN(new_n296_));
  NOR3_X1   g095(.A1(new_n283_), .A2(G141gat), .A3(G148gat), .ZN(new_n297_));
  AOI21_X1  g096(.A(KEYINPUT3), .B1(new_n262_), .B2(new_n263_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n296_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  OAI21_X1  g098(.A(KEYINPUT86), .B1(new_n295_), .B2(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n300_), .A2(new_n286_), .A3(new_n290_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n301_), .A2(new_n272_), .A3(new_n251_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n294_), .A2(KEYINPUT4), .A3(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G225gat), .A2(G233gat), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n251_), .B1(new_n301_), .B2(new_n272_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT94), .B(KEYINPUT4), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n304_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n303_), .A2(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n294_), .A2(new_n302_), .A3(new_n304_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G1gat), .B(G29gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(G85gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT0), .B(G57gat), .ZN(new_n313_));
  XOR2_X1   g112(.A(new_n312_), .B(new_n313_), .Z(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n310_), .A2(new_n315_), .ZN(new_n316_));
  AND3_X1   g115(.A1(new_n294_), .A2(KEYINPUT4), .A3(new_n302_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n293_), .A2(new_n252_), .A3(new_n306_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n304_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  OAI211_X1 g119(.A(new_n309_), .B(new_n314_), .C1(new_n317_), .C2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n316_), .A2(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n260_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT29), .ZN(new_n324_));
  OAI211_X1 g123(.A(new_n324_), .B(new_n272_), .C1(new_n291_), .C2(new_n292_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(KEYINPUT28), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT28), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n301_), .A2(new_n327_), .A3(new_n324_), .A4(new_n272_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G22gat), .B(G50gat), .ZN(new_n329_));
  AND3_X1   g128(.A1(new_n326_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n329_), .B1(new_n326_), .B2(new_n328_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT90), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G228gat), .A2(G233gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT88), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n324_), .B1(new_n301_), .B2(new_n272_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT89), .ZN(new_n338_));
  INV_X1    g137(.A(G204gat), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n338_), .B1(new_n339_), .B2(G197gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(G197gat), .ZN(new_n341_));
  INV_X1    g140(.A(G197gat), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n342_), .A2(KEYINPUT89), .A3(G204gat), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n340_), .A2(new_n341_), .A3(new_n343_), .ZN(new_n344_));
  OR2_X1    g143(.A1(new_n344_), .A2(KEYINPUT21), .ZN(new_n345_));
  XOR2_X1   g144(.A(G211gat), .B(G218gat), .Z(new_n346_));
  NAND2_X1  g145(.A1(new_n342_), .A2(G204gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(new_n341_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n346_), .B1(KEYINPUT21), .B2(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G211gat), .B(G218gat), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT21), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  AOI22_X1  g151(.A1(new_n345_), .A2(new_n349_), .B1(new_n344_), .B2(new_n352_), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n333_), .B(new_n336_), .C1(new_n337_), .C2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n293_), .A2(KEYINPUT29), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n353_), .B1(KEYINPUT90), .B2(new_n335_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n336_), .A2(new_n333_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n355_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n354_), .A2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G78gat), .B(G106gat), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n354_), .A2(new_n358_), .A3(new_n360_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n332_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT92), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n360_), .B1(new_n354_), .B2(new_n358_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT91), .ZN(new_n367_));
  OAI211_X1 g166(.A(new_n332_), .B(new_n363_), .C1(new_n366_), .C2(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n362_), .A2(KEYINPUT91), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n365_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n330_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n331_), .ZN(new_n372_));
  AND3_X1   g171(.A1(new_n371_), .A2(new_n363_), .A3(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n362_), .A2(KEYINPUT91), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n366_), .A2(new_n367_), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n373_), .A2(new_n374_), .A3(KEYINPUT92), .A4(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n364_), .B1(new_n370_), .B2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G226gat), .A2(G233gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT19), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n353_), .B1(new_n233_), .B2(new_n244_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(G183gat), .A2(G190gat), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n207_), .A2(KEYINPUT23), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n205_), .A2(KEYINPUT81), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n203_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n204_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n381_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n219_), .B1(new_n235_), .B2(new_n237_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(KEYINPUT93), .A2(KEYINPUT24), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(KEYINPUT93), .A2(KEYINPUT24), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n211_), .B(new_n219_), .C1(new_n389_), .C2(new_n390_), .ZN(new_n391_));
  AND2_X1   g190(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n392_));
  OAI211_X1 g191(.A(new_n228_), .B(new_n230_), .C1(new_n392_), .C2(new_n224_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n390_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(G169gat), .A2(G176gat), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n394_), .A2(new_n395_), .A3(new_n388_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n391_), .A2(new_n393_), .A3(new_n396_), .ZN(new_n397_));
  OAI22_X1  g196(.A1(new_n386_), .A2(new_n387_), .B1(new_n397_), .B2(new_n243_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n348_), .A2(KEYINPUT21), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n399_), .B(new_n350_), .C1(new_n344_), .C2(KEYINPUT21), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n352_), .A2(new_n344_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(KEYINPUT20), .B1(new_n398_), .B2(new_n402_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n379_), .B1(new_n380_), .B2(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n233_), .A2(new_n244_), .A3(new_n353_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT20), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n406_), .B1(new_n398_), .B2(new_n402_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n405_), .A2(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n404_), .B1(new_n379_), .B2(new_n408_), .ZN(new_n409_));
  XOR2_X1   g208(.A(G8gat), .B(G36gat), .Z(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(KEYINPUT18), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G64gat), .B(G92gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n409_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n408_), .A2(new_n379_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n245_), .A2(new_n402_), .ZN(new_n417_));
  OAI22_X1  g216(.A1(new_n217_), .A2(new_n204_), .B1(G183gat), .B2(G190gat), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n391_), .A2(new_n393_), .A3(new_n396_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n243_), .ZN(new_n420_));
  AOI22_X1  g219(.A1(new_n239_), .A2(new_n418_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n406_), .B1(new_n421_), .B2(new_n353_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n379_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n417_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n416_), .A2(new_n424_), .A3(new_n413_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n415_), .A2(KEYINPUT27), .A3(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT98), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NOR3_X1   g227(.A1(new_n380_), .A2(new_n403_), .A3(new_n379_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n423_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n414_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(new_n425_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT27), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n415_), .A2(KEYINPUT98), .A3(KEYINPUT27), .A4(new_n425_), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n428_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n377_), .A2(new_n436_), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n323_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT99), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n370_), .A2(new_n376_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n364_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n413_), .A2(KEYINPUT32), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n443_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n444_), .B1(new_n409_), .B2(new_n443_), .ZN(new_n445_));
  AND3_X1   g244(.A1(new_n308_), .A2(new_n309_), .A3(new_n314_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n314_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n445_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT97), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n322_), .A2(KEYINPUT97), .A3(new_n445_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT33), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n321_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT95), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT95), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n321_), .A2(new_n455_), .A3(new_n452_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n454_), .A2(new_n456_), .ZN(new_n457_));
  AND2_X1   g256(.A1(new_n431_), .A2(new_n425_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n294_), .A2(new_n302_), .A3(new_n319_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(new_n315_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT96), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT96), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n459_), .A2(new_n462_), .A3(new_n315_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n303_), .A2(new_n304_), .A3(new_n318_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n461_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n308_), .A2(KEYINPUT33), .A3(new_n309_), .A4(new_n314_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n458_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  OAI211_X1 g266(.A(new_n450_), .B(new_n451_), .C1(new_n457_), .C2(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n260_), .B1(new_n442_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n322_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n377_), .B1(new_n470_), .B2(new_n436_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n439_), .B1(new_n469_), .B2(new_n471_), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n470_), .A2(new_n428_), .A3(new_n434_), .A4(new_n435_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n442_), .A2(new_n473_), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n458_), .A2(new_n465_), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n475_), .A2(new_n466_), .A3(new_n454_), .A4(new_n456_), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n377_), .A2(new_n476_), .A3(new_n450_), .A4(new_n451_), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n474_), .A2(new_n477_), .A3(KEYINPUT99), .A4(new_n260_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n438_), .B1(new_n472_), .B2(new_n478_), .ZN(new_n479_));
  XOR2_X1   g278(.A(G127gat), .B(G155gat), .Z(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT16), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G183gat), .B(G211gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n481_), .B(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT17), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G57gat), .B(G64gat), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT67), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT11), .ZN(new_n489_));
  XOR2_X1   g288(.A(G71gat), .B(G78gat), .Z(new_n490_));
  OR2_X1    g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n486_), .B(KEYINPUT67), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT11), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n489_), .A2(new_n494_), .A3(new_n490_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n491_), .A2(new_n495_), .ZN(new_n496_));
  AND2_X1   g295(.A1(G231gat), .A2(G233gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT77), .ZN(new_n499_));
  OR2_X1    g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G15gat), .B(G22gat), .ZN(new_n501_));
  INV_X1    g300(.A(G1gat), .ZN(new_n502_));
  INV_X1    g301(.A(G8gat), .ZN(new_n503_));
  OAI21_X1  g302(.A(KEYINPUT14), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n501_), .A2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G1gat), .B(G8gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n498_), .A2(new_n499_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n500_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n508_), .B1(new_n500_), .B2(new_n509_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n485_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n500_), .A2(new_n509_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(new_n507_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n483_), .B(KEYINPUT17), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n515_), .A2(new_n510_), .A3(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n513_), .A2(new_n517_), .A3(KEYINPUT78), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT78), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n515_), .A2(new_n519_), .A3(new_n510_), .A4(new_n516_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT37), .ZN(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G232gat), .A2(G233gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n523_), .B(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT35), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT74), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  OAI21_X1  g329(.A(KEYINPUT74), .B1(new_n526_), .B2(new_n527_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(KEYINPUT64), .B(G92gat), .ZN(new_n532_));
  AOI21_X1  g331(.A(KEYINPUT9), .B1(new_n532_), .B2(G85gat), .ZN(new_n533_));
  NAND3_X1  g332(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT65), .B1(new_n533_), .B2(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(KEYINPUT65), .B1(G85gat), .B2(G92gat), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n536_), .B1(new_n535_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G99gat), .A2(G106gat), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT6), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(G106gat), .ZN(new_n543_));
  XOR2_X1   g342(.A(KEYINPUT10), .B(G99gat), .Z(new_n544_));
  AOI21_X1  g343(.A(new_n542_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n539_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT8), .ZN(new_n547_));
  NOR2_X1   g346(.A1(G99gat), .A2(G106gat), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT7), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n542_), .B1(new_n550_), .B2(KEYINPUT66), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n551_), .B1(KEYINPUT66), .B2(new_n550_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G85gat), .B(G92gat), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n547_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n555_));
  OAI211_X1 g354(.A(new_n547_), .B(new_n554_), .C1(new_n550_), .C2(new_n542_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n546_), .B1(new_n555_), .B2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT68), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  XOR2_X1   g359(.A(G29gat), .B(G36gat), .Z(new_n561_));
  XOR2_X1   g360(.A(G43gat), .B(G50gat), .Z(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G29gat), .B(G36gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G43gat), .B(G50gat), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n563_), .A2(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT15), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n546_), .B(KEYINPUT68), .C1(new_n555_), .C2(new_n557_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n560_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n570_), .A2(KEYINPUT73), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT73), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n560_), .A2(new_n572_), .A3(new_n568_), .A4(new_n569_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n552_), .A2(new_n554_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(KEYINPUT8), .ZN(new_n575_));
  AOI22_X1  g374(.A1(new_n575_), .A2(new_n556_), .B1(new_n539_), .B2(new_n545_), .ZN(new_n576_));
  AOI22_X1  g375(.A1(new_n576_), .A2(new_n567_), .B1(new_n527_), .B2(new_n526_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n573_), .A2(new_n577_), .ZN(new_n578_));
  OAI211_X1 g377(.A(new_n530_), .B(new_n531_), .C1(new_n571_), .C2(new_n578_), .ZN(new_n579_));
  AND2_X1   g378(.A1(new_n573_), .A2(new_n577_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n570_), .A2(KEYINPUT73), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n580_), .A2(new_n529_), .A3(new_n528_), .A4(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G190gat), .B(G218gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT75), .ZN(new_n584_));
  XOR2_X1   g383(.A(G134gat), .B(G162gat), .Z(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT36), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n579_), .A2(new_n582_), .A3(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT36), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n586_), .A2(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n590_), .B1(new_n579_), .B2(new_n582_), .ZN(new_n591_));
  OAI211_X1 g390(.A(KEYINPUT76), .B(new_n522_), .C1(new_n588_), .C2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n579_), .A2(new_n582_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n590_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n579_), .A2(new_n582_), .A3(new_n587_), .ZN(new_n596_));
  OR2_X1    g395(.A1(new_n522_), .A2(KEYINPUT76), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n522_), .A2(KEYINPUT76), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n595_), .A2(new_n596_), .A3(new_n597_), .A4(new_n598_), .ZN(new_n599_));
  AND3_X1   g398(.A1(new_n521_), .A2(new_n592_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n568_), .A2(new_n507_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n508_), .A2(new_n567_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G229gat), .A2(G233gat), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n602_), .A2(new_n603_), .A3(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n507_), .A2(new_n566_), .A3(new_n563_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n603_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n604_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n605_), .A2(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G113gat), .B(G141gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G169gat), .B(G197gat), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n611_), .B(new_n612_), .Z(new_n613_));
  OR2_X1    g412(.A1(new_n613_), .A2(KEYINPUT79), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n610_), .B(new_n614_), .Z(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT71), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT13), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(KEYINPUT71), .A2(KEYINPUT13), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT12), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n496_), .A2(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n560_), .A2(new_n569_), .A3(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n621_), .B1(new_n576_), .B2(new_n496_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(G230gat), .A2(G233gat), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n576_), .A2(new_n496_), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n623_), .A2(new_n624_), .A3(new_n625_), .A4(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n576_), .A2(new_n496_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n491_), .A2(new_n495_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n558_), .A2(new_n629_), .ZN(new_n630_));
  OAI211_X1 g429(.A(G230gat), .B(G233gat), .C1(new_n628_), .C2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n627_), .A2(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(G120gat), .B(G148gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT5), .ZN(new_n634_));
  XNOR2_X1  g433(.A(G176gat), .B(G204gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT69), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n632_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT70), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n627_), .A2(new_n631_), .A3(new_n636_), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n639_), .A2(new_n640_), .A3(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n640_), .B1(new_n639_), .B2(new_n641_), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n619_), .B(new_n620_), .C1(new_n642_), .C2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n639_), .A2(new_n641_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(KEYINPUT70), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n639_), .A2(new_n640_), .A3(new_n641_), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n646_), .A2(new_n647_), .A3(new_n617_), .A4(new_n618_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n644_), .A2(new_n648_), .ZN(new_n649_));
  NOR4_X1   g448(.A1(new_n479_), .A2(new_n601_), .A3(new_n616_), .A4(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n650_), .A2(new_n502_), .A3(new_n322_), .ZN(new_n651_));
  XOR2_X1   g450(.A(new_n651_), .B(KEYINPUT100), .Z(new_n652_));
  OR2_X1    g451(.A1(new_n652_), .A2(KEYINPUT38), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(KEYINPUT38), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n588_), .A2(new_n591_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n479_), .A2(new_n655_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n644_), .A2(new_n648_), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n656_), .A2(new_n615_), .A3(new_n657_), .A4(new_n521_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT101), .ZN(new_n659_));
  OAI21_X1  g458(.A(G1gat), .B1(new_n659_), .B2(new_n470_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n653_), .A2(new_n654_), .A3(new_n660_), .ZN(G1324gat));
  OAI21_X1  g460(.A(G8gat), .B1(new_n658_), .B2(new_n436_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT39), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n436_), .A2(G8gat), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n650_), .A2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n663_), .A2(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n666_), .B(new_n667_), .ZN(G1325gat));
  INV_X1    g467(.A(KEYINPUT41), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT103), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT101), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n658_), .B(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(new_n259_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n670_), .B1(new_n673_), .B2(G15gat), .ZN(new_n674_));
  AOI211_X1 g473(.A(KEYINPUT103), .B(new_n255_), .C1(new_n672_), .C2(new_n259_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n669_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(G15gat), .B1(new_n659_), .B2(new_n260_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(KEYINPUT103), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n673_), .A2(new_n670_), .A3(G15gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n678_), .A2(KEYINPUT41), .A3(new_n679_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n650_), .A2(new_n255_), .A3(new_n259_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n676_), .A2(new_n680_), .A3(new_n681_), .ZN(G1326gat));
  INV_X1    g481(.A(G22gat), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n650_), .A2(new_n683_), .A3(new_n442_), .ZN(new_n684_));
  OAI21_X1  g483(.A(G22gat), .B1(new_n659_), .B2(new_n377_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n685_), .A2(KEYINPUT42), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n685_), .A2(KEYINPUT42), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n684_), .B1(new_n686_), .B2(new_n687_), .ZN(G1327gat));
  INV_X1    g487(.A(new_n438_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n450_), .A2(new_n451_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n455_), .B1(new_n321_), .B2(new_n452_), .ZN(new_n691_));
  AND3_X1   g490(.A1(new_n321_), .A2(new_n455_), .A3(new_n452_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n467_), .A2(new_n691_), .A3(new_n692_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n690_), .A2(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n259_), .B1(new_n694_), .B2(new_n377_), .ZN(new_n695_));
  AOI21_X1  g494(.A(KEYINPUT99), .B1(new_n695_), .B2(new_n474_), .ZN(new_n696_));
  AND4_X1   g495(.A1(KEYINPUT99), .A2(new_n474_), .A3(new_n477_), .A4(new_n260_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n689_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n655_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n699_), .A2(new_n521_), .ZN(new_n700_));
  AND4_X1   g499(.A1(new_n698_), .A2(new_n615_), .A3(new_n657_), .A4(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(G29gat), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n701_), .A2(new_n702_), .A3(new_n322_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT43), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n592_), .A2(new_n599_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n698_), .A2(new_n704_), .A3(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n705_), .ZN(new_n707_));
  OAI21_X1  g506(.A(KEYINPUT43), .B1(new_n479_), .B2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n708_), .ZN(new_n709_));
  NOR3_X1   g508(.A1(new_n649_), .A2(new_n616_), .A3(new_n521_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT104), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n711_), .B(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n702_), .B1(new_n714_), .B2(new_n322_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n715_), .A2(KEYINPUT105), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n715_), .A2(KEYINPUT105), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n703_), .B1(new_n716_), .B2(new_n717_), .ZN(G1328gat));
  INV_X1    g517(.A(G36gat), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT106), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n436_), .B(new_n720_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n701_), .A2(new_n719_), .A3(new_n721_), .ZN(new_n722_));
  XOR2_X1   g521(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n723_));
  XNOR2_X1  g522(.A(new_n722_), .B(new_n723_), .ZN(new_n724_));
  OR2_X1    g523(.A1(new_n711_), .A2(new_n713_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n711_), .A2(new_n713_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n436_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n724_), .B1(new_n727_), .B2(new_n719_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT46), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  OAI211_X1 g529(.A(KEYINPUT46), .B(new_n724_), .C1(new_n727_), .C2(new_n719_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(G1329gat));
  INV_X1    g531(.A(G43gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n701_), .A2(new_n733_), .A3(new_n259_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n260_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n734_), .B1(new_n735_), .B2(new_n733_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT47), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  OAI211_X1 g537(.A(KEYINPUT47), .B(new_n734_), .C1(new_n735_), .C2(new_n733_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(G1330gat));
  INV_X1    g539(.A(G50gat), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n701_), .A2(new_n741_), .A3(new_n442_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n377_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n742_), .B1(new_n743_), .B2(new_n741_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT108), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT108), .ZN(new_n746_));
  OAI211_X1 g545(.A(new_n746_), .B(new_n742_), .C1(new_n743_), .C2(new_n741_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n747_), .ZN(G1331gat));
  NOR4_X1   g547(.A1(new_n479_), .A2(new_n601_), .A3(new_n615_), .A4(new_n657_), .ZN(new_n749_));
  INV_X1    g548(.A(G57gat), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n749_), .A2(new_n750_), .A3(new_n322_), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n656_), .A2(new_n616_), .A3(new_n649_), .A4(new_n521_), .ZN(new_n752_));
  XOR2_X1   g551(.A(new_n752_), .B(KEYINPUT109), .Z(new_n753_));
  AND2_X1   g552(.A1(new_n753_), .A2(new_n322_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n751_), .B1(new_n754_), .B2(new_n750_), .ZN(G1332gat));
  INV_X1    g554(.A(G64gat), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n749_), .A2(new_n756_), .A3(new_n721_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n753_), .A2(new_n721_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(G64gat), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n759_), .A2(KEYINPUT48), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n759_), .A2(KEYINPUT48), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n757_), .B1(new_n760_), .B2(new_n761_), .ZN(G1333gat));
  INV_X1    g561(.A(G71gat), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n749_), .A2(new_n763_), .A3(new_n259_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n753_), .A2(new_n259_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(G71gat), .ZN(new_n766_));
  XOR2_X1   g565(.A(KEYINPUT110), .B(KEYINPUT49), .Z(new_n767_));
  AND2_X1   g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n766_), .A2(new_n767_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n764_), .B1(new_n768_), .B2(new_n769_), .ZN(G1334gat));
  INV_X1    g569(.A(G78gat), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n749_), .A2(new_n771_), .A3(new_n442_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n753_), .A2(new_n442_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(G78gat), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n774_), .A2(KEYINPUT50), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n774_), .A2(KEYINPUT50), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n772_), .B1(new_n775_), .B2(new_n776_), .ZN(G1335gat));
  INV_X1    g576(.A(new_n521_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n649_), .A2(new_n616_), .A3(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT111), .ZN(new_n780_));
  OR2_X1    g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n780_), .ZN(new_n782_));
  AOI22_X1  g581(.A1(new_n706_), .A2(new_n708_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  XOR2_X1   g582(.A(new_n783_), .B(KEYINPUT112), .Z(new_n784_));
  OAI21_X1  g583(.A(G85gat), .B1(new_n784_), .B2(new_n470_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n479_), .A2(new_n615_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n700_), .A2(new_n649_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  OR3_X1    g587(.A1(new_n788_), .A2(G85gat), .A3(new_n470_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n785_), .A2(new_n789_), .ZN(G1336gat));
  INV_X1    g589(.A(G92gat), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n791_), .B1(new_n788_), .B2(new_n436_), .ZN(new_n792_));
  XOR2_X1   g591(.A(new_n792_), .B(KEYINPUT113), .Z(new_n793_));
  INV_X1    g592(.A(new_n784_), .ZN(new_n794_));
  AND2_X1   g593(.A1(new_n721_), .A2(new_n532_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n793_), .B1(new_n794_), .B2(new_n795_), .ZN(G1337gat));
  OAI21_X1  g595(.A(G99gat), .B1(new_n784_), .B2(new_n260_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n788_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n798_), .A2(new_n259_), .A3(new_n544_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n797_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT51), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT51), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n797_), .A2(new_n802_), .A3(new_n799_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n801_), .A2(new_n803_), .ZN(G1338gat));
  NAND2_X1  g603(.A1(new_n781_), .A2(new_n782_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n709_), .A2(KEYINPUT114), .A3(new_n442_), .A4(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(G106gat), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT114), .B1(new_n783_), .B2(new_n442_), .ZN(new_n808_));
  OAI21_X1  g607(.A(KEYINPUT115), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n709_), .A2(new_n442_), .A3(new_n805_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT114), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT115), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n812_), .A2(new_n813_), .A3(G106gat), .A4(new_n806_), .ZN(new_n814_));
  AND3_X1   g613(.A1(new_n809_), .A2(KEYINPUT52), .A3(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n816_));
  OAI211_X1 g615(.A(KEYINPUT115), .B(new_n816_), .C1(new_n807_), .C2(new_n808_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n798_), .A2(new_n543_), .A3(new_n442_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(KEYINPUT53), .B1(new_n815_), .B2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n809_), .A2(KEYINPUT52), .A3(new_n814_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT53), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n821_), .A2(new_n822_), .A3(new_n817_), .A4(new_n818_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n820_), .A2(new_n823_), .ZN(G1339gat));
  INV_X1    g623(.A(KEYINPUT58), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT12), .B1(new_n558_), .B2(new_n629_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n826_), .A2(new_n630_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n625_), .B1(new_n827_), .B2(new_n623_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n627_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n827_), .A2(KEYINPUT55), .A3(new_n625_), .A4(new_n623_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n637_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT56), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n602_), .A2(new_n603_), .A3(new_n608_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n607_), .A2(new_n604_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n613_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n837_), .B1(new_n613_), .B2(new_n610_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(KEYINPUT120), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n839_), .A2(new_n641_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n834_), .A2(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n832_), .A2(new_n833_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n825_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n830_), .A2(new_n831_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n638_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(KEYINPUT56), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n846_), .A2(KEYINPUT58), .A3(new_n834_), .A4(new_n840_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n843_), .A2(new_n705_), .A3(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT119), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n845_), .A2(new_n849_), .A3(KEYINPUT56), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n833_), .B1(new_n832_), .B2(KEYINPUT119), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n641_), .A2(new_n615_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(KEYINPUT118), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n850_), .A2(new_n851_), .A3(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n646_), .A2(new_n647_), .A3(new_n839_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n655_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n848_), .B1(new_n856_), .B2(KEYINPUT57), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n858_));
  AOI211_X1 g657(.A(new_n858_), .B(new_n655_), .C1(new_n854_), .C2(new_n855_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n778_), .B1(new_n857_), .B2(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n600_), .A2(new_n616_), .A3(new_n657_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(KEYINPUT117), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT117), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n600_), .A2(new_n657_), .A3(new_n863_), .A4(new_n616_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(KEYINPUT116), .B(KEYINPUT54), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n862_), .A2(new_n864_), .A3(new_n866_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n861_), .A2(KEYINPUT117), .A3(new_n865_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n860_), .A2(new_n867_), .A3(new_n868_), .ZN(new_n869_));
  AND3_X1   g668(.A1(new_n437_), .A2(new_n322_), .A3(new_n259_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT59), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n869_), .A2(KEYINPUT59), .A3(new_n870_), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(G113gat), .B1(new_n875_), .B2(new_n616_), .ZN(new_n876_));
  OR3_X1    g675(.A1(new_n871_), .A2(G113gat), .A3(new_n616_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(G1340gat));
  INV_X1    g677(.A(new_n871_), .ZN(new_n879_));
  XOR2_X1   g678(.A(KEYINPUT121), .B(G120gat), .Z(new_n880_));
  OAI21_X1  g679(.A(new_n880_), .B1(new_n657_), .B2(KEYINPUT60), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n879_), .B(new_n881_), .C1(KEYINPUT60), .C2(new_n880_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n875_), .A2(new_n657_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n883_), .B2(new_n880_), .ZN(G1341gat));
  INV_X1    g683(.A(G127gat), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n879_), .A2(new_n885_), .A3(new_n521_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n778_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n887_), .B2(new_n885_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(KEYINPUT122), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT122), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n890_), .B(new_n886_), .C1(new_n887_), .C2(new_n885_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n891_), .ZN(G1342gat));
  OAI21_X1  g691(.A(G134gat), .B1(new_n875_), .B2(new_n707_), .ZN(new_n893_));
  OR3_X1    g692(.A1(new_n871_), .A2(G134gat), .A3(new_n699_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(G1343gat));
  NOR4_X1   g694(.A1(new_n721_), .A2(new_n377_), .A3(new_n470_), .A4(new_n259_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n869_), .A2(new_n896_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n897_), .A2(new_n616_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(new_n262_), .ZN(G1344gat));
  NOR2_X1   g698(.A1(new_n897_), .A2(new_n657_), .ZN(new_n900_));
  XOR2_X1   g699(.A(KEYINPUT123), .B(G148gat), .Z(new_n901_));
  XNOR2_X1  g700(.A(new_n900_), .B(new_n901_), .ZN(G1345gat));
  NAND3_X1  g701(.A1(new_n869_), .A2(new_n521_), .A3(new_n896_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(KEYINPUT124), .ZN(new_n904_));
  XNOR2_X1  g703(.A(KEYINPUT61), .B(G155gat), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n904_), .B(new_n905_), .ZN(G1346gat));
  OAI21_X1  g705(.A(G162gat), .B1(new_n897_), .B2(new_n707_), .ZN(new_n907_));
  OR2_X1    g706(.A1(new_n699_), .A2(G162gat), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n907_), .B1(new_n897_), .B2(new_n908_), .ZN(G1347gat));
  AND3_X1   g708(.A1(new_n721_), .A2(new_n377_), .A3(new_n323_), .ZN(new_n910_));
  AND2_X1   g709(.A1(new_n869_), .A2(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n615_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n912_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n913_), .B1(new_n237_), .B2(new_n912_), .ZN(new_n914_));
  AOI21_X1  g713(.A(KEYINPUT62), .B1(new_n912_), .B2(G169gat), .ZN(new_n915_));
  OR2_X1    g714(.A1(new_n914_), .A2(new_n915_), .ZN(G1348gat));
  INV_X1    g715(.A(new_n911_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n917_), .A2(new_n657_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n918_), .A2(new_n235_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n919_), .B1(G176gat), .B2(new_n918_), .ZN(G1349gat));
  NOR2_X1   g719(.A1(new_n917_), .A2(new_n778_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n921_), .A2(new_n240_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n392_), .A2(new_n224_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n922_), .B1(new_n923_), .B2(new_n921_), .ZN(G1350gat));
  NAND3_X1  g723(.A1(new_n911_), .A2(new_n231_), .A3(new_n655_), .ZN(new_n925_));
  OAI21_X1  g724(.A(G190gat), .B1(new_n917_), .B2(new_n707_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT125), .ZN(new_n927_));
  AND2_X1   g726(.A1(new_n926_), .A2(new_n927_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n926_), .A2(new_n927_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n925_), .B1(new_n928_), .B2(new_n929_), .ZN(G1351gat));
  NAND3_X1  g729(.A1(new_n442_), .A2(new_n260_), .A3(new_n470_), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT126), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n721_), .B1(new_n931_), .B2(new_n932_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n933_), .B1(new_n932_), .B2(new_n931_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n869_), .A2(new_n934_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n935_), .A2(new_n616_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n936_), .B(new_n342_), .ZN(G1352gat));
  NOR2_X1   g736(.A1(new_n935_), .A2(new_n657_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n938_), .A2(new_n939_), .ZN(new_n940_));
  XOR2_X1   g739(.A(KEYINPUT127), .B(G204gat), .Z(new_n941_));
  OAI21_X1  g740(.A(new_n940_), .B1(new_n938_), .B2(new_n941_), .ZN(G1353gat));
  NAND3_X1  g741(.A1(new_n869_), .A2(new_n521_), .A3(new_n934_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n944_));
  AND2_X1   g743(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n945_));
  NOR3_X1   g744(.A1(new_n943_), .A2(new_n944_), .A3(new_n945_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n946_), .B1(new_n943_), .B2(new_n944_), .ZN(G1354gat));
  OAI21_X1  g746(.A(G218gat), .B1(new_n935_), .B2(new_n707_), .ZN(new_n948_));
  OR2_X1    g747(.A1(new_n699_), .A2(G218gat), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n948_), .B1(new_n935_), .B2(new_n949_), .ZN(G1355gat));
endmodule


