//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 0 0 1 0 1 1 0 1 1 1 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 0 1 0 0 1 0 1 1 1 1 0 1 1 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n739_, new_n740_, new_n741_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n770_,
    new_n771_, new_n772_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n781_, new_n782_, new_n784_, new_n785_,
    new_n786_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n857_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n873_, new_n874_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n907_, new_n908_, new_n909_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n918_,
    new_n919_, new_n920_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n932_,
    new_n933_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n944_, new_n945_;
  XNOR2_X1  g000(.A(G211gat), .B(G218gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT21), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G197gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT87), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT87), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(G197gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G204gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(G197gat), .A2(G204gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n204_), .A2(new_n210_), .A3(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT88), .B(KEYINPUT21), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n215_), .B1(new_n210_), .B2(new_n212_), .ZN(new_n216_));
  INV_X1    g015(.A(G204gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n206_), .A2(new_n208_), .A3(new_n217_), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n203_), .B1(G197gat), .B2(G204gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(new_n202_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n213_), .B1(new_n216_), .B2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT89), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n217_), .B1(new_n206_), .B2(new_n208_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n214_), .B1(new_n224_), .B2(new_n211_), .ZN(new_n225_));
  INV_X1    g024(.A(G218gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(G211gat), .ZN(new_n227_));
  INV_X1    g026(.A(G211gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(G218gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n227_), .A2(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n230_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n224_), .A2(new_n211_), .ZN(new_n232_));
  AOI22_X1  g031(.A1(new_n225_), .A2(new_n231_), .B1(new_n232_), .B2(new_n204_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT89), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G228gat), .A2(G233gat), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G155gat), .A2(G162gat), .ZN(new_n238_));
  NOR2_X1   g037(.A1(G155gat), .A2(G162gat), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n238_), .B1(new_n239_), .B2(KEYINPUT1), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT1), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n241_), .A2(KEYINPUT85), .A3(G155gat), .A4(G162gat), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT85), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n243_), .B1(new_n238_), .B2(KEYINPUT1), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n240_), .A2(new_n242_), .A3(new_n244_), .ZN(new_n245_));
  XOR2_X1   g044(.A(G141gat), .B(G148gat), .Z(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n248_));
  INV_X1    g047(.A(G141gat), .ZN(new_n249_));
  INV_X1    g048(.A(G148gat), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n248_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G141gat), .A2(G148gat), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT2), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n255_));
  OAI21_X1  g054(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n251_), .A2(new_n254_), .A3(new_n255_), .A4(new_n256_), .ZN(new_n257_));
  XOR2_X1   g056(.A(G155gat), .B(G162gat), .Z(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n247_), .A2(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n237_), .B1(new_n260_), .B2(KEYINPUT29), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n223_), .A2(new_n235_), .A3(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(G78gat), .ZN(new_n263_));
  AOI22_X1  g062(.A1(new_n245_), .A2(new_n246_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n264_));
  XOR2_X1   g063(.A(KEYINPUT90), .B(KEYINPUT29), .Z(new_n265_));
  NOR2_X1   g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n237_), .B1(new_n266_), .B2(new_n233_), .ZN(new_n267_));
  AND3_X1   g066(.A1(new_n262_), .A2(new_n263_), .A3(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n263_), .B1(new_n262_), .B2(new_n267_), .ZN(new_n269_));
  OAI21_X1  g068(.A(G106gat), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  XOR2_X1   g069(.A(G22gat), .B(G50gat), .Z(new_n271_));
  XOR2_X1   g070(.A(KEYINPUT86), .B(KEYINPUT28), .Z(new_n272_));
  OAI21_X1  g071(.A(new_n272_), .B1(new_n260_), .B2(KEYINPUT29), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT29), .ZN(new_n274_));
  INV_X1    g073(.A(new_n272_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n264_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n271_), .B1(new_n273_), .B2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT91), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n273_), .A2(new_n271_), .A3(new_n276_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n278_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n225_), .A2(new_n231_), .ZN(new_n283_));
  AND3_X1   g082(.A1(new_n283_), .A2(new_n234_), .A3(new_n213_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n234_), .B1(new_n283_), .B2(new_n213_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n236_), .B1(new_n264_), .B2(new_n274_), .ZN(new_n286_));
  NOR3_X1   g085(.A1(new_n284_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  OR2_X1    g086(.A1(new_n264_), .A2(new_n265_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n236_), .B1(new_n288_), .B2(new_n222_), .ZN(new_n289_));
  OAI21_X1  g088(.A(G78gat), .B1(new_n287_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(G106gat), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n262_), .A2(new_n263_), .A3(new_n267_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n290_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  AND3_X1   g092(.A1(new_n270_), .A2(new_n282_), .A3(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n280_), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT91), .B1(new_n295_), .B2(new_n277_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(new_n281_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n297_), .B1(new_n270_), .B2(new_n293_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n294_), .A2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G1gat), .B(G29gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(G85gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT0), .B(G57gat), .ZN(new_n302_));
  XOR2_X1   g101(.A(new_n301_), .B(new_n302_), .Z(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G225gat), .A2(G233gat), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(G134gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(G127gat), .ZN(new_n308_));
  INV_X1    g107(.A(G127gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(G134gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(G120gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(G113gat), .ZN(new_n313_));
  INV_X1    g112(.A(G113gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(G120gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n311_), .A2(new_n316_), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n308_), .A2(new_n310_), .A3(new_n313_), .A4(new_n315_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n260_), .A2(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n306_), .B1(new_n321_), .B2(KEYINPUT4), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n247_), .A2(new_n319_), .A3(new_n259_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n321_), .A2(KEYINPUT95), .A3(new_n323_), .ZN(new_n324_));
  NOR3_X1   g123(.A1(new_n264_), .A2(KEYINPUT95), .A3(new_n319_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n324_), .A2(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n322_), .B1(new_n327_), .B2(KEYINPUT4), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n306_), .B1(new_n324_), .B2(new_n326_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n304_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n327_), .A2(new_n305_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT4), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n332_), .B1(new_n324_), .B2(new_n326_), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n331_), .B(new_n303_), .C1(new_n333_), .C2(new_n322_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n330_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(G190gat), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT79), .B1(new_n337_), .B2(KEYINPUT26), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT79), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT26), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n339_), .A2(new_n340_), .A3(G190gat), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n338_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT78), .ZN(new_n343_));
  INV_X1    g142(.A(G183gat), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n343_), .B1(new_n344_), .B2(KEYINPUT25), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT25), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n346_), .A2(KEYINPUT78), .A3(G183gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n337_), .A2(KEYINPUT26), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n344_), .A2(KEYINPUT25), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n345_), .A2(new_n347_), .A3(new_n348_), .A4(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT80), .B1(new_n342_), .B2(new_n350_), .ZN(new_n351_));
  AND3_X1   g150(.A1(new_n347_), .A2(new_n348_), .A3(new_n349_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT80), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n338_), .A2(new_n341_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n352_), .A2(new_n353_), .A3(new_n354_), .A4(new_n345_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G183gat), .A2(G190gat), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT23), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(G169gat), .ZN(new_n361_));
  INV_X1    g160(.A(G176gat), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n361_), .A2(new_n362_), .A3(KEYINPUT81), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT81), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n364_), .B1(G169gat), .B2(G176gat), .ZN(new_n365_));
  AND2_X1   g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT24), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n367_), .B1(G169gat), .B2(G176gat), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n360_), .B1(new_n366_), .B2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n363_), .A2(new_n365_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(new_n367_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n351_), .A2(new_n355_), .A3(new_n369_), .A4(new_n371_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(G169gat), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n358_), .B(new_n359_), .C1(G183gat), .C2(G190gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n372_), .A2(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G71gat), .B(G99gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(G43gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n377_), .B(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G227gat), .A2(G233gat), .ZN(new_n381_));
  INV_X1    g180(.A(G15gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(KEYINPUT30), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n380_), .B(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT83), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n319_), .B(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n386_), .A2(new_n387_), .A3(new_n389_), .ZN(new_n390_));
  OR2_X1    g189(.A1(new_n380_), .A2(new_n384_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n380_), .A2(new_n384_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n391_), .A2(new_n387_), .A3(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n389_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n386_), .A2(new_n387_), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n336_), .B(new_n390_), .C1(new_n395_), .C2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G226gat), .A2(G233gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT19), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT93), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n374_), .A2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n373_), .B(new_n361_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT93), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n402_), .A2(new_n404_), .A3(new_n375_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n367_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n369_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n346_), .A2(G183gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(new_n349_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n340_), .A2(G190gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(new_n348_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT92), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n410_), .A2(new_n348_), .A3(KEYINPUT92), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n409_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n405_), .B1(new_n407_), .B2(new_n415_), .ZN(new_n416_));
  OAI211_X1 g215(.A(KEYINPUT20), .B(new_n400_), .C1(new_n416_), .C2(new_n222_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n284_), .A2(new_n285_), .ZN(new_n419_));
  AOI21_X1  g218(.A(KEYINPUT94), .B1(new_n419_), .B2(new_n377_), .ZN(new_n420_));
  AND4_X1   g219(.A1(KEYINPUT94), .A2(new_n377_), .A3(new_n223_), .A4(new_n235_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n418_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  OAI211_X1 g221(.A(new_n376_), .B(new_n372_), .C1(new_n284_), .C2(new_n285_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT20), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n424_), .B1(new_n416_), .B2(new_n222_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n400_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G8gat), .B(G36gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(KEYINPUT18), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G64gat), .B(G92gat), .ZN(new_n430_));
  XOR2_X1   g229(.A(new_n429_), .B(new_n430_), .Z(new_n431_));
  NAND3_X1  g230(.A1(new_n422_), .A2(new_n427_), .A3(new_n431_), .ZN(new_n432_));
  AND3_X1   g231(.A1(new_n423_), .A2(new_n425_), .A3(new_n400_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n416_), .A2(new_n222_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n434_), .A2(new_n424_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n435_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n433_), .B1(new_n436_), .B2(new_n399_), .ZN(new_n437_));
  OAI211_X1 g236(.A(KEYINPUT27), .B(new_n432_), .C1(new_n437_), .C2(new_n431_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(KEYINPUT97), .B(KEYINPUT27), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n377_), .A2(new_n223_), .A3(new_n235_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT94), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n419_), .A2(KEYINPUT94), .A3(new_n377_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n417_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n431_), .ZN(new_n446_));
  NOR3_X1   g245(.A1(new_n445_), .A2(new_n426_), .A3(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n431_), .B1(new_n422_), .B2(new_n427_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n440_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n438_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT99), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT99), .ZN(new_n452_));
  INV_X1    g251(.A(new_n438_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n449_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n452_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  AOI211_X1 g254(.A(new_n299_), .B(new_n397_), .C1(new_n451_), .C2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n390_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT84), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT84), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n459_), .B(new_n390_), .C1(new_n395_), .C2(new_n396_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n458_), .A2(new_n460_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n299_), .A2(new_n449_), .A3(new_n438_), .A4(new_n336_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n431_), .A2(KEYINPUT32), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n422_), .A2(new_n427_), .A3(new_n463_), .ZN(new_n464_));
  OAI211_X1 g263(.A(new_n335_), .B(new_n464_), .C1(new_n437_), .C2(new_n463_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n446_), .B1(new_n445_), .B2(new_n426_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n323_), .A2(KEYINPUT95), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n264_), .A2(new_n319_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(KEYINPUT4), .B1(new_n469_), .B2(new_n325_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n322_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n329_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT33), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n304_), .A2(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n306_), .B1(new_n468_), .B2(new_n332_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n470_), .A2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n303_), .B1(new_n327_), .B2(new_n306_), .ZN(new_n477_));
  AOI22_X1  g276(.A1(new_n472_), .A2(new_n474_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n334_), .A2(new_n473_), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n466_), .A2(new_n478_), .A3(new_n432_), .A4(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n270_), .A2(new_n293_), .A3(new_n282_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n270_), .A2(new_n293_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n297_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  AOI22_X1  g283(.A1(new_n465_), .A2(new_n480_), .B1(new_n481_), .B2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n462_), .B1(new_n485_), .B2(KEYINPUT96), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n465_), .A2(new_n480_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n484_), .A2(new_n481_), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n487_), .A2(new_n488_), .A3(KEYINPUT96), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n461_), .B1(new_n486_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(KEYINPUT98), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT98), .ZN(new_n492_));
  OAI211_X1 g291(.A(new_n492_), .B(new_n461_), .C1(new_n486_), .C2(new_n489_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n456_), .B1(new_n491_), .B2(new_n493_), .ZN(new_n494_));
  XOR2_X1   g293(.A(KEYINPUT72), .B(G1gat), .Z(new_n495_));
  INV_X1    g294(.A(G8gat), .ZN(new_n496_));
  OAI21_X1  g295(.A(KEYINPUT14), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G15gat), .B(G22gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G1gat), .B(G8gat), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n497_), .A2(new_n498_), .A3(new_n500_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G29gat), .B(G36gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G43gat), .B(G50gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n504_), .A2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT75), .ZN(new_n509_));
  OR2_X1    g308(.A1(new_n504_), .A2(new_n507_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G229gat), .A2(G233gat), .ZN(new_n513_));
  OAI21_X1  g312(.A(KEYINPUT76), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT76), .ZN(new_n515_));
  INV_X1    g314(.A(new_n513_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n511_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n507_), .B(KEYINPUT15), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n518_), .A2(new_n503_), .A3(new_n502_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n509_), .A2(new_n513_), .A3(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n514_), .A2(new_n517_), .A3(new_n520_), .ZN(new_n521_));
  XOR2_X1   g320(.A(G113gat), .B(G141gat), .Z(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(KEYINPUT77), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G169gat), .B(G197gat), .ZN(new_n524_));
  XOR2_X1   g323(.A(new_n523_), .B(new_n524_), .Z(new_n525_));
  NAND2_X1  g324(.A1(new_n521_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n525_), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n514_), .A2(new_n517_), .A3(new_n520_), .A4(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n526_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT67), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT12), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G85gat), .B(G92gat), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n533_), .B1(KEYINPUT9), .B2(G92gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n535_));
  OR2_X1    g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(new_n535_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G99gat), .A2(G106gat), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT6), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  XOR2_X1   g339(.A(KEYINPUT10), .B(G99gat), .Z(new_n541_));
  AOI21_X1  g340(.A(new_n540_), .B1(new_n291_), .B2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n536_), .A2(new_n537_), .A3(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(G99gat), .A2(G106gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT7), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n538_), .B(KEYINPUT6), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT65), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n545_), .A2(KEYINPUT65), .A3(new_n546_), .ZN(new_n550_));
  AOI211_X1 g349(.A(KEYINPUT8), .B(new_n533_), .C1(new_n549_), .C2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT8), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT66), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n540_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n546_), .A2(KEYINPUT66), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n554_), .A2(new_n555_), .A3(new_n545_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n533_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n552_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n543_), .B1(new_n551_), .B2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G57gat), .B(G64gat), .ZN(new_n560_));
  OR2_X1    g359(.A1(new_n560_), .A2(KEYINPUT11), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(KEYINPUT11), .ZN(new_n562_));
  XOR2_X1   g361(.A(G71gat), .B(G78gat), .Z(new_n563_));
  NAND3_X1  g362(.A1(new_n561_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n562_), .A2(new_n563_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n532_), .B1(new_n559_), .B2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n543_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n549_), .A2(new_n550_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n570_), .A2(new_n552_), .A3(new_n557_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n556_), .A2(new_n557_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(KEYINPUT8), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n569_), .B1(new_n571_), .B2(new_n573_), .ZN(new_n574_));
  OAI22_X1  g373(.A1(new_n574_), .A2(new_n566_), .B1(new_n531_), .B2(KEYINPUT12), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n531_), .A2(KEYINPUT12), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n559_), .A2(new_n567_), .A3(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n568_), .B1(new_n575_), .B2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G230gat), .A2(G233gat), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n574_), .B(new_n566_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n581_), .A2(G230gat), .A3(G233gat), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  XOR2_X1   g382(.A(G120gat), .B(G148gat), .Z(new_n584_));
  XNOR2_X1  g383(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G176gat), .B(G204gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n583_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n588_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n580_), .A2(new_n582_), .A3(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n589_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n593_), .A2(KEYINPUT13), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(KEYINPUT13), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n559_), .A2(new_n518_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n574_), .A2(new_n507_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(G232gat), .A2(G233gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT34), .ZN(new_n600_));
  OR2_X1    g399(.A1(new_n600_), .A2(KEYINPUT35), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n597_), .A2(new_n598_), .A3(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(KEYINPUT35), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n603_), .B(KEYINPUT69), .Z(new_n604_));
  OR2_X1    g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n602_), .A2(new_n604_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  XOR2_X1   g406(.A(G190gat), .B(G218gat), .Z(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT70), .ZN(new_n609_));
  XOR2_X1   g408(.A(G134gat), .B(G162gat), .Z(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT36), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n607_), .A2(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n611_), .B(new_n612_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n605_), .A2(new_n615_), .A3(new_n606_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n614_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT71), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n617_), .A2(new_n618_), .A3(KEYINPUT37), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n618_), .A2(KEYINPUT37), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(KEYINPUT37), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n614_), .A2(new_n616_), .A3(new_n620_), .A4(new_n621_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n619_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(G231gat), .A2(G233gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n566_), .B(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(new_n504_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(KEYINPUT74), .ZN(new_n627_));
  XOR2_X1   g426(.A(G127gat), .B(G155gat), .Z(new_n628_));
  XNOR2_X1  g427(.A(G183gat), .B(G211gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n628_), .B(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(KEYINPUT17), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n627_), .B(new_n633_), .ZN(new_n634_));
  OR3_X1    g433(.A1(new_n626_), .A2(KEYINPUT17), .A3(new_n632_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n623_), .A2(new_n636_), .ZN(new_n637_));
  NOR4_X1   g436(.A1(new_n494_), .A2(new_n530_), .A3(new_n596_), .A4(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n638_), .A2(new_n335_), .A3(new_n495_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT38), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT100), .ZN(new_n642_));
  INV_X1    g441(.A(new_n596_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(new_n529_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n636_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n494_), .A2(new_n617_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  OAI21_X1  g447(.A(G1gat), .B1(new_n648_), .B2(new_n336_), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n649_), .B(KEYINPUT101), .Z(new_n650_));
  NAND2_X1  g449(.A1(new_n639_), .A2(new_n640_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT102), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n642_), .A2(new_n650_), .A3(new_n652_), .ZN(G1324gat));
  INV_X1    g452(.A(new_n451_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n455_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  OAI21_X1  g456(.A(G8gat), .B1(new_n648_), .B2(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT39), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n638_), .A2(new_n496_), .A3(new_n656_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n661_), .B(new_n662_), .ZN(G1325gat));
  OAI21_X1  g462(.A(G15gat), .B1(new_n648_), .B2(new_n461_), .ZN(new_n664_));
  XOR2_X1   g463(.A(new_n664_), .B(KEYINPUT41), .Z(new_n665_));
  INV_X1    g464(.A(new_n461_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n638_), .A2(new_n382_), .A3(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(G1326gat));
  OAI21_X1  g467(.A(G22gat), .B1(new_n648_), .B2(new_n488_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT42), .ZN(new_n670_));
  INV_X1    g469(.A(G22gat), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n638_), .A2(new_n671_), .A3(new_n299_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n672_), .ZN(G1327gat));
  INV_X1    g472(.A(KEYINPUT106), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n491_), .A2(new_n493_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n456_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n623_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT43), .ZN(new_n679_));
  AOI21_X1  g478(.A(KEYINPUT104), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT104), .ZN(new_n681_));
  NOR4_X1   g480(.A1(new_n494_), .A2(new_n681_), .A3(KEYINPUT43), .A4(new_n623_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n487_), .A2(new_n488_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT96), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n485_), .A2(KEYINPUT96), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n685_), .A2(new_n686_), .A3(new_n462_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n492_), .B1(new_n687_), .B2(new_n461_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n493_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n677_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n623_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n679_), .B1(new_n690_), .B2(new_n691_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n680_), .A2(new_n682_), .A3(new_n692_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n644_), .A2(new_n636_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n675_), .B1(new_n693_), .B2(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n690_), .A2(new_n679_), .A3(new_n691_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(new_n681_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n678_), .A2(KEYINPUT104), .A3(new_n679_), .ZN(new_n699_));
  OAI21_X1  g498(.A(KEYINPUT43), .B1(new_n494_), .B2(new_n623_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n698_), .A2(new_n699_), .A3(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n701_), .A2(KEYINPUT44), .A3(new_n694_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n696_), .A2(new_n335_), .A3(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(G29gat), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n494_), .A2(new_n530_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n645_), .A2(new_n617_), .ZN(new_n706_));
  XOR2_X1   g505(.A(new_n706_), .B(KEYINPUT105), .Z(new_n707_));
  AND2_X1   g506(.A1(new_n707_), .A2(new_n643_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n705_), .A2(new_n708_), .ZN(new_n709_));
  NOR3_X1   g508(.A1(new_n709_), .A2(G29gat), .A3(new_n336_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n674_), .B1(new_n704_), .B2(new_n711_), .ZN(new_n712_));
  AOI211_X1 g511(.A(KEYINPUT106), .B(new_n710_), .C1(new_n703_), .C2(G29gat), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1328gat));
  INV_X1    g513(.A(new_n709_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT107), .ZN(new_n716_));
  INV_X1    g515(.A(G36gat), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n656_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n715_), .A2(new_n716_), .A3(new_n719_), .ZN(new_n720_));
  OAI21_X1  g519(.A(KEYINPUT107), .B1(new_n709_), .B2(new_n718_), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n720_), .A2(KEYINPUT45), .A3(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(KEYINPUT45), .B1(new_n720_), .B2(new_n721_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n701_), .A2(KEYINPUT44), .A3(new_n694_), .ZN(new_n725_));
  AOI21_X1  g524(.A(KEYINPUT44), .B1(new_n701_), .B2(new_n694_), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n725_), .A2(new_n726_), .A3(new_n657_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n724_), .B1(new_n727_), .B2(new_n717_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT46), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n724_), .B(KEYINPUT46), .C1(new_n727_), .C2(new_n717_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(G1329gat));
  OAI211_X1 g531(.A(G43gat), .B(new_n390_), .C1(new_n395_), .C2(new_n396_), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n725_), .A2(new_n726_), .A3(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(G43gat), .B1(new_n715_), .B2(new_n666_), .ZN(new_n735_));
  OR3_X1    g534(.A1(new_n734_), .A2(KEYINPUT47), .A3(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(KEYINPUT47), .B1(new_n734_), .B2(new_n735_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(G1330gat));
  AOI21_X1  g537(.A(G50gat), .B1(new_n715_), .B2(new_n299_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n725_), .A2(new_n726_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n299_), .A2(G50gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n739_), .B1(new_n740_), .B2(new_n741_), .ZN(G1331gat));
  AND4_X1   g541(.A1(new_n647_), .A2(new_n636_), .A3(new_n530_), .A4(new_n596_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n743_), .A2(G57gat), .A3(new_n335_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT109), .ZN(new_n745_));
  NOR4_X1   g544(.A1(new_n494_), .A2(new_n529_), .A3(new_n643_), .A4(new_n637_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT108), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n747_), .A2(new_n336_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n745_), .B1(new_n748_), .B2(G57gat), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT110), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT110), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n745_), .B(new_n751_), .C1(G57gat), .C2(new_n748_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(G1332gat));
  INV_X1    g552(.A(G64gat), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n754_), .B1(new_n743_), .B2(new_n656_), .ZN(new_n755_));
  XOR2_X1   g554(.A(new_n755_), .B(KEYINPUT48), .Z(new_n756_));
  NAND2_X1  g555(.A1(new_n656_), .A2(new_n754_), .ZN(new_n757_));
  XOR2_X1   g556(.A(new_n757_), .B(KEYINPUT111), .Z(new_n758_));
  OAI21_X1  g557(.A(new_n756_), .B1(new_n747_), .B2(new_n758_), .ZN(G1333gat));
  NAND2_X1  g558(.A1(new_n743_), .A2(new_n666_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(G71gat), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT112), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT49), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT112), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n761_), .B(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT49), .ZN(new_n767_));
  OR3_X1    g566(.A1(new_n747_), .A2(G71gat), .A3(new_n461_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n764_), .A2(new_n767_), .A3(new_n768_), .ZN(G1334gat));
  AOI21_X1  g568(.A(new_n263_), .B1(new_n743_), .B2(new_n299_), .ZN(new_n770_));
  XOR2_X1   g569(.A(new_n770_), .B(KEYINPUT50), .Z(new_n771_));
  NAND2_X1  g570(.A1(new_n299_), .A2(new_n263_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n771_), .B1(new_n747_), .B2(new_n772_), .ZN(G1335gat));
  NOR3_X1   g572(.A1(new_n643_), .A2(new_n636_), .A3(new_n529_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n701_), .A2(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(G85gat), .B1(new_n775_), .B2(new_n336_), .ZN(new_n776_));
  NOR3_X1   g575(.A1(new_n494_), .A2(new_n529_), .A3(new_n643_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(new_n707_), .ZN(new_n778_));
  OR2_X1    g577(.A1(new_n336_), .A2(G85gat), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n776_), .B1(new_n778_), .B2(new_n779_), .ZN(G1336gat));
  OAI21_X1  g579(.A(G92gat), .B1(new_n775_), .B2(new_n657_), .ZN(new_n781_));
  OR2_X1    g580(.A1(new_n657_), .A2(G92gat), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n781_), .B1(new_n778_), .B2(new_n782_), .ZN(G1337gat));
  OAI21_X1  g582(.A(G99gat), .B1(new_n775_), .B2(new_n461_), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n390_), .B(new_n541_), .C1(new_n395_), .C2(new_n396_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n784_), .B1(new_n778_), .B2(new_n785_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g586(.A1(new_n777_), .A2(new_n291_), .A3(new_n299_), .A4(new_n707_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n701_), .A2(new_n299_), .A3(new_n774_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT52), .ZN(new_n790_));
  AND3_X1   g589(.A1(new_n789_), .A2(new_n790_), .A3(G106gat), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n789_), .B2(G106gat), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n788_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT53), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT53), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n795_), .B(new_n788_), .C1(new_n791_), .C2(new_n792_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(G1339gat));
  OAI21_X1  g596(.A(KEYINPUT55), .B1(new_n578_), .B2(new_n579_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(new_n580_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n578_), .A2(KEYINPUT55), .A3(new_n579_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n590_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n801_), .A2(KEYINPUT56), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT56), .ZN(new_n803_));
  AOI211_X1 g602(.A(new_n803_), .B(new_n590_), .C1(new_n799_), .C2(new_n800_), .ZN(new_n804_));
  OR2_X1    g603(.A1(new_n802_), .A2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n509_), .A2(new_n516_), .A3(new_n519_), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n525_), .B(new_n806_), .C1(new_n512_), .C2(new_n516_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n528_), .A2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n591_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n805_), .A2(KEYINPUT117), .A3(KEYINPUT58), .A4(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n810_), .B1(new_n802_), .B2(new_n804_), .ZN(new_n812_));
  XOR2_X1   g611(.A(KEYINPUT116), .B(KEYINPUT58), .Z(new_n813_));
  AOI21_X1  g612(.A(new_n623_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT117), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT58), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n815_), .B1(new_n812_), .B2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n811_), .A2(new_n814_), .A3(new_n817_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n530_), .A2(new_n809_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n799_), .A2(new_n800_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n588_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n803_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n801_), .A2(KEYINPUT114), .A3(KEYINPUT56), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n804_), .A2(KEYINPUT114), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n819_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT115), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(new_n593_), .B2(new_n808_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n592_), .A2(KEYINPUT115), .A3(new_n528_), .A4(new_n807_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n617_), .B1(new_n826_), .B2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n818_), .B1(new_n832_), .B2(KEYINPUT57), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT114), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n834_), .B1(new_n821_), .B2(new_n803_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n835_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n830_), .B1(new_n836_), .B2(new_n819_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT57), .ZN(new_n838_));
  NOR3_X1   g637(.A1(new_n837_), .A2(new_n838_), .A3(new_n617_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n645_), .B1(new_n833_), .B2(new_n839_), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n637_), .A2(new_n596_), .A3(new_n529_), .ZN(new_n841_));
  OR2_X1    g640(.A1(KEYINPUT113), .A2(KEYINPUT54), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  XOR2_X1   g642(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n844_));
  AOI21_X1  g643(.A(new_n843_), .B1(new_n841_), .B2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n840_), .A2(new_n845_), .ZN(new_n846_));
  NOR4_X1   g645(.A1(new_n656_), .A2(new_n336_), .A3(new_n457_), .A4(new_n299_), .ZN(new_n847_));
  XOR2_X1   g646(.A(new_n847_), .B(KEYINPUT118), .Z(new_n848_));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n848_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(KEYINPUT59), .ZN(new_n850_));
  OAI21_X1  g649(.A(G113gat), .B1(new_n850_), .B2(new_n530_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n846_), .A2(new_n848_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n852_), .A2(new_n314_), .A3(new_n529_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n853_), .ZN(G1340gat));
  OAI21_X1  g653(.A(G120gat), .B1(new_n850_), .B2(new_n643_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n312_), .B1(new_n643_), .B2(KEYINPUT60), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n852_), .B(new_n856_), .C1(KEYINPUT60), .C2(new_n312_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n857_), .ZN(G1341gat));
  OAI21_X1  g657(.A(new_n309_), .B1(new_n849_), .B2(new_n645_), .ZN(new_n859_));
  OR2_X1    g658(.A1(new_n859_), .A2(KEYINPUT119), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(KEYINPUT119), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n852_), .B(KEYINPUT59), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n645_), .A2(new_n309_), .ZN(new_n863_));
  AOI22_X1  g662(.A1(new_n860_), .A2(new_n861_), .B1(new_n862_), .B2(new_n863_), .ZN(G1342gat));
  OAI21_X1  g663(.A(G134gat), .B1(new_n850_), .B2(new_n623_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n852_), .A2(new_n307_), .A3(new_n617_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(G1343gat));
  NAND2_X1  g666(.A1(new_n846_), .A2(new_n461_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n657_), .A2(new_n335_), .A3(new_n299_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n529_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g671(.A1(new_n870_), .A2(new_n596_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(KEYINPUT120), .B(G148gat), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n873_), .B(new_n874_), .ZN(G1345gat));
  NAND2_X1  g674(.A1(new_n870_), .A2(new_n636_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(KEYINPUT61), .B(G155gat), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n876_), .B(new_n877_), .ZN(G1346gat));
  INV_X1    g677(.A(G162gat), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n870_), .A2(new_n879_), .A3(new_n617_), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n868_), .A2(new_n623_), .A3(new_n869_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n881_), .B2(new_n879_), .ZN(G1347gat));
  NAND4_X1  g681(.A1(new_n656_), .A2(new_n336_), .A3(new_n666_), .A4(new_n488_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n883_), .A2(new_n530_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n885_), .B1(new_n840_), .B2(new_n845_), .ZN(new_n886_));
  OAI21_X1  g685(.A(KEYINPUT121), .B1(new_n886_), .B2(new_n361_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT121), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n841_), .A2(new_n844_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n889_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n832_), .A2(KEYINPUT57), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n838_), .B1(new_n837_), .B2(new_n617_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n891_), .A2(new_n892_), .A3(new_n818_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n890_), .B1(new_n893_), .B2(new_n645_), .ZN(new_n894_));
  OAI211_X1 g693(.A(new_n888_), .B(G169gat), .C1(new_n894_), .C2(new_n885_), .ZN(new_n895_));
  AND3_X1   g694(.A1(new_n887_), .A2(KEYINPUT62), .A3(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT62), .ZN(new_n897_));
  OAI211_X1 g696(.A(KEYINPUT121), .B(new_n897_), .C1(new_n886_), .C2(new_n361_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(KEYINPUT22), .B(G169gat), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n886_), .A2(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n900_), .ZN(new_n901_));
  OAI21_X1  g700(.A(KEYINPUT122), .B1(new_n896_), .B2(new_n901_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n887_), .A2(KEYINPUT62), .A3(new_n895_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n904_));
  NAND4_X1  g703(.A1(new_n903_), .A2(new_n904_), .A3(new_n898_), .A4(new_n900_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n902_), .A2(new_n905_), .ZN(G1348gat));
  NOR2_X1   g705(.A1(new_n894_), .A2(new_n883_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(new_n596_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(KEYINPUT123), .B(G176gat), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n908_), .B(new_n909_), .ZN(G1349gat));
  NOR3_X1   g709(.A1(new_n894_), .A2(new_n645_), .A3(new_n883_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n409_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n912_), .B1(G183gat), .B2(new_n911_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(KEYINPUT124), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT124), .ZN(new_n915_));
  OAI211_X1 g714(.A(new_n912_), .B(new_n915_), .C1(G183gat), .C2(new_n911_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n914_), .A2(new_n916_), .ZN(G1350gat));
  NAND2_X1  g716(.A1(new_n413_), .A2(new_n414_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n907_), .A2(new_n918_), .A3(new_n617_), .ZN(new_n919_));
  NOR3_X1   g718(.A1(new_n894_), .A2(new_n623_), .A3(new_n883_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n919_), .B1(new_n920_), .B2(new_n337_), .ZN(G1351gat));
  NOR2_X1   g720(.A1(new_n894_), .A2(new_n666_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n488_), .A2(new_n335_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n656_), .A2(new_n923_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n924_), .ZN(new_n925_));
  NAND4_X1  g724(.A1(new_n922_), .A2(G197gat), .A3(new_n529_), .A4(new_n925_), .ZN(new_n926_));
  AND2_X1   g725(.A1(new_n926_), .A2(KEYINPUT125), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n926_), .A2(KEYINPUT125), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n868_), .A2(new_n924_), .ZN(new_n929_));
  AOI21_X1  g728(.A(G197gat), .B1(new_n929_), .B2(new_n529_), .ZN(new_n930_));
  NOR3_X1   g729(.A1(new_n927_), .A2(new_n928_), .A3(new_n930_), .ZN(G1352gat));
  NAND2_X1  g730(.A1(new_n929_), .A2(new_n596_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n217_), .A2(KEYINPUT126), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n932_), .B(new_n933_), .ZN(G1353gat));
  XNOR2_X1  g733(.A(KEYINPUT63), .B(G211gat), .ZN(new_n935_));
  NAND4_X1  g734(.A1(new_n922_), .A2(new_n636_), .A3(new_n925_), .A4(new_n935_), .ZN(new_n936_));
  NOR3_X1   g735(.A1(new_n868_), .A2(new_n645_), .A3(new_n924_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n936_), .B1(new_n937_), .B2(new_n938_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n939_), .A2(KEYINPUT127), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT127), .ZN(new_n941_));
  OAI211_X1 g740(.A(new_n941_), .B(new_n936_), .C1(new_n937_), .C2(new_n938_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n940_), .A2(new_n942_), .ZN(G1354gat));
  NAND3_X1  g742(.A1(new_n929_), .A2(new_n226_), .A3(new_n617_), .ZN(new_n944_));
  NOR3_X1   g743(.A1(new_n868_), .A2(new_n623_), .A3(new_n924_), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n944_), .B1(new_n945_), .B2(new_n226_), .ZN(G1355gat));
endmodule


