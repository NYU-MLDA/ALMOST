//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 0 0 1 0 0 1 0 1 0 1 0 1 1 1 0 1 0 0 1 1 1 0 0 1 0 1 0 1 1 1 0 1 1 0 1 0 0 1 0 1 1 0 1 1 1 0 1 0 1 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n734_, new_n735_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n769_, new_n770_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n864_, new_n865_, new_n867_, new_n868_, new_n869_,
    new_n871_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n904_, new_n905_, new_n906_,
    new_n907_, new_n909_, new_n910_, new_n911_, new_n912_, new_n914_,
    new_n915_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_, new_n925_;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT71), .ZN(new_n203_));
  AOI21_X1  g002(.A(KEYINPUT65), .B1(G85gat), .B2(G92gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT66), .ZN(new_n205_));
  OR2_X1    g004(.A1(new_n205_), .A2(KEYINPUT9), .ZN(new_n206_));
  NOR2_X1   g005(.A1(G85gat), .A2(G92gat), .ZN(new_n207_));
  AND2_X1   g006(.A1(G85gat), .A2(G92gat), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n207_), .B1(new_n208_), .B2(KEYINPUT66), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n205_), .A2(KEYINPUT9), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n206_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT6), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT67), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  XOR2_X1   g014(.A(KEYINPUT10), .B(G99gat), .Z(new_n216_));
  INV_X1    g015(.A(G106gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n211_), .A2(new_n215_), .A3(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n208_), .A2(new_n207_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT8), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(G99gat), .A2(G106gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n223_), .B(KEYINPUT7), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n222_), .B1(new_n215_), .B2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(new_n213_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(new_n220_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT68), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT68), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n227_), .A2(new_n230_), .A3(new_n220_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n229_), .A2(KEYINPUT8), .A3(new_n231_), .ZN(new_n232_));
  AND3_X1   g031(.A1(new_n226_), .A2(KEYINPUT70), .A3(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(KEYINPUT70), .B1(new_n226_), .B2(new_n232_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n219_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G57gat), .B(G64gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT69), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT11), .ZN(new_n238_));
  XOR2_X1   g037(.A(G71gat), .B(G78gat), .Z(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n238_), .A2(new_n240_), .ZN(new_n241_));
  XOR2_X1   g040(.A(new_n237_), .B(KEYINPUT11), .Z(new_n242_));
  OAI21_X1  g041(.A(new_n241_), .B1(new_n242_), .B2(new_n240_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n235_), .A2(KEYINPUT12), .A3(new_n243_), .ZN(new_n244_));
  AND3_X1   g043(.A1(new_n229_), .A2(KEYINPUT8), .A3(new_n231_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n219_), .B1(new_n245_), .B2(new_n225_), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT12), .B1(new_n246_), .B2(new_n243_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n243_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G230gat), .A2(G233gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT64), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n244_), .A2(new_n249_), .A3(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n251_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n248_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n246_), .A2(new_n243_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n253_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT5), .B(G176gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(G204gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G120gat), .B(G148gat), .ZN(new_n259_));
  XOR2_X1   g058(.A(new_n258_), .B(new_n259_), .Z(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  AND3_X1   g060(.A1(new_n252_), .A2(new_n256_), .A3(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n261_), .B1(new_n252_), .B2(new_n256_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n203_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n252_), .A2(new_n256_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(new_n260_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n252_), .A2(new_n256_), .A3(new_n261_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n266_), .A2(KEYINPUT71), .A3(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n264_), .A2(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n202_), .B1(new_n269_), .B2(KEYINPUT13), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT13), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n264_), .A2(new_n268_), .A3(KEYINPUT72), .A4(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT73), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n274_), .B1(new_n269_), .B2(KEYINPUT13), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n269_), .A2(new_n274_), .A3(KEYINPUT13), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n273_), .B1(new_n275_), .B2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT74), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT85), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G169gat), .A2(G176gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT24), .ZN(new_n283_));
  NOR2_X1   g082(.A1(G169gat), .A2(G176gat), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n281_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(G169gat), .ZN(new_n286_));
  INV_X1    g085(.A(G176gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n288_), .A2(KEYINPUT85), .A3(KEYINPUT24), .A4(new_n282_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n285_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G183gat), .A2(G190gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT23), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT23), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n293_), .A2(G183gat), .A3(G190gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT24), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n284_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(KEYINPUT25), .B(G183gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(KEYINPUT84), .A2(G190gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT26), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT26), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n301_), .A2(KEYINPUT84), .A3(G190gat), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n298_), .A2(new_n300_), .A3(new_n302_), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n290_), .A2(new_n295_), .A3(new_n297_), .A4(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n287_), .A2(KEYINPUT86), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT86), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(G176gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(KEYINPUT22), .B(G169gat), .ZN(new_n309_));
  AOI22_X1  g108(.A1(new_n308_), .A2(new_n309_), .B1(G169gat), .B2(G176gat), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n293_), .B1(G183gat), .B2(G190gat), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT87), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n294_), .A2(new_n312_), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n293_), .A2(KEYINPUT87), .A3(G183gat), .A4(G190gat), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n311_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(G183gat), .A2(G190gat), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n310_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n304_), .A2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT30), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G127gat), .B(G134gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G113gat), .B(G120gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n319_), .B(new_n323_), .ZN(new_n324_));
  XOR2_X1   g123(.A(G15gat), .B(G43gat), .Z(new_n325_));
  NAND2_X1  g124(.A1(G227gat), .A2(G233gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n324_), .B(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G71gat), .B(G99gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT88), .B(KEYINPUT31), .ZN(new_n330_));
  XOR2_X1   g129(.A(new_n329_), .B(new_n330_), .Z(new_n331_));
  OR2_X1    g130(.A1(new_n328_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n328_), .A2(new_n331_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(G155gat), .A2(G162gat), .ZN(new_n336_));
  AND2_X1   g135(.A1(G155gat), .A2(G162gat), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT1), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n336_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT89), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n340_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G155gat), .A2(G162gat), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n342_), .A2(KEYINPUT89), .A3(KEYINPUT1), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n339_), .A2(new_n341_), .A3(new_n343_), .ZN(new_n344_));
  XOR2_X1   g143(.A(G141gat), .B(G148gat), .Z(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT3), .ZN(new_n347_));
  INV_X1    g146(.A(G141gat), .ZN(new_n348_));
  INV_X1    g147(.A(G148gat), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n347_), .A2(new_n348_), .A3(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G141gat), .A2(G148gat), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT2), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n350_), .A2(new_n353_), .A3(new_n354_), .A4(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n336_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n356_), .A2(new_n342_), .A3(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n346_), .A2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(new_n322_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(KEYINPUT4), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G225gat), .A2(G233gat), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  AND2_X1   g162(.A1(new_n356_), .A2(new_n342_), .ZN(new_n364_));
  AOI22_X1  g163(.A1(new_n364_), .A2(new_n357_), .B1(new_n345_), .B2(new_n344_), .ZN(new_n365_));
  OR3_X1    g164(.A1(new_n365_), .A2(KEYINPUT4), .A3(new_n322_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n361_), .A2(new_n363_), .A3(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n360_), .A2(new_n362_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G1gat), .B(G29gat), .ZN(new_n370_));
  INV_X1    g169(.A(G85gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(KEYINPUT0), .B(G57gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n372_), .B(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n369_), .B(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n315_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(KEYINPUT26), .B(G190gat), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n296_), .B1(G169gat), .B2(G176gat), .ZN(new_n379_));
  AOI22_X1  g178(.A1(new_n298_), .A2(new_n378_), .B1(new_n379_), .B2(new_n288_), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n377_), .A2(KEYINPUT95), .A3(new_n297_), .A4(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT95), .ZN(new_n382_));
  NOR2_X1   g181(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n383_));
  AND2_X1   g182(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n384_));
  AND2_X1   g183(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n385_));
  NOR2_X1   g184(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n386_));
  OAI22_X1  g185(.A1(new_n383_), .A2(new_n384_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n379_), .A2(new_n288_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n387_), .A2(new_n388_), .A3(new_n297_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n382_), .B1(new_n389_), .B2(new_n315_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n381_), .A2(new_n390_), .ZN(new_n391_));
  AND2_X1   g190(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n392_));
  NOR2_X1   g191(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT86), .B(G176gat), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n282_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT96), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n316_), .B1(new_n292_), .B2(new_n294_), .ZN(new_n398_));
  NOR3_X1   g197(.A1(new_n396_), .A2(new_n397_), .A3(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n398_), .ZN(new_n400_));
  AOI21_X1  g199(.A(KEYINPUT96), .B1(new_n310_), .B2(new_n400_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n391_), .A2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G197gat), .B(G204gat), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT21), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(G197gat), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n407_), .A2(G204gat), .ZN(new_n408_));
  INV_X1    g207(.A(G204gat), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n409_), .A2(G197gat), .ZN(new_n410_));
  OAI21_X1  g209(.A(KEYINPUT21), .B1(new_n408_), .B2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G211gat), .B(G218gat), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n406_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n413_));
  XOR2_X1   g212(.A(G211gat), .B(G218gat), .Z(new_n414_));
  OAI211_X1 g213(.A(new_n414_), .B(KEYINPUT21), .C1(new_n408_), .C2(new_n410_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(KEYINPUT97), .B1(new_n403_), .B2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT97), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n413_), .A2(new_n415_), .ZN(new_n419_));
  AOI211_X1 g218(.A(new_n418_), .B(new_n419_), .C1(new_n391_), .C2(new_n402_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n419_), .A2(new_n317_), .A3(new_n304_), .ZN(new_n421_));
  AOI21_X1  g220(.A(KEYINPUT94), .B1(new_n421_), .B2(KEYINPUT20), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n421_), .A2(KEYINPUT94), .A3(KEYINPUT20), .ZN(new_n423_));
  OAI22_X1  g222(.A1(new_n417_), .A2(new_n420_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G226gat), .A2(G233gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n425_), .B(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n424_), .A2(new_n428_), .ZN(new_n429_));
  XOR2_X1   g228(.A(G64gat), .B(G92gat), .Z(new_n430_));
  XNOR2_X1  g229(.A(G8gat), .B(G36gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n430_), .B(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n432_), .B(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT32), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n391_), .A2(new_n402_), .A3(new_n419_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n318_), .A2(new_n416_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n436_), .A2(KEYINPUT20), .A3(new_n427_), .A4(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n429_), .A2(new_n435_), .A3(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT20), .B1(new_n318_), .B2(new_n416_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT94), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n421_), .A2(KEYINPUT94), .A3(KEYINPUT20), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n444_), .B(new_n427_), .C1(new_n417_), .C2(new_n420_), .ZN(new_n445_));
  OAI22_X1  g244(.A1(new_n389_), .A2(new_n315_), .B1(new_n396_), .B2(new_n398_), .ZN(new_n446_));
  OAI21_X1  g245(.A(KEYINPUT20), .B1(new_n446_), .B2(new_n416_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT100), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT100), .ZN(new_n449_));
  OAI211_X1 g248(.A(new_n449_), .B(KEYINPUT20), .C1(new_n446_), .C2(new_n416_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n448_), .A2(new_n437_), .A3(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(new_n428_), .ZN(new_n452_));
  AND2_X1   g251(.A1(new_n445_), .A2(new_n452_), .ZN(new_n453_));
  OAI211_X1 g252(.A(new_n376_), .B(new_n439_), .C1(new_n435_), .C2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n367_), .A2(new_n368_), .A3(new_n374_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(KEYINPUT33), .ZN(new_n456_));
  AND3_X1   g255(.A1(new_n361_), .A2(new_n362_), .A3(new_n366_), .ZN(new_n457_));
  OR2_X1    g256(.A1(new_n457_), .A2(KEYINPUT99), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n374_), .B1(new_n360_), .B2(new_n363_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(KEYINPUT99), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n458_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n397_), .B1(new_n396_), .B2(new_n398_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n310_), .A2(new_n400_), .A3(KEYINPUT96), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n464_), .B1(new_n390_), .B2(new_n381_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n418_), .B1(new_n465_), .B2(new_n419_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n403_), .A2(KEYINPUT97), .A3(new_n416_), .ZN(new_n467_));
  AOI22_X1  g266(.A1(new_n466_), .A2(new_n467_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n468_));
  OAI211_X1 g267(.A(new_n434_), .B(new_n438_), .C1(new_n468_), .C2(new_n427_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n434_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n466_), .A2(new_n467_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n427_), .B1(new_n471_), .B2(new_n444_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n438_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n470_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n456_), .A2(new_n461_), .A3(new_n469_), .A4(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n454_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT29), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n477_), .B1(new_n346_), .B2(new_n358_), .ZN(new_n478_));
  AND2_X1   g277(.A1(G228gat), .A2(G233gat), .ZN(new_n479_));
  NOR3_X1   g278(.A1(new_n478_), .A2(new_n419_), .A3(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  XOR2_X1   g280(.A(KEYINPUT91), .B(KEYINPUT29), .Z(new_n482_));
  OAI21_X1  g281(.A(new_n416_), .B1(new_n365_), .B2(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(KEYINPUT92), .B1(new_n483_), .B2(new_n479_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n482_), .B1(new_n346_), .B2(new_n358_), .ZN(new_n485_));
  OAI211_X1 g284(.A(KEYINPUT92), .B(new_n479_), .C1(new_n485_), .C2(new_n419_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n481_), .B1(new_n484_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(G22gat), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n479_), .B1(new_n485_), .B2(new_n419_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT92), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(new_n486_), .ZN(new_n493_));
  INV_X1    g292(.A(G22gat), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n493_), .A2(new_n494_), .A3(new_n481_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n489_), .A2(G50gat), .A3(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(G50gat), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n494_), .B1(new_n493_), .B2(new_n481_), .ZN(new_n498_));
  AOI211_X1 g297(.A(G22gat), .B(new_n480_), .C1(new_n492_), .C2(new_n486_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n497_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n496_), .A2(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n359_), .A2(KEYINPUT29), .ZN(new_n502_));
  XNOR2_X1  g301(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n502_), .B(new_n503_), .ZN(new_n504_));
  XOR2_X1   g303(.A(G78gat), .B(G106gat), .Z(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n501_), .A2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n496_), .A2(new_n500_), .A3(new_n506_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n476_), .A2(new_n510_), .ZN(new_n511_));
  AOI211_X1 g310(.A(new_n470_), .B(new_n473_), .C1(new_n424_), .C2(new_n428_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT27), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n434_), .B1(new_n445_), .B2(new_n452_), .ZN(new_n514_));
  NOR3_X1   g313(.A1(new_n512_), .A2(new_n513_), .A3(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(KEYINPUT27), .B1(new_n474_), .B2(new_n469_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  AND3_X1   g316(.A1(new_n496_), .A2(new_n500_), .A3(new_n506_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n506_), .B1(new_n496_), .B2(new_n500_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n517_), .A2(new_n375_), .A3(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n335_), .B1(new_n511_), .B2(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n332_), .A2(new_n375_), .A3(new_n333_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n434_), .B1(new_n429_), .B2(new_n438_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n513_), .B1(new_n525_), .B2(new_n512_), .ZN(new_n526_));
  OAI211_X1 g325(.A(KEYINPUT27), .B(new_n469_), .C1(new_n453_), .C2(new_n434_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NOR3_X1   g327(.A1(new_n528_), .A2(new_n520_), .A3(KEYINPUT101), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT101), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n530_), .B1(new_n517_), .B2(new_n510_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n524_), .B1(new_n529_), .B2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(KEYINPUT102), .ZN(new_n533_));
  OAI21_X1  g332(.A(KEYINPUT101), .B1(new_n528_), .B2(new_n520_), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n510_), .A2(new_n530_), .A3(new_n526_), .A4(new_n527_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT102), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n536_), .A2(new_n537_), .A3(new_n524_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n522_), .B1(new_n533_), .B2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G15gat), .B(G22gat), .ZN(new_n540_));
  INV_X1    g339(.A(G1gat), .ZN(new_n541_));
  INV_X1    g340(.A(G8gat), .ZN(new_n542_));
  OAI21_X1  g341(.A(KEYINPUT14), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n540_), .A2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G1gat), .B(G8gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G29gat), .B(G36gat), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G43gat), .B(G50gat), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n549_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(new_n547_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n546_), .A2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(KEYINPUT76), .B(KEYINPUT15), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n553_), .B(new_n555_), .Z(new_n556_));
  AOI21_X1  g355(.A(new_n554_), .B1(new_n556_), .B2(new_n546_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G229gat), .A2(G233gat), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n546_), .B(new_n553_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n560_), .A2(G229gat), .A3(G233gat), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n559_), .B1(KEYINPUT81), .B2(new_n561_), .ZN(new_n562_));
  AND2_X1   g361(.A1(new_n561_), .A2(KEYINPUT81), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G113gat), .B(G141gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G169gat), .B(G197gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  OR3_X1    g365(.A1(new_n562_), .A2(new_n563_), .A3(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n566_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT82), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n567_), .A2(KEYINPUT82), .A3(new_n568_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT83), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n571_), .A2(KEYINPUT83), .A3(new_n572_), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n539_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT37), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G190gat), .B(G218gat), .ZN(new_n580_));
  INV_X1    g379(.A(G162gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(KEYINPUT77), .B(G134gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT36), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(KEYINPUT75), .B(KEYINPUT34), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G232gat), .A2(G233gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT35), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n553_), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n219_), .B(new_n593_), .C1(new_n245_), .C2(new_n225_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n219_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT70), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n596_), .B1(new_n245_), .B2(new_n225_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n226_), .A2(KEYINPUT70), .A3(new_n232_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n595_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n556_), .ZN(new_n600_));
  OAI211_X1 g399(.A(new_n592_), .B(new_n594_), .C1(new_n599_), .C2(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n590_), .A2(new_n591_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n235_), .A2(new_n556_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n602_), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n604_), .A2(new_n605_), .A3(new_n592_), .A4(new_n594_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n585_), .B1(new_n603_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n584_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n587_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n603_), .A2(new_n606_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(KEYINPUT78), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n609_), .A2(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n609_), .A2(new_n612_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n579_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(G231gat), .A2(G233gat), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n546_), .B(new_n616_), .Z(new_n617_));
  XNOR2_X1  g416(.A(new_n243_), .B(new_n617_), .ZN(new_n618_));
  XOR2_X1   g417(.A(G183gat), .B(G211gat), .Z(new_n619_));
  XNOR2_X1  g418(.A(G127gat), .B(G155gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  OR2_X1    g422(.A1(new_n623_), .A2(KEYINPUT17), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(KEYINPUT17), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n618_), .A2(new_n624_), .A3(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT80), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(KEYINPUT80), .B1(new_n618_), .B2(new_n625_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n628_), .B1(new_n629_), .B2(new_n626_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n609_), .A2(new_n612_), .ZN(new_n631_));
  OAI211_X1 g430(.A(new_n611_), .B(new_n587_), .C1(new_n607_), .C2(new_n608_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n631_), .A2(KEYINPUT37), .A3(new_n632_), .ZN(new_n633_));
  AND3_X1   g432(.A1(new_n615_), .A2(new_n630_), .A3(new_n633_), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n280_), .A2(new_n578_), .A3(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n635_), .B1(KEYINPUT103), .B2(KEYINPUT38), .ZN(new_n636_));
  NOR3_X1   g435(.A1(new_n636_), .A2(G1gat), .A3(new_n375_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(KEYINPUT103), .A2(KEYINPUT38), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n637_), .B(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n573_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n278_), .A2(new_n640_), .A3(new_n630_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT104), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n642_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n613_), .A2(new_n614_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n539_), .A2(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n643_), .A2(new_n644_), .A3(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(G1gat), .B1(new_n647_), .B2(new_n375_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT105), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n639_), .A2(new_n649_), .ZN(G1324gat));
  OAI21_X1  g449(.A(G8gat), .B1(new_n647_), .B2(new_n517_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT106), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n652_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n653_), .A2(KEYINPUT39), .A3(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n635_), .A2(new_n542_), .A3(new_n528_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT39), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n651_), .A2(new_n652_), .A3(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n655_), .A2(new_n656_), .A3(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT40), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n655_), .A2(KEYINPUT40), .A3(new_n656_), .A4(new_n658_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1325gat));
  OAI21_X1  g462(.A(G15gat), .B1(new_n647_), .B2(new_n334_), .ZN(new_n664_));
  XOR2_X1   g463(.A(new_n664_), .B(KEYINPUT41), .Z(new_n665_));
  INV_X1    g464(.A(G15gat), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n635_), .A2(new_n666_), .A3(new_n335_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(G1326gat));
  OAI21_X1  g467(.A(G22gat), .B1(new_n647_), .B2(new_n510_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT42), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n635_), .A2(new_n494_), .A3(new_n520_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(G1327gat));
  INV_X1    g471(.A(KEYINPUT108), .ZN(new_n673_));
  INV_X1    g472(.A(new_n630_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n278_), .A2(new_n640_), .A3(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n615_), .A2(new_n633_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  OAI21_X1  g476(.A(KEYINPUT43), .B1(new_n539_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n521_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n520_), .B1(new_n454_), .B2(new_n475_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n334_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n537_), .B1(new_n536_), .B2(new_n524_), .ZN(new_n682_));
  AOI211_X1 g481(.A(KEYINPUT102), .B(new_n523_), .C1(new_n534_), .C2(new_n535_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n681_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT43), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n684_), .A2(new_n685_), .A3(new_n676_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n675_), .B1(new_n678_), .B2(new_n686_), .ZN(new_n687_));
  XOR2_X1   g486(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n688_));
  OAI21_X1  g487(.A(new_n673_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n675_), .ZN(new_n690_));
  AND3_X1   g489(.A1(new_n684_), .A2(new_n685_), .A3(new_n676_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n685_), .B1(new_n684_), .B2(new_n676_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n690_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n688_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n693_), .A2(KEYINPUT108), .A3(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n687_), .A2(KEYINPUT44), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n689_), .A2(new_n695_), .A3(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(G29gat), .B1(new_n697_), .B2(new_n375_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n645_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n699_), .A2(new_n630_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n578_), .A2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(new_n278_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n375_), .A2(G29gat), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT109), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n698_), .B1(new_n702_), .B2(new_n704_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT110), .ZN(G1328gat));
  NOR3_X1   g505(.A1(new_n687_), .A2(new_n673_), .A3(new_n688_), .ZN(new_n707_));
  AOI21_X1  g506(.A(KEYINPUT108), .B1(new_n693_), .B2(new_n694_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n709_), .A2(KEYINPUT111), .A3(new_n528_), .A4(new_n696_), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n689_), .A2(new_n695_), .A3(new_n528_), .A4(new_n696_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT111), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n710_), .A2(G36gat), .A3(new_n713_), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n702_), .A2(G36gat), .A3(new_n517_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT45), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n715_), .B(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n714_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT46), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n714_), .A2(KEYINPUT46), .A3(new_n717_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1329gat));
  INV_X1    g521(.A(G43gat), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n723_), .B1(new_n702_), .B2(new_n334_), .ZN(new_n724_));
  AND4_X1   g523(.A1(G43gat), .A2(new_n689_), .A3(new_n696_), .A4(new_n695_), .ZN(new_n725_));
  AOI21_X1  g524(.A(KEYINPUT112), .B1(new_n725_), .B2(new_n335_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT112), .ZN(new_n727_));
  NOR4_X1   g526(.A1(new_n697_), .A2(new_n727_), .A3(new_n723_), .A4(new_n334_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n724_), .B1(new_n726_), .B2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(KEYINPUT47), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT47), .ZN(new_n731_));
  OAI211_X1 g530(.A(new_n731_), .B(new_n724_), .C1(new_n726_), .C2(new_n728_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n730_), .A2(new_n732_), .ZN(G1330gat));
  OAI21_X1  g532(.A(G50gat), .B1(new_n697_), .B2(new_n510_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n701_), .A2(new_n497_), .A3(new_n278_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n734_), .B1(new_n510_), .B2(new_n735_), .ZN(G1331gat));
  NOR2_X1   g535(.A1(new_n539_), .A2(new_n640_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n269_), .A2(KEYINPUT13), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(KEYINPUT73), .ZN(new_n739_));
  AOI22_X1  g538(.A1(new_n739_), .A2(new_n276_), .B1(new_n270_), .B2(new_n272_), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n737_), .A2(new_n740_), .A3(new_n634_), .ZN(new_n741_));
  AOI21_X1  g540(.A(G57gat), .B1(new_n741_), .B2(new_n376_), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n279_), .A2(new_n646_), .A3(new_n630_), .A4(new_n577_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n743_), .A2(new_n375_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n742_), .B1(new_n744_), .B2(G57gat), .ZN(G1332gat));
  OAI21_X1  g544(.A(G64gat), .B1(new_n743_), .B2(new_n517_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT48), .ZN(new_n747_));
  INV_X1    g546(.A(G64gat), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n741_), .A2(new_n748_), .A3(new_n528_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(G1333gat));
  OAI21_X1  g549(.A(G71gat), .B1(new_n743_), .B2(new_n334_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT49), .ZN(new_n752_));
  INV_X1    g551(.A(G71gat), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n741_), .A2(new_n753_), .A3(new_n335_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n752_), .A2(new_n754_), .ZN(G1334gat));
  OAI21_X1  g554(.A(G78gat), .B1(new_n743_), .B2(new_n510_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT50), .ZN(new_n757_));
  INV_X1    g556(.A(G78gat), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n741_), .A2(new_n758_), .A3(new_n520_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(G1335gat));
  NOR2_X1   g559(.A1(new_n278_), .A2(new_n630_), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n573_), .B(new_n761_), .C1(new_n691_), .C2(new_n692_), .ZN(new_n762_));
  NOR3_X1   g561(.A1(new_n762_), .A2(new_n371_), .A3(new_n375_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n279_), .A2(new_n700_), .A3(new_n737_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT113), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n764_), .B(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(new_n376_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n763_), .B1(new_n767_), .B2(new_n371_), .ZN(G1336gat));
  AOI21_X1  g567(.A(G92gat), .B1(new_n766_), .B2(new_n528_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n762_), .A2(new_n517_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(G92gat), .B2(new_n770_), .ZN(G1337gat));
  NAND3_X1  g570(.A1(new_n766_), .A2(new_n216_), .A3(new_n335_), .ZN(new_n772_));
  OAI21_X1  g571(.A(G99gat), .B1(new_n762_), .B2(new_n334_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT51), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n772_), .B(new_n773_), .C1(KEYINPUT114), .C2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(KEYINPUT114), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n775_), .B(new_n776_), .ZN(G1338gat));
  NAND3_X1  g576(.A1(new_n766_), .A2(new_n217_), .A3(new_n520_), .ZN(new_n778_));
  OAI21_X1  g577(.A(G106gat), .B1(new_n762_), .B2(new_n510_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT52), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g581(.A(G113gat), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n251_), .B1(new_n244_), .B2(new_n249_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n252_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n244_), .A2(new_n249_), .A3(KEYINPUT55), .A4(new_n251_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n260_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n262_), .B1(new_n789_), .B2(KEYINPUT56), .ZN(new_n790_));
  AOI211_X1 g589(.A(new_n558_), .B(new_n554_), .C1(new_n556_), .C2(new_n546_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n566_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n792_), .B1(new_n560_), .B2(new_n558_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT118), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n567_), .B1(new_n791_), .B2(new_n794_), .ZN(new_n795_));
  XOR2_X1   g594(.A(new_n795_), .B(KEYINPUT119), .Z(new_n796_));
  INV_X1    g595(.A(KEYINPUT56), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n788_), .A2(new_n797_), .A3(new_n260_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n790_), .A2(new_n796_), .A3(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT58), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n790_), .A2(new_n796_), .A3(KEYINPUT58), .A4(new_n798_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n801_), .A2(new_n676_), .A3(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT121), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n801_), .A2(new_n676_), .A3(KEYINPUT121), .A4(new_n802_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n789_), .A2(KEYINPUT56), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n807_), .A2(new_n640_), .A3(new_n267_), .A4(new_n798_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n796_), .A2(new_n269_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n699_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT120), .ZN(new_n812_));
  AOI21_X1  g611(.A(KEYINPUT57), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n645_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT57), .ZN(new_n815_));
  NOR3_X1   g614(.A1(new_n814_), .A2(KEYINPUT120), .A3(new_n815_), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n805_), .B(new_n806_), .C1(new_n813_), .C2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n674_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n278_), .A2(new_n634_), .A3(new_n577_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n819_), .B1(new_n820_), .B2(KEYINPUT116), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT117), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n615_), .A2(new_n577_), .A3(new_n630_), .A4(new_n633_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n740_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT116), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n822_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  NOR4_X1   g625(.A1(new_n740_), .A2(new_n823_), .A3(KEYINPUT116), .A4(KEYINPUT117), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n821_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(KEYINPUT117), .B1(new_n820_), .B2(KEYINPUT116), .ZN(new_n829_));
  INV_X1    g628(.A(new_n819_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n830_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n824_), .A2(new_n825_), .A3(new_n822_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n829_), .A2(new_n831_), .A3(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n818_), .A2(new_n828_), .A3(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n536_), .A2(new_n376_), .A3(new_n335_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n783_), .B1(new_n837_), .B2(new_n573_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(KEYINPUT122), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n837_), .A2(KEYINPUT59), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n803_), .B1(new_n813_), .B2(new_n816_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n674_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n828_), .A2(new_n833_), .A3(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT59), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n843_), .A2(new_n844_), .A3(new_n836_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n840_), .A2(new_n845_), .ZN(new_n846_));
  NOR3_X1   g645(.A1(new_n846_), .A2(new_n783_), .A3(new_n577_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n839_), .A2(new_n847_), .ZN(G1340gat));
  NAND3_X1  g647(.A1(new_n840_), .A2(new_n279_), .A3(new_n845_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(KEYINPUT123), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT123), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n840_), .A2(new_n851_), .A3(new_n279_), .A4(new_n845_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n850_), .A2(G120gat), .A3(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n834_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n854_), .A2(new_n835_), .ZN(new_n855_));
  INV_X1    g654(.A(G120gat), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n856_), .B1(new_n278_), .B2(KEYINPUT60), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n855_), .B(new_n857_), .C1(KEYINPUT60), .C2(new_n856_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n853_), .A2(new_n858_), .ZN(G1341gat));
  AOI21_X1  g658(.A(G127gat), .B1(new_n855_), .B2(new_n630_), .ZN(new_n860_));
  INV_X1    g659(.A(G127gat), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n846_), .A2(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n860_), .B1(new_n862_), .B2(new_n630_), .ZN(G1342gat));
  AOI21_X1  g662(.A(G134gat), .B1(new_n855_), .B2(new_n645_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n846_), .A2(new_n677_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n864_), .B1(new_n865_), .B2(G134gat), .ZN(G1343gat));
  NOR2_X1   g665(.A1(new_n528_), .A2(new_n375_), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n834_), .A2(new_n520_), .A3(new_n334_), .A4(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n868_), .A2(new_n573_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(new_n348_), .ZN(G1344gat));
  NOR2_X1   g669(.A1(new_n868_), .A2(new_n280_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(new_n349_), .ZN(G1345gat));
  AND3_X1   g671(.A1(new_n834_), .A2(new_n520_), .A3(new_n334_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT124), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n873_), .A2(new_n874_), .A3(new_n630_), .A4(new_n867_), .ZN(new_n875_));
  OAI21_X1  g674(.A(KEYINPUT124), .B1(new_n868_), .B2(new_n674_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(KEYINPUT61), .B(G155gat), .ZN(new_n877_));
  AND3_X1   g676(.A1(new_n875_), .A2(new_n876_), .A3(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n877_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1346gat));
  NAND4_X1  g679(.A1(new_n873_), .A2(new_n581_), .A3(new_n645_), .A4(new_n867_), .ZN(new_n881_));
  OAI21_X1  g680(.A(G162gat), .B1(new_n868_), .B2(new_n677_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(KEYINPUT125), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT125), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n881_), .A2(new_n885_), .A3(new_n882_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n884_), .A2(new_n886_), .ZN(G1347gat));
  NOR3_X1   g686(.A1(new_n523_), .A2(new_n520_), .A3(new_n517_), .ZN(new_n888_));
  AND2_X1   g687(.A1(new_n843_), .A2(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n286_), .B1(new_n889_), .B2(new_n640_), .ZN(new_n890_));
  OR2_X1    g689(.A1(new_n890_), .A2(KEYINPUT62), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n889_), .A2(new_n309_), .A3(new_n640_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n890_), .A2(KEYINPUT62), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n891_), .A2(new_n892_), .A3(new_n893_), .ZN(G1348gat));
  AOI21_X1  g693(.A(new_n395_), .B1(new_n889_), .B2(new_n740_), .ZN(new_n895_));
  NOR3_X1   g694(.A1(new_n854_), .A2(new_n287_), .A3(new_n280_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n895_), .B1(new_n888_), .B2(new_n896_), .ZN(G1349gat));
  NAND2_X1  g696(.A1(new_n828_), .A2(new_n833_), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n898_), .A2(new_n888_), .ZN(new_n899_));
  AOI21_X1  g698(.A(G183gat), .B1(new_n899_), .B2(new_n630_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n843_), .A2(new_n888_), .ZN(new_n901_));
  NOR3_X1   g700(.A1(new_n901_), .A2(new_n298_), .A3(new_n674_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n900_), .A2(new_n902_), .ZN(G1350gat));
  NAND3_X1  g702(.A1(new_n889_), .A2(new_n645_), .A3(new_n378_), .ZN(new_n904_));
  OAI21_X1  g703(.A(G190gat), .B1(new_n901_), .B2(new_n677_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT126), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n906_), .B(new_n907_), .ZN(G1351gat));
  AND4_X1   g707(.A1(new_n375_), .A2(new_n834_), .A3(new_n520_), .A4(new_n334_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(new_n528_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n407_), .B1(new_n910_), .B2(new_n573_), .ZN(new_n911_));
  NAND4_X1  g710(.A1(new_n909_), .A2(G197gat), .A3(new_n528_), .A4(new_n640_), .ZN(new_n912_));
  AND2_X1   g711(.A1(new_n911_), .A2(new_n912_), .ZN(G1352gat));
  OAI211_X1 g712(.A(KEYINPUT127), .B(G204gat), .C1(new_n910_), .C2(new_n280_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n915_));
  NAND4_X1  g714(.A1(new_n909_), .A2(new_n528_), .A3(new_n279_), .A4(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n914_), .A2(new_n916_), .ZN(G1353gat));
  NOR2_X1   g716(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n918_), .B1(new_n910_), .B2(new_n674_), .ZN(new_n919_));
  XOR2_X1   g718(.A(KEYINPUT63), .B(G211gat), .Z(new_n920_));
  NAND4_X1  g719(.A1(new_n909_), .A2(new_n528_), .A3(new_n630_), .A4(new_n920_), .ZN(new_n921_));
  AND2_X1   g720(.A1(new_n919_), .A2(new_n921_), .ZN(G1354gat));
  INV_X1    g721(.A(G218gat), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n923_), .B1(new_n910_), .B2(new_n699_), .ZN(new_n924_));
  NAND4_X1  g723(.A1(new_n909_), .A2(G218gat), .A3(new_n528_), .A4(new_n676_), .ZN(new_n925_));
  AND2_X1   g724(.A1(new_n924_), .A2(new_n925_), .ZN(G1355gat));
endmodule


