//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0 0 1 1 0 0 0 0 0 1 0 1 0 1 0 0 1 0 1 1 1 1 1 1 0 0 0 0 0 1 1 1 1 0 1 1 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n744_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n854_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n864_,
    new_n865_, new_n867_, new_n868_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n884_, new_n885_, new_n887_, new_n888_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n913_, new_n914_, new_n915_;
  XOR2_X1   g000(.A(KEYINPUT66), .B(G71gat), .Z(new_n202_));
  INV_X1    g001(.A(G78gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT66), .B(G71gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G78gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G57gat), .B(G64gat), .ZN(new_n207_));
  OAI211_X1 g006(.A(new_n204_), .B(new_n206_), .C1(KEYINPUT11), .C2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT67), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n207_), .A2(KEYINPUT11), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n210_), .A2(new_n211_), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT68), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n210_), .A2(new_n211_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT68), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n216_), .A2(new_n217_), .A3(new_n212_), .ZN(new_n218_));
  AND2_X1   g017(.A1(new_n215_), .A2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(G15gat), .B(G22gat), .ZN(new_n220_));
  INV_X1    g019(.A(G1gat), .ZN(new_n221_));
  INV_X1    g020(.A(G8gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT14), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n220_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G1gat), .B(G8gat), .ZN(new_n225_));
  XOR2_X1   g024(.A(new_n224_), .B(new_n225_), .Z(new_n226_));
  NAND2_X1  g025(.A1(G231gat), .A2(G233gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n226_), .B(new_n227_), .ZN(new_n228_));
  AND2_X1   g027(.A1(new_n219_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT17), .ZN(new_n230_));
  XOR2_X1   g029(.A(G127gat), .B(G155gat), .Z(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(KEYINPUT16), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G183gat), .B(G211gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  NOR3_X1   g033(.A1(new_n229_), .A2(new_n230_), .A3(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n235_), .B1(new_n219_), .B2(new_n228_), .ZN(new_n236_));
  OR3_X1    g035(.A1(new_n213_), .A2(new_n214_), .A3(new_n228_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n228_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n234_), .B(KEYINPUT17), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n237_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n236_), .A2(new_n240_), .ZN(new_n241_));
  AND2_X1   g040(.A1(G155gat), .A2(G162gat), .ZN(new_n242_));
  NOR2_X1   g041(.A1(G155gat), .A2(G162gat), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(KEYINPUT90), .A2(KEYINPUT3), .ZN(new_n245_));
  NOR2_X1   g044(.A1(G141gat), .A2(G148gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(KEYINPUT90), .A2(KEYINPUT3), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n245_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  AND2_X1   g047(.A1(new_n246_), .A2(new_n245_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G141gat), .A2(G148gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT2), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT2), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n253_), .A2(G141gat), .A3(G148gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(KEYINPUT91), .B1(new_n250_), .B2(new_n255_), .ZN(new_n256_));
  OR2_X1    g055(.A1(KEYINPUT90), .A2(KEYINPUT3), .ZN(new_n257_));
  INV_X1    g056(.A(G141gat), .ZN(new_n258_));
  INV_X1    g057(.A(G148gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  AND2_X1   g059(.A1(KEYINPUT90), .A2(KEYINPUT3), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n257_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n246_), .A2(new_n245_), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n262_), .A2(new_n255_), .A3(KEYINPUT91), .A4(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n244_), .B1(new_n256_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT92), .ZN(new_n267_));
  OR2_X1    g066(.A1(new_n246_), .A2(KEYINPUT89), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n246_), .A2(KEYINPUT89), .ZN(new_n269_));
  AOI22_X1  g068(.A1(new_n268_), .A2(new_n269_), .B1(G141gat), .B2(G148gat), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT1), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n242_), .A2(new_n271_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n243_), .A2(KEYINPUT1), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n272_), .B1(new_n273_), .B2(new_n242_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n270_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n266_), .A2(new_n267_), .A3(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n244_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n262_), .A2(new_n255_), .A3(new_n263_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT91), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n277_), .B1(new_n280_), .B2(new_n264_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n275_), .ZN(new_n282_));
  OAI21_X1  g081(.A(KEYINPUT92), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n276_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT29), .ZN(new_n285_));
  AOI21_X1  g084(.A(KEYINPUT93), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT93), .ZN(new_n287_));
  AOI211_X1 g086(.A(new_n287_), .B(KEYINPUT29), .C1(new_n276_), .C2(new_n283_), .ZN(new_n288_));
  OAI21_X1  g087(.A(KEYINPUT28), .B1(new_n286_), .B2(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n267_), .B1(new_n266_), .B2(new_n275_), .ZN(new_n290_));
  NOR3_X1   g089(.A1(new_n281_), .A2(KEYINPUT92), .A3(new_n282_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n285_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(new_n287_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT28), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n284_), .A2(KEYINPUT93), .A3(new_n285_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n293_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  XOR2_X1   g095(.A(G22gat), .B(G50gat), .Z(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  AND3_X1   g097(.A1(new_n289_), .A2(new_n296_), .A3(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n298_), .B1(new_n289_), .B2(new_n296_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G78gat), .B(G106gat), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n276_), .A2(new_n283_), .A3(KEYINPUT29), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G211gat), .B(G218gat), .ZN(new_n304_));
  INV_X1    g103(.A(G197gat), .ZN(new_n305_));
  OAI21_X1  g104(.A(KEYINPUT94), .B1(new_n305_), .B2(G204gat), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n304_), .A2(KEYINPUT21), .A3(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G197gat), .B(G204gat), .ZN(new_n308_));
  OR2_X1    g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n308_), .ZN(new_n310_));
  OR2_X1    g109(.A1(new_n304_), .A2(KEYINPUT21), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n309_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n312_), .B1(G228gat), .B2(G233gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n303_), .A2(KEYINPUT95), .A3(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n285_), .B1(new_n266_), .B2(new_n275_), .ZN(new_n315_));
  OAI211_X1 g114(.A(G228gat), .B(G233gat), .C1(new_n315_), .C2(new_n312_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(KEYINPUT95), .B1(new_n303_), .B2(new_n313_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n302_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(KEYINPUT96), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT97), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n303_), .A2(new_n313_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT95), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n302_), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n325_), .A2(new_n314_), .A3(new_n316_), .A4(new_n326_), .ZN(new_n327_));
  AND3_X1   g126(.A1(new_n319_), .A2(new_n322_), .A3(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n322_), .B1(new_n319_), .B2(new_n327_), .ZN(new_n329_));
  OAI22_X1  g128(.A1(new_n301_), .A2(new_n321_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n289_), .A2(new_n296_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(new_n297_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n289_), .A2(new_n296_), .A3(new_n298_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n319_), .A2(new_n327_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(KEYINPUT97), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n319_), .A2(new_n322_), .A3(new_n327_), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n334_), .A2(new_n336_), .A3(new_n320_), .A4(new_n337_), .ZN(new_n338_));
  AND2_X1   g137(.A1(new_n330_), .A2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G127gat), .B(G134gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G113gat), .B(G120gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  OR2_X1    g141(.A1(new_n340_), .A2(new_n341_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT87), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n342_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n345_), .B1(new_n344_), .B2(new_n343_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n276_), .A2(new_n283_), .A3(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n343_), .A2(new_n342_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n266_), .A2(new_n275_), .A3(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G225gat), .A2(G233gat), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n347_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G1gat), .B(G29gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT0), .ZN(new_n353_));
  INV_X1    g152(.A(G57gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(G85gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  AND3_X1   g157(.A1(new_n347_), .A2(KEYINPUT4), .A3(new_n349_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n350_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n360_), .B1(new_n347_), .B2(KEYINPUT4), .ZN(new_n361_));
  OAI211_X1 g160(.A(new_n351_), .B(new_n358_), .C1(new_n359_), .C2(new_n361_), .ZN(new_n362_));
  OR2_X1    g161(.A1(KEYINPUT101), .A2(KEYINPUT33), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT98), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT20), .ZN(new_n366_));
  INV_X1    g165(.A(G190gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT81), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT81), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(G190gat), .ZN(new_n370_));
  AND3_X1   g169(.A1(new_n368_), .A2(new_n370_), .A3(KEYINPUT26), .ZN(new_n371_));
  INV_X1    g170(.A(G183gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(KEYINPUT25), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT25), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(G183gat), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n373_), .B(new_n375_), .C1(KEYINPUT26), .C2(new_n367_), .ZN(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT82), .B1(new_n371_), .B2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G169gat), .A2(G176gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(KEYINPUT24), .ZN(new_n379_));
  NOR2_X1   g178(.A1(G169gat), .A2(G176gat), .ZN(new_n380_));
  MUX2_X1   g179(.A(new_n379_), .B(KEYINPUT24), .S(new_n380_), .Z(new_n381_));
  NAND2_X1  g180(.A1(G183gat), .A2(G190gat), .ZN(new_n382_));
  AOI21_X1  g181(.A(KEYINPUT83), .B1(new_n382_), .B2(KEYINPUT23), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT23), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n385_), .A2(G183gat), .A3(G190gat), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n382_), .A2(KEYINPUT83), .A3(KEYINPUT23), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n384_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n368_), .A2(new_n370_), .A3(KEYINPUT26), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT82), .ZN(new_n390_));
  OR2_X1    g189(.A1(new_n367_), .A2(KEYINPUT26), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT25), .B(G183gat), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n389_), .A2(new_n390_), .A3(new_n391_), .A4(new_n392_), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n377_), .A2(new_n381_), .A3(new_n388_), .A4(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n368_), .A2(new_n370_), .A3(new_n372_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n382_), .A2(KEYINPUT23), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(new_n386_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n395_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(G169gat), .ZN(new_n399_));
  OR3_X1    g198(.A1(new_n399_), .A2(KEYINPUT84), .A3(KEYINPUT22), .ZN(new_n400_));
  INV_X1    g199(.A(G176gat), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT22), .B1(new_n399_), .B2(KEYINPUT84), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n400_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n398_), .A2(new_n403_), .A3(new_n378_), .ZN(new_n404_));
  AND3_X1   g203(.A1(new_n394_), .A2(KEYINPUT85), .A3(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(KEYINPUT85), .B1(new_n394_), .B2(new_n404_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n312_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n392_), .ZN(new_n408_));
  XOR2_X1   g207(.A(KEYINPUT26), .B(G190gat), .Z(new_n409_));
  OAI211_X1 g208(.A(new_n381_), .B(new_n397_), .C1(new_n408_), .C2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n387_), .A2(new_n386_), .ZN(new_n411_));
  OAI22_X1  g210(.A1(new_n411_), .A2(new_n383_), .B1(G183gat), .B2(G190gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT22), .B(G169gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(new_n401_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n412_), .A2(new_n378_), .A3(new_n414_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n410_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n312_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n366_), .B1(new_n407_), .B2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G226gat), .A2(G233gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(KEYINPUT19), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n365_), .B1(new_n419_), .B2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n394_), .A2(new_n404_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT85), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n394_), .A2(KEYINPUT85), .A3(new_n404_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n417_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n418_), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT20), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n430_), .A2(KEYINPUT98), .A3(new_n421_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n417_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n421_), .B1(new_n416_), .B2(new_n312_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n432_), .A2(KEYINPUT20), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT99), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n432_), .A2(KEYINPUT99), .A3(KEYINPUT20), .A4(new_n433_), .ZN(new_n437_));
  AOI22_X1  g236(.A1(new_n423_), .A2(new_n431_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G8gat), .B(G36gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(KEYINPUT18), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT100), .ZN(new_n441_));
  XOR2_X1   g240(.A(G64gat), .B(G92gat), .Z(new_n442_));
  XNOR2_X1  g241(.A(new_n441_), .B(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n438_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n436_), .A2(new_n437_), .ZN(new_n445_));
  NOR3_X1   g244(.A1(new_n419_), .A2(new_n365_), .A3(new_n422_), .ZN(new_n446_));
  AOI21_X1  g245(.A(KEYINPUT98), .B1(new_n430_), .B2(new_n421_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n445_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n443_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n347_), .A2(new_n349_), .ZN(new_n451_));
  OR2_X1    g250(.A1(new_n451_), .A2(KEYINPUT102), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(KEYINPUT102), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n350_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  OR2_X1    g253(.A1(new_n347_), .A2(KEYINPUT4), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n347_), .A2(KEYINPUT4), .A3(new_n349_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n360_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n357_), .B1(new_n454_), .B2(new_n457_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n364_), .A2(new_n444_), .A3(new_n450_), .A4(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n351_), .B1(new_n359_), .B2(new_n361_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(new_n357_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(new_n362_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n443_), .A2(KEYINPUT32), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n445_), .B(new_n463_), .C1(new_n446_), .C2(new_n447_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n463_), .ZN(new_n465_));
  AND3_X1   g264(.A1(new_n410_), .A2(new_n415_), .A3(KEYINPUT103), .ZN(new_n466_));
  AOI21_X1  g265(.A(KEYINPUT103), .B1(new_n410_), .B2(new_n415_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n312_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n432_), .A2(new_n468_), .A3(KEYINPUT20), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n469_), .A2(KEYINPUT104), .A3(new_n421_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n419_), .A2(new_n422_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(KEYINPUT104), .B1(new_n469_), .B2(new_n421_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n465_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n462_), .A2(new_n464_), .A3(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT105), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n462_), .A2(new_n464_), .A3(new_n474_), .A4(KEYINPUT105), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n459_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n462_), .B1(new_n330_), .B2(new_n338_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n450_), .A2(new_n444_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT27), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n449_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n482_), .B1(new_n438_), .B2(new_n443_), .ZN(new_n484_));
  AOI22_X1  g283(.A1(new_n481_), .A2(new_n482_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  AOI22_X1  g284(.A1(new_n339_), .A2(new_n479_), .B1(new_n480_), .B2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n426_), .A2(new_n427_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(KEYINPUT30), .ZN(new_n488_));
  XOR2_X1   g287(.A(G71gat), .B(G99gat), .Z(new_n489_));
  NAND2_X1  g288(.A1(G227gat), .A2(G233gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G15gat), .B(G43gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT86), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n491_), .B(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n488_), .B(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT88), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n346_), .B(KEYINPUT31), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  OAI21_X1  g298(.A(KEYINPUT106), .B1(new_n486_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n339_), .A2(new_n479_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n330_), .A2(new_n338_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n462_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n502_), .A2(new_n485_), .A3(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n501_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT106), .ZN(new_n506_));
  INV_X1    g305(.A(new_n499_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n505_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n485_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n509_), .A2(new_n502_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n507_), .A2(new_n462_), .ZN(new_n511_));
  AOI22_X1  g310(.A1(new_n500_), .A2(new_n508_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G232gat), .A2(G233gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT34), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT35), .ZN(new_n515_));
  XOR2_X1   g314(.A(new_n515_), .B(KEYINPUT71), .Z(new_n516_));
  NOR2_X1   g315(.A1(new_n514_), .A2(KEYINPUT35), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT72), .ZN(new_n518_));
  NOR2_X1   g317(.A1(G99gat), .A2(G106gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT7), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G99gat), .A2(G106gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT6), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  XOR2_X1   g322(.A(G85gat), .B(G92gat), .Z(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT8), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n523_), .A2(KEYINPUT8), .A3(new_n524_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(KEYINPUT10), .B(G99gat), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT64), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(G106gat), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT9), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(KEYINPUT65), .ZN(new_n535_));
  OR2_X1    g334(.A1(new_n534_), .A2(KEYINPUT65), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n524_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G85gat), .A2(G92gat), .ZN(new_n538_));
  OAI211_X1 g337(.A(new_n537_), .B(new_n522_), .C1(new_n538_), .C2(new_n535_), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n527_), .B(new_n528_), .C1(new_n533_), .C2(new_n539_), .ZN(new_n540_));
  XOR2_X1   g339(.A(G29gat), .B(G36gat), .Z(new_n541_));
  XNOR2_X1  g340(.A(G43gat), .B(G50gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n518_), .B1(new_n540_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT15), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n543_), .B(new_n545_), .ZN(new_n546_));
  AOI211_X1 g345(.A(new_n516_), .B(new_n544_), .C1(new_n546_), .C2(new_n540_), .ZN(new_n547_));
  AND2_X1   g346(.A1(new_n544_), .A2(KEYINPUT73), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n540_), .A2(new_n546_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n549_), .B1(new_n544_), .B2(KEYINPUT73), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n516_), .B1(new_n548_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT74), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n551_), .A2(new_n552_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n547_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G190gat), .B(G218gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT75), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G134gat), .B(G162gat), .ZN(new_n558_));
  XOR2_X1   g357(.A(new_n557_), .B(new_n558_), .Z(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n560_), .A2(KEYINPUT36), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n555_), .A2(new_n561_), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n559_), .B(KEYINPUT36), .Z(new_n563_));
  OAI21_X1  g362(.A(new_n562_), .B1(new_n563_), .B2(new_n555_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT108), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(KEYINPUT109), .B1(new_n512_), .B2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n510_), .A2(new_n511_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n506_), .B1(new_n505_), .B2(new_n507_), .ZN(new_n570_));
  AOI211_X1 g369(.A(KEYINPUT106), .B(new_n499_), .C1(new_n501_), .C2(new_n504_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n569_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT109), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n572_), .A2(new_n573_), .A3(new_n566_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n241_), .B1(new_n568_), .B2(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n216_), .A2(new_n540_), .A3(new_n212_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n540_), .B1(new_n216_), .B2(new_n212_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT12), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n576_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G230gat), .A2(G233gat), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n540_), .A2(KEYINPUT12), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n215_), .A2(new_n218_), .A3(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n579_), .A2(new_n580_), .A3(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n576_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n584_), .A2(new_n577_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n583_), .B1(new_n580_), .B2(new_n585_), .ZN(new_n586_));
  XOR2_X1   g385(.A(G120gat), .B(G148gat), .Z(new_n587_));
  XNOR2_X1  g386(.A(G176gat), .B(G204gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(KEYINPUT69), .B(KEYINPUT5), .Z(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT70), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n589_), .B(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n586_), .A2(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n586_), .A2(new_n593_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  OR2_X1    g395(.A1(new_n596_), .A2(KEYINPUT13), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(KEYINPUT13), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n543_), .B(KEYINPUT78), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(new_n226_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n226_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n546_), .A2(new_n602_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n601_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(G229gat), .A2(G233gat), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n600_), .B(new_n602_), .ZN(new_n607_));
  OAI22_X1  g406(.A1(new_n606_), .A2(KEYINPUT79), .B1(new_n605_), .B2(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n608_), .B1(KEYINPUT79), .B2(new_n606_), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n609_), .A2(KEYINPUT80), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G113gat), .B(G141gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G169gat), .B(G197gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n610_), .B(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n599_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n575_), .A2(new_n617_), .ZN(new_n618_));
  OAI21_X1  g417(.A(G1gat), .B1(new_n618_), .B2(new_n503_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n617_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n512_), .A2(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n563_), .B(KEYINPUT76), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n555_), .A2(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n623_), .B1(new_n561_), .B2(new_n555_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT37), .ZN(new_n625_));
  XOR2_X1   g424(.A(KEYINPUT77), .B(KEYINPUT37), .Z(new_n626_));
  OAI22_X1  g425(.A1(new_n624_), .A2(new_n625_), .B1(new_n564_), .B2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n628_), .A2(new_n241_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n621_), .A2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n630_), .A2(new_n221_), .A3(new_n462_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT107), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n632_), .A2(KEYINPUT38), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n632_), .A2(KEYINPUT38), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n619_), .B1(new_n633_), .B2(new_n634_), .ZN(G1324gat));
  NAND3_X1  g434(.A1(new_n630_), .A2(new_n222_), .A3(new_n509_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n575_), .A2(new_n617_), .A3(new_n509_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT39), .ZN(new_n638_));
  AND3_X1   g437(.A1(new_n637_), .A2(new_n638_), .A3(G8gat), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n638_), .B1(new_n637_), .B2(G8gat), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n636_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT40), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  OAI211_X1 g442(.A(KEYINPUT40), .B(new_n636_), .C1(new_n639_), .C2(new_n640_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(G1325gat));
  OAI21_X1  g444(.A(G15gat), .B1(new_n618_), .B2(new_n507_), .ZN(new_n646_));
  XOR2_X1   g445(.A(KEYINPUT110), .B(KEYINPUT41), .Z(new_n647_));
  OR2_X1    g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n647_), .ZN(new_n649_));
  INV_X1    g448(.A(G15gat), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n630_), .A2(new_n650_), .A3(new_n499_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n648_), .A2(new_n649_), .A3(new_n651_), .ZN(G1326gat));
  INV_X1    g451(.A(G22gat), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n630_), .A2(new_n653_), .A3(new_n502_), .ZN(new_n654_));
  OAI21_X1  g453(.A(G22gat), .B1(new_n618_), .B2(new_n339_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n655_), .A2(KEYINPUT42), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n655_), .A2(KEYINPUT42), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n654_), .B1(new_n656_), .B2(new_n657_), .ZN(G1327gat));
  INV_X1    g457(.A(new_n241_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n659_), .A2(new_n564_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n621_), .A2(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(G29gat), .B1(new_n661_), .B2(new_n462_), .ZN(new_n662_));
  OAI21_X1  g461(.A(KEYINPUT43), .B1(new_n512_), .B2(new_n627_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT43), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n572_), .A2(new_n664_), .A3(new_n628_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n663_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT111), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT44), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n620_), .A2(new_n659_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n666_), .A2(new_n669_), .A3(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n669_), .B1(new_n666_), .B2(new_n670_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n462_), .A2(G29gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n662_), .B1(new_n674_), .B2(new_n675_), .ZN(G1328gat));
  INV_X1    g475(.A(KEYINPUT45), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n485_), .A2(G36gat), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n621_), .A2(new_n677_), .A3(new_n660_), .A4(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT112), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n621_), .A2(new_n660_), .A3(new_n678_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n681_), .B1(KEYINPUT45), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n673_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n684_), .A2(new_n509_), .A3(new_n671_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n680_), .A2(G36gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n683_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT46), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  AOI211_X1 g488(.A(KEYINPUT46), .B(new_n683_), .C1(new_n685_), .C2(new_n686_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n689_), .A2(new_n690_), .ZN(G1329gat));
  INV_X1    g490(.A(G43gat), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n661_), .A2(new_n692_), .A3(new_n499_), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n672_), .A2(new_n673_), .A3(new_n507_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n693_), .B1(new_n694_), .B2(new_n692_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT47), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  OAI211_X1 g496(.A(KEYINPUT47), .B(new_n693_), .C1(new_n694_), .C2(new_n692_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(G1330gat));
  AOI21_X1  g498(.A(G50gat), .B1(new_n661_), .B2(new_n502_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n502_), .A2(G50gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n700_), .B1(new_n674_), .B2(new_n701_), .ZN(G1331gat));
  INV_X1    g501(.A(new_n599_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n703_), .A2(new_n615_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n572_), .A2(new_n704_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n705_), .A2(new_n629_), .ZN(new_n706_));
  AOI21_X1  g505(.A(G57gat), .B1(new_n706_), .B2(new_n462_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n575_), .A2(new_n704_), .ZN(new_n708_));
  NOR3_X1   g507(.A1(new_n708_), .A2(new_n354_), .A3(new_n503_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT113), .ZN(new_n710_));
  OR2_X1    g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n709_), .A2(new_n710_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n707_), .B1(new_n711_), .B2(new_n712_), .ZN(G1332gat));
  INV_X1    g512(.A(G64gat), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n706_), .A2(new_n714_), .A3(new_n509_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT48), .ZN(new_n716_));
  INV_X1    g515(.A(new_n708_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(new_n509_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n716_), .B1(new_n718_), .B2(G64gat), .ZN(new_n719_));
  AOI211_X1 g518(.A(KEYINPUT48), .B(new_n714_), .C1(new_n717_), .C2(new_n509_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n715_), .B1(new_n719_), .B2(new_n720_), .ZN(G1333gat));
  INV_X1    g520(.A(G71gat), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n706_), .A2(new_n722_), .A3(new_n499_), .ZN(new_n723_));
  OAI21_X1  g522(.A(G71gat), .B1(new_n708_), .B2(new_n507_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n724_), .A2(KEYINPUT49), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n724_), .A2(KEYINPUT49), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n723_), .B1(new_n725_), .B2(new_n726_), .ZN(G1334gat));
  NAND3_X1  g526(.A1(new_n706_), .A2(new_n203_), .A3(new_n502_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n575_), .A2(new_n502_), .A3(new_n704_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT50), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n729_), .A2(new_n730_), .A3(G78gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n729_), .B2(G78gat), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n728_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(KEYINPUT114), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT114), .ZN(new_n735_));
  OAI211_X1 g534(.A(new_n735_), .B(new_n728_), .C1(new_n731_), .C2(new_n732_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(G1335gat));
  NOR3_X1   g536(.A1(new_n703_), .A2(new_n615_), .A3(new_n659_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n666_), .A2(new_n738_), .ZN(new_n739_));
  OAI21_X1  g538(.A(G85gat), .B1(new_n739_), .B2(new_n503_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n705_), .A2(new_n660_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n741_), .A2(new_n356_), .A3(new_n462_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(G1336gat));
  OAI21_X1  g542(.A(G92gat), .B1(new_n739_), .B2(new_n485_), .ZN(new_n744_));
  INV_X1    g543(.A(G92gat), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n741_), .A2(new_n745_), .A3(new_n509_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(new_n746_), .ZN(G1337gat));
  NOR2_X1   g546(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n748_));
  OAI21_X1  g547(.A(G99gat), .B1(new_n739_), .B2(new_n507_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n741_), .A2(new_n531_), .A3(new_n499_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n748_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n752_));
  XOR2_X1   g551(.A(new_n751_), .B(new_n752_), .Z(G1338gat));
  NOR3_X1   g552(.A1(new_n512_), .A2(KEYINPUT43), .A3(new_n627_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n664_), .B1(new_n572_), .B2(new_n628_), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n502_), .B(new_n738_), .C1(new_n754_), .C2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT52), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n756_), .A2(new_n757_), .A3(G106gat), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT116), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n756_), .A2(KEYINPUT116), .A3(new_n757_), .A4(G106gat), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n756_), .A2(G106gat), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(KEYINPUT52), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n760_), .A2(new_n761_), .A3(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n741_), .A2(new_n532_), .A3(new_n502_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT53), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT53), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n764_), .A2(new_n768_), .A3(new_n765_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(G1339gat));
  NOR2_X1   g569(.A1(new_n599_), .A2(new_n615_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n629_), .A2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT54), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n629_), .A2(KEYINPUT54), .A3(new_n771_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT121), .ZN(new_n777_));
  INV_X1    g576(.A(new_n595_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n605_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n607_), .A2(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(KEYINPUT119), .B1(new_n780_), .B2(new_n614_), .ZN(new_n781_));
  NOR3_X1   g580(.A1(new_n780_), .A2(KEYINPUT119), .A3(new_n614_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n782_), .B1(new_n779_), .B2(new_n604_), .ZN(new_n783_));
  AOI22_X1  g582(.A1(new_n781_), .A2(new_n783_), .B1(new_n609_), .B2(new_n614_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n579_), .A2(KEYINPUT55), .A3(new_n582_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n580_), .A2(KEYINPUT117), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n583_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n786_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n579_), .A2(new_n582_), .A3(KEYINPUT55), .A4(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n787_), .A2(new_n789_), .A3(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT118), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT118), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n787_), .A2(new_n789_), .A3(new_n794_), .A4(new_n791_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n793_), .A2(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(KEYINPUT56), .B1(new_n796_), .B2(new_n593_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT56), .ZN(new_n798_));
  AOI211_X1 g597(.A(new_n798_), .B(new_n592_), .C1(new_n793_), .C2(new_n795_), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n778_), .B(new_n784_), .C1(new_n797_), .C2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT58), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n777_), .B1(new_n802_), .B2(new_n627_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n800_), .A2(new_n801_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n627_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n804_), .B1(new_n805_), .B2(KEYINPUT121), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n803_), .A2(new_n806_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n615_), .B(new_n778_), .C1(new_n797_), .C2(new_n799_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n784_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n809_));
  XOR2_X1   g608(.A(new_n809_), .B(KEYINPUT120), .Z(new_n810_));
  NAND2_X1  g609(.A1(new_n808_), .A2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT57), .B1(new_n811_), .B2(new_n564_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT57), .ZN(new_n813_));
  INV_X1    g612(.A(new_n564_), .ZN(new_n814_));
  AOI211_X1 g613(.A(new_n813_), .B(new_n814_), .C1(new_n808_), .C2(new_n810_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n812_), .A2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n807_), .A2(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n776_), .B1(new_n817_), .B2(new_n241_), .ZN(new_n818_));
  NOR4_X1   g617(.A1(new_n509_), .A2(new_n507_), .A3(new_n503_), .A4(new_n502_), .ZN(new_n819_));
  XOR2_X1   g618(.A(new_n819_), .B(KEYINPUT122), .Z(new_n820_));
  NOR2_X1   g619(.A1(new_n818_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(G113gat), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n821_), .A2(new_n822_), .A3(new_n615_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n805_), .A2(KEYINPUT121), .ZN(new_n824_));
  AOI211_X1 g623(.A(new_n777_), .B(new_n627_), .C1(new_n800_), .C2(new_n801_), .ZN(new_n825_));
  NOR3_X1   g624(.A1(new_n824_), .A2(new_n825_), .A3(new_n804_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n814_), .B1(new_n808_), .B2(new_n810_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(KEYINPUT57), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n241_), .B1(new_n826_), .B2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n776_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n820_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n831_), .A2(KEYINPUT59), .A3(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT59), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n834_), .B1(new_n818_), .B2(new_n820_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n616_), .B1(new_n833_), .B2(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n823_), .B1(new_n836_), .B2(new_n822_), .ZN(G1340gat));
  INV_X1    g636(.A(KEYINPUT60), .ZN(new_n838_));
  XNOR2_X1  g637(.A(KEYINPUT123), .B(G120gat), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n599_), .A2(new_n838_), .A3(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n821_), .A2(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n703_), .B1(new_n833_), .B2(new_n835_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(new_n839_), .ZN(G1341gat));
  NAND2_X1  g643(.A1(new_n659_), .A2(G127gat), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n845_), .B1(new_n833_), .B2(new_n835_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n659_), .B1(new_n807_), .B2(new_n816_), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n659_), .B(new_n832_), .C1(new_n847_), .C2(new_n776_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT124), .ZN(new_n849_));
  INV_X1    g648(.A(G127gat), .ZN(new_n850_));
  AND3_X1   g649(.A1(new_n848_), .A2(new_n849_), .A3(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n849_), .B1(new_n848_), .B2(new_n850_), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n846_), .A2(new_n851_), .A3(new_n852_), .ZN(G1342gat));
  INV_X1    g652(.A(G134gat), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n821_), .A2(new_n854_), .A3(new_n567_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n627_), .B1(new_n833_), .B2(new_n835_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n855_), .B1(new_n856_), .B2(new_n854_), .ZN(G1343gat));
  NOR4_X1   g656(.A1(new_n509_), .A2(new_n339_), .A3(new_n503_), .A4(new_n499_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n831_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n860_), .A2(new_n258_), .A3(new_n615_), .ZN(new_n861_));
  OAI21_X1  g660(.A(G141gat), .B1(new_n859_), .B2(new_n616_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(G1344gat));
  NAND3_X1  g662(.A1(new_n860_), .A2(new_n259_), .A3(new_n599_), .ZN(new_n864_));
  OAI21_X1  g663(.A(G148gat), .B1(new_n859_), .B2(new_n703_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(G1345gat));
  NAND3_X1  g665(.A1(new_n831_), .A2(new_n659_), .A3(new_n858_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(KEYINPUT61), .B(G155gat), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n867_), .B(new_n868_), .ZN(G1346gat));
  OR3_X1    g668(.A1(new_n859_), .A2(G162gat), .A3(new_n566_), .ZN(new_n870_));
  OAI21_X1  g669(.A(G162gat), .B1(new_n859_), .B2(new_n627_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(G1347gat));
  NOR4_X1   g671(.A1(new_n507_), .A2(new_n502_), .A3(new_n485_), .A4(new_n462_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n831_), .A2(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(G169gat), .B1(new_n874_), .B2(new_n616_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT62), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  OAI211_X1 g676(.A(KEYINPUT62), .B(G169gat), .C1(new_n874_), .C2(new_n616_), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n831_), .A2(new_n873_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n879_), .A2(new_n615_), .A3(new_n413_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n877_), .A2(new_n878_), .A3(new_n880_), .ZN(G1348gat));
  NAND3_X1  g680(.A1(new_n831_), .A2(new_n599_), .A3(new_n873_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g682(.A1(new_n879_), .A2(new_n659_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(G183gat), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n885_), .B1(new_n408_), .B2(new_n884_), .ZN(G1350gat));
  OAI21_X1  g685(.A(G190gat), .B1(new_n874_), .B2(new_n627_), .ZN(new_n887_));
  OR2_X1    g686(.A1(new_n566_), .A2(new_n409_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n874_), .B2(new_n888_), .ZN(G1351gat));
  INV_X1    g688(.A(KEYINPUT125), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n509_), .A2(new_n507_), .A3(new_n480_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n818_), .B2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n891_), .ZN(new_n893_));
  OAI211_X1 g692(.A(KEYINPUT125), .B(new_n893_), .C1(new_n847_), .C2(new_n776_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n894_), .ZN(new_n895_));
  AOI21_X1  g694(.A(G197gat), .B1(new_n895_), .B2(new_n615_), .ZN(new_n896_));
  AOI211_X1 g695(.A(new_n305_), .B(new_n616_), .C1(new_n892_), .C2(new_n894_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n896_), .A2(new_n897_), .ZN(G1352gat));
  AOI21_X1  g697(.A(KEYINPUT125), .B1(new_n831_), .B2(new_n893_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n894_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n599_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n901_));
  XOR2_X1   g700(.A(KEYINPUT126), .B(G204gat), .Z(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n902_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n895_), .A2(new_n599_), .A3(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n903_), .A2(new_n905_), .ZN(G1353gat));
  AOI21_X1  g705(.A(new_n241_), .B1(new_n892_), .B2(new_n894_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(KEYINPUT63), .B(G211gat), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n909_), .B1(new_n907_), .B2(new_n910_), .ZN(G1354gat));
  NAND2_X1  g710(.A1(new_n895_), .A2(new_n567_), .ZN(new_n912_));
  INV_X1    g711(.A(G218gat), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n628_), .A2(G218gat), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(KEYINPUT127), .ZN(new_n915_));
  AOI22_X1  g714(.A1(new_n912_), .A2(new_n913_), .B1(new_n895_), .B2(new_n915_), .ZN(G1355gat));
endmodule


