//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 0 1 0 0 0 1 0 0 1 1 0 0 0 1 1 1 0 1 1 0 1 1 1 1 1 1 1 1 0 0 0 1 1 1 0 1 1 0 1 1 1 0 1 1 1 1 0 1 1 0 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n575_,
    new_n576_, new_n577_, new_n578_, new_n579_, new_n581_, new_n582_,
    new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n629_, new_n630_, new_n631_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n655_, new_n656_,
    new_n657_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n667_, new_n668_, new_n669_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n782_, new_n783_, new_n784_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n792_,
    new_n793_, new_n795_, new_n796_, new_n798_, new_n799_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n811_, new_n812_, new_n813_, new_n815_,
    new_n816_, new_n818_, new_n819_, new_n821_, new_n822_, new_n823_,
    new_n825_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n833_, new_n834_, new_n835_;
  XNOR2_X1  g000(.A(KEYINPUT22), .B(G169gat), .ZN(new_n202_));
  INV_X1    g001(.A(G176gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT83), .ZN(new_n206_));
  AND2_X1   g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT84), .B(KEYINPUT23), .ZN(new_n208_));
  INV_X1    g007(.A(G183gat), .ZN(new_n209_));
  INV_X1    g008(.A(G190gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n208_), .A2(new_n211_), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n212_), .B1(KEYINPUT23), .B2(new_n211_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n207_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT85), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n208_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT23), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n211_), .A2(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n216_), .B1(new_n217_), .B2(new_n219_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n220_), .B1(new_n216_), .B2(new_n219_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n222_), .B(KEYINPUT82), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(KEYINPUT24), .A3(new_n206_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT26), .B(G190gat), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT25), .B1(new_n209_), .B2(KEYINPUT81), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n209_), .A2(KEYINPUT25), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n225_), .B(new_n226_), .C1(new_n227_), .C2(KEYINPUT81), .ZN(new_n228_));
  OAI211_X1 g027(.A(new_n224_), .B(new_n228_), .C1(KEYINPUT24), .C2(new_n223_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n215_), .B1(new_n221_), .B2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G71gat), .B(G99gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(G43gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n230_), .B(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G127gat), .B(G134gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G113gat), .B(G120gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n233_), .B(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G227gat), .A2(G233gat), .ZN(new_n238_));
  XOR2_X1   g037(.A(new_n238_), .B(G15gat), .Z(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT30), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(KEYINPUT31), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n237_), .B(new_n241_), .ZN(new_n242_));
  XOR2_X1   g041(.A(G155gat), .B(G162gat), .Z(new_n243_));
  OR2_X1    g042(.A1(G141gat), .A2(G148gat), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT2), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G141gat), .A2(G148gat), .ZN(new_n246_));
  AOI22_X1  g045(.A1(new_n244_), .A2(KEYINPUT3), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n247_), .B1(KEYINPUT3), .B2(new_n244_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT86), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n243_), .B1(new_n248_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT1), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n243_), .A2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n253_), .A2(new_n254_), .A3(new_n244_), .A4(new_n246_), .ZN(new_n255_));
  AND2_X1   g054(.A1(new_n251_), .A2(new_n255_), .ZN(new_n256_));
  OR2_X1    g055(.A1(new_n256_), .A2(new_n236_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n236_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G225gat), .A2(G233gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n257_), .A2(KEYINPUT4), .A3(new_n258_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT95), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT95), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n257_), .A2(new_n264_), .A3(KEYINPUT4), .A4(new_n258_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n257_), .ZN(new_n266_));
  XOR2_X1   g065(.A(KEYINPUT96), .B(KEYINPUT4), .Z(new_n267_));
  AOI22_X1  g066(.A1(new_n263_), .A2(new_n265_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n261_), .B1(new_n268_), .B2(new_n260_), .ZN(new_n269_));
  XOR2_X1   g068(.A(G1gat), .B(G29gat), .Z(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT97), .B(G85gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT0), .B(G57gat), .ZN(new_n273_));
  XOR2_X1   g072(.A(new_n272_), .B(new_n273_), .Z(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n269_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT33), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n269_), .A2(KEYINPUT33), .A3(new_n275_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n268_), .A2(new_n260_), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n280_), .B(new_n274_), .C1(new_n260_), .C2(new_n259_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n278_), .A2(new_n279_), .A3(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n207_), .B(KEYINPUT91), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n283_), .B1(new_n221_), .B2(new_n214_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n223_), .A2(KEYINPUT24), .A3(new_n205_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT25), .B(G183gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n225_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  OR2_X1    g087(.A1(new_n288_), .A2(KEYINPUT90), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(KEYINPUT90), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT24), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n213_), .B1(new_n291_), .B2(new_n222_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n289_), .A2(new_n290_), .A3(new_n292_), .ZN(new_n293_));
  XOR2_X1   g092(.A(G197gat), .B(G204gat), .Z(new_n294_));
  OR2_X1    g093(.A1(new_n294_), .A2(KEYINPUT21), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(KEYINPUT21), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G211gat), .B(G218gat), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n295_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  OR2_X1    g097(.A1(new_n296_), .A2(new_n297_), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n284_), .A2(new_n293_), .A3(new_n298_), .A4(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G226gat), .A2(G233gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT19), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT20), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n298_), .A2(new_n299_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n304_), .B1(new_n230_), .B2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n300_), .A2(new_n303_), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT92), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  AOI22_X1  g108(.A1(new_n284_), .A2(new_n293_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n310_));
  OAI21_X1  g109(.A(KEYINPUT20), .B1(new_n230_), .B2(new_n305_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n302_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n300_), .A2(KEYINPUT92), .A3(new_n303_), .A4(new_n306_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n309_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  XOR2_X1   g113(.A(G8gat), .B(G36gat), .Z(new_n315_));
  XNOR2_X1  g114(.A(G64gat), .B(G92gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n314_), .A2(new_n320_), .ZN(new_n321_));
  NAND4_X1  g120(.A1(new_n309_), .A2(new_n319_), .A3(new_n312_), .A4(new_n313_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n321_), .A2(KEYINPUT94), .A3(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT94), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n314_), .A2(new_n324_), .A3(new_n320_), .ZN(new_n325_));
  AND2_X1   g124(.A1(new_n323_), .A2(new_n325_), .ZN(new_n326_));
  OAI211_X1 g125(.A(new_n274_), .B(new_n261_), .C1(new_n268_), .C2(new_n260_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n276_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n319_), .A2(KEYINPUT32), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NOR3_X1   g130(.A1(new_n310_), .A2(new_n302_), .A3(new_n311_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n303_), .B1(new_n300_), .B2(new_n306_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n331_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n334_), .B1(new_n314_), .B2(new_n331_), .ZN(new_n335_));
  OAI22_X1  g134(.A1(new_n282_), .A2(new_n326_), .B1(new_n329_), .B2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT29), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n305_), .B1(new_n256_), .B2(new_n337_), .ZN(new_n338_));
  AND3_X1   g137(.A1(KEYINPUT88), .A2(G228gat), .A3(G233gat), .ZN(new_n339_));
  AOI21_X1  g138(.A(KEYINPUT88), .B1(G228gat), .B2(G233gat), .ZN(new_n340_));
  OR2_X1    g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n338_), .A2(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n338_), .A2(new_n339_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G78gat), .B(G106gat), .ZN(new_n344_));
  OR3_X1    g143(.A1(new_n342_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT89), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n256_), .A2(new_n337_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G22gat), .B(G50gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n347_), .B(new_n350_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n344_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n352_));
  AOI22_X1  g151(.A1(new_n346_), .A2(new_n351_), .B1(new_n352_), .B2(new_n345_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT89), .ZN(new_n354_));
  AND4_X1   g153(.A1(new_n354_), .A2(new_n345_), .A3(new_n352_), .A4(new_n351_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n353_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT27), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n323_), .A2(new_n357_), .A3(new_n325_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n356_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n320_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n322_), .A2(KEYINPUT27), .A3(new_n360_), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n358_), .A2(new_n359_), .A3(new_n329_), .A4(new_n361_), .ZN(new_n362_));
  AOI22_X1  g161(.A1(new_n336_), .A2(new_n356_), .B1(new_n362_), .B2(KEYINPUT98), .ZN(new_n363_));
  OR2_X1    g162(.A1(new_n362_), .A2(KEYINPUT98), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n242_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n358_), .A2(new_n361_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n366_), .A2(new_n359_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n242_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n368_), .A2(new_n328_), .ZN(new_n369_));
  AND2_X1   g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n365_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT65), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT6), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT64), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT64), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT6), .ZN(new_n376_));
  AND2_X1   g175(.A1(G99gat), .A2(G106gat), .ZN(new_n377_));
  AND3_X1   g176(.A1(new_n374_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n377_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n372_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G99gat), .A2(G106gat), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n375_), .A2(KEYINPUT6), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n373_), .A2(KEYINPUT64), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n381_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n374_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n384_), .A2(KEYINPUT65), .A3(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NOR3_X1   g187(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n380_), .A2(new_n386_), .A3(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G85gat), .B(G92gat), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n392_), .A2(KEYINPUT8), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n391_), .A2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n390_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n392_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT8), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n394_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT9), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n400_), .A2(G85gat), .A3(G92gat), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n401_), .B1(new_n392_), .B2(new_n400_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(KEYINPUT10), .B(G99gat), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n403_), .A2(G106gat), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n405_), .A2(new_n386_), .A3(new_n380_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n399_), .A2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G29gat), .B(G36gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G43gat), .B(G50gat), .ZN(new_n409_));
  XOR2_X1   g208(.A(new_n408_), .B(new_n409_), .Z(new_n410_));
  XOR2_X1   g209(.A(new_n410_), .B(KEYINPUT15), .Z(new_n411_));
  NAND2_X1  g210(.A1(new_n407_), .A2(new_n411_), .ZN(new_n412_));
  AOI22_X1  g211(.A1(new_n391_), .A2(new_n393_), .B1(new_n397_), .B2(KEYINPUT8), .ZN(new_n413_));
  INV_X1    g212(.A(new_n406_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n410_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  XOR2_X1   g216(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n418_));
  NAND2_X1  g217(.A1(G232gat), .A2(G233gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  OR2_X1    g219(.A1(new_n420_), .A2(KEYINPUT35), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n412_), .A2(new_n417_), .A3(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n420_), .A2(KEYINPUT35), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n412_), .A2(new_n417_), .A3(new_n423_), .A4(new_n421_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(new_n426_), .A3(KEYINPUT71), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G190gat), .B(G218gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G134gat), .B(G162gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n428_), .B(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n430_), .A2(KEYINPUT36), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n427_), .A2(new_n432_), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n425_), .A2(new_n426_), .A3(KEYINPUT71), .A4(new_n431_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n425_), .A2(new_n426_), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n430_), .A2(KEYINPUT36), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n435_), .A2(new_n438_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n371_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT13), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G230gat), .A2(G233gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G57gat), .B(G64gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT11), .ZN(new_n444_));
  XNOR2_X1  g243(.A(KEYINPUT66), .B(G71gat), .ZN(new_n445_));
  INV_X1    g244(.A(G78gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n445_), .B(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n444_), .A2(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n445_), .B(G78gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n443_), .A2(KEYINPUT11), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n448_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n399_), .A2(new_n453_), .A3(new_n406_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n452_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n442_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  OR2_X1    g255(.A1(new_n456_), .A2(KEYINPUT67), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(KEYINPUT67), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n453_), .B1(new_n399_), .B2(new_n406_), .ZN(new_n460_));
  NOR3_X1   g259(.A1(new_n413_), .A2(new_n414_), .A3(new_n452_), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT12), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT12), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n463_), .B1(new_n415_), .B2(new_n453_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n462_), .A2(new_n442_), .A3(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(KEYINPUT69), .B1(new_n459_), .B2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G120gat), .B(G148gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(KEYINPUT5), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G176gat), .B(G204gat), .ZN(new_n470_));
  XOR2_X1   g269(.A(new_n469_), .B(new_n470_), .Z(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n472_), .A2(KEYINPUT68), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT69), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n457_), .A2(new_n465_), .A3(new_n474_), .A4(new_n458_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n467_), .A2(new_n473_), .A3(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n473_), .B1(new_n467_), .B2(new_n475_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n441_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n478_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n480_), .A2(KEYINPUT13), .A3(new_n476_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G15gat), .B(G22gat), .ZN(new_n484_));
  INV_X1    g283(.A(G1gat), .ZN(new_n485_));
  INV_X1    g284(.A(G8gat), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT14), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n484_), .A2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G1gat), .B(G8gat), .ZN(new_n489_));
  XOR2_X1   g288(.A(new_n488_), .B(new_n489_), .Z(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(new_n416_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT77), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n488_), .B(new_n489_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(new_n410_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n491_), .A2(new_n492_), .A3(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G229gat), .A2(G233gat), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n493_), .A2(KEYINPUT77), .A3(new_n410_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n495_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT78), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT78), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n495_), .A2(new_n501_), .A3(new_n497_), .A4(new_n498_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n500_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n411_), .A2(new_n493_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n496_), .B(KEYINPUT79), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n504_), .A2(new_n491_), .A3(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G113gat), .B(G141gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G169gat), .B(G197gat), .ZN(new_n508_));
  XOR2_X1   g307(.A(new_n507_), .B(new_n508_), .Z(new_n509_));
  AND3_X1   g308(.A1(new_n503_), .A2(new_n506_), .A3(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n509_), .B1(new_n503_), .B2(new_n506_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n512_), .A2(KEYINPUT80), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT80), .ZN(new_n514_));
  NOR3_X1   g313(.A1(new_n510_), .A2(new_n511_), .A3(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  XOR2_X1   g315(.A(G127gat), .B(G155gat), .Z(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT16), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G183gat), .B(G211gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT17), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT76), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G231gat), .A2(G233gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n493_), .B(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(new_n452_), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n525_), .A2(KEYINPUT75), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n525_), .A2(KEYINPUT75), .ZN(new_n527_));
  NOR3_X1   g326(.A1(new_n522_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n528_));
  OR2_X1    g327(.A1(new_n525_), .A2(KEYINPUT73), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n525_), .A2(KEYINPUT73), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT17), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n520_), .A2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n529_), .A2(new_n530_), .A3(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT74), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n534_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n528_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NOR3_X1   g337(.A1(new_n483_), .A2(new_n516_), .A3(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT100), .ZN(new_n540_));
  OR2_X1    g339(.A1(new_n539_), .A2(KEYINPUT100), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n440_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  OAI21_X1  g341(.A(G1gat), .B1(new_n542_), .B2(new_n329_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n371_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n516_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT72), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n439_), .A2(new_n548_), .A3(KEYINPUT37), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT37), .ZN(new_n550_));
  AOI22_X1  g349(.A1(new_n433_), .A2(new_n434_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n550_), .B1(new_n551_), .B2(KEYINPUT72), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n549_), .A2(new_n552_), .A3(new_n537_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n553_), .B1(new_n481_), .B2(new_n479_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n547_), .A2(new_n554_), .ZN(new_n555_));
  NOR3_X1   g354(.A1(new_n555_), .A2(G1gat), .A3(new_n329_), .ZN(new_n556_));
  AND3_X1   g355(.A1(new_n556_), .A2(KEYINPUT99), .A3(KEYINPUT38), .ZN(new_n557_));
  AOI21_X1  g356(.A(KEYINPUT99), .B1(new_n556_), .B2(KEYINPUT38), .ZN(new_n558_));
  OAI221_X1 g357(.A(new_n543_), .B1(KEYINPUT38), .B2(new_n556_), .C1(new_n557_), .C2(new_n558_), .ZN(G1324gat));
  INV_X1    g358(.A(KEYINPUT40), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT101), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n440_), .A2(new_n366_), .A3(new_n540_), .A4(new_n541_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n561_), .B1(new_n562_), .B2(G8gat), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n562_), .A2(new_n561_), .A3(G8gat), .ZN(new_n565_));
  AND3_X1   g364(.A1(new_n564_), .A2(KEYINPUT39), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT39), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n563_), .A2(new_n567_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n547_), .A2(new_n486_), .A3(new_n366_), .A4(new_n554_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n560_), .B1(new_n566_), .B2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n564_), .A2(KEYINPUT39), .A3(new_n565_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n572_), .A2(KEYINPUT40), .A3(new_n568_), .A4(new_n569_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n571_), .A2(new_n573_), .ZN(G1325gat));
  OAI21_X1  g373(.A(G15gat), .B1(new_n542_), .B2(new_n368_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(KEYINPUT102), .B(KEYINPUT41), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  OR3_X1    g376(.A1(new_n555_), .A2(G15gat), .A3(new_n368_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n575_), .A2(new_n576_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n577_), .A2(new_n578_), .A3(new_n579_), .ZN(G1326gat));
  XOR2_X1   g379(.A(new_n356_), .B(KEYINPUT103), .Z(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  OR3_X1    g381(.A1(new_n555_), .A2(G22gat), .A3(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(G22gat), .B1(new_n542_), .B2(new_n582_), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n584_), .A2(KEYINPUT42), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n584_), .A2(KEYINPUT42), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n583_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT104), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  OAI211_X1 g388(.A(new_n583_), .B(KEYINPUT104), .C1(new_n585_), .C2(new_n586_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(G1327gat));
  NAND2_X1  g390(.A1(new_n549_), .A2(new_n552_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n592_), .B1(new_n365_), .B2(new_n370_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT43), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n537_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n483_), .A2(new_n516_), .ZN(new_n596_));
  OAI211_X1 g395(.A(KEYINPUT43), .B(new_n592_), .C1(new_n365_), .C2(new_n370_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n595_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n598_));
  XOR2_X1   g397(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n595_), .A2(KEYINPUT44), .A3(new_n596_), .A4(new_n597_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n600_), .A2(new_n328_), .A3(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(G29gat), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n538_), .A2(new_n439_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n483_), .A2(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n544_), .A2(new_n545_), .A3(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n329_), .A2(G29gat), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n607_), .B(KEYINPUT106), .Z(new_n608_));
  OAI21_X1  g407(.A(new_n603_), .B1(new_n606_), .B2(new_n608_), .ZN(G1328gat));
  NAND3_X1  g408(.A1(new_n600_), .A2(new_n366_), .A3(new_n601_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(G36gat), .ZN(new_n611_));
  INV_X1    g410(.A(new_n366_), .ZN(new_n612_));
  OR2_X1    g411(.A1(new_n612_), .A2(G36gat), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n606_), .A2(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n611_), .A2(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(KEYINPUT108), .B(KEYINPUT46), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n611_), .A2(new_n616_), .A3(new_n618_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(G1329gat));
  NAND4_X1  g421(.A1(new_n600_), .A2(G43gat), .A3(new_n242_), .A4(new_n601_), .ZN(new_n623_));
  INV_X1    g422(.A(G43gat), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n624_), .B1(new_n606_), .B2(new_n368_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(G1330gat));
  NAND4_X1  g427(.A1(new_n600_), .A2(G50gat), .A3(new_n359_), .A4(new_n601_), .ZN(new_n629_));
  INV_X1    g428(.A(G50gat), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n630_), .B1(new_n606_), .B2(new_n582_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n629_), .A2(new_n631_), .ZN(G1331gat));
  NOR2_X1   g431(.A1(new_n482_), .A2(new_n545_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n544_), .A2(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n634_), .A2(new_n553_), .ZN(new_n635_));
  INV_X1    g434(.A(G57gat), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n635_), .A2(new_n636_), .A3(new_n328_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n440_), .A2(new_n537_), .A3(new_n633_), .ZN(new_n638_));
  OAI21_X1  g437(.A(G57gat), .B1(new_n638_), .B2(new_n329_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(G1332gat));
  OAI21_X1  g439(.A(G64gat), .B1(new_n638_), .B2(new_n612_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT48), .ZN(new_n642_));
  INV_X1    g441(.A(G64gat), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n635_), .A2(new_n643_), .A3(new_n366_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n644_), .ZN(G1333gat));
  INV_X1    g444(.A(G71gat), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n635_), .A2(new_n646_), .A3(new_n242_), .ZN(new_n647_));
  OAI21_X1  g446(.A(G71gat), .B1(new_n638_), .B2(new_n368_), .ZN(new_n648_));
  OR2_X1    g447(.A1(new_n648_), .A2(KEYINPUT111), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(KEYINPUT111), .ZN(new_n650_));
  XNOR2_X1  g449(.A(KEYINPUT110), .B(KEYINPUT49), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n649_), .A2(new_n650_), .A3(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n651_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n647_), .B1(new_n652_), .B2(new_n653_), .ZN(G1334gat));
  OAI21_X1  g453(.A(G78gat), .B1(new_n638_), .B2(new_n582_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT50), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n635_), .A2(new_n446_), .A3(new_n581_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(G1335gat));
  NOR2_X1   g457(.A1(new_n634_), .A2(new_n604_), .ZN(new_n659_));
  INV_X1    g458(.A(G85gat), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n659_), .A2(new_n660_), .A3(new_n328_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n595_), .A2(new_n597_), .A3(new_n633_), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n662_), .A2(KEYINPUT112), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(KEYINPUT112), .ZN(new_n664_));
  AND3_X1   g463(.A1(new_n663_), .A2(new_n328_), .A3(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n661_), .B1(new_n665_), .B2(new_n660_), .ZN(G1336gat));
  INV_X1    g465(.A(G92gat), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n659_), .A2(new_n667_), .A3(new_n366_), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n663_), .A2(new_n366_), .A3(new_n664_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n668_), .B1(new_n669_), .B2(new_n667_), .ZN(G1337gat));
  OAI21_X1  g469(.A(G99gat), .B1(new_n662_), .B2(new_n368_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n368_), .A2(new_n403_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n659_), .A2(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n671_), .A2(KEYINPUT113), .A3(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n674_), .B(new_n675_), .ZN(G1338gat));
  INV_X1    g475(.A(G106gat), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n659_), .A2(new_n677_), .A3(new_n359_), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n595_), .A2(new_n359_), .A3(new_n597_), .A4(new_n633_), .ZN(new_n679_));
  XOR2_X1   g478(.A(KEYINPUT115), .B(KEYINPUT52), .Z(new_n680_));
  NAND3_X1  g479(.A1(new_n679_), .A2(G106gat), .A3(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n680_), .B1(new_n679_), .B2(G106gat), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n678_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(new_n687_));
  OAI211_X1 g486(.A(new_n678_), .B(new_n685_), .C1(new_n682_), .C2(new_n683_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1339gat));
  INV_X1    g488(.A(KEYINPUT121), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n367_), .A2(new_n328_), .A3(new_n242_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT120), .ZN(new_n693_));
  INV_X1    g492(.A(new_n442_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n463_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n695_));
  AOI21_X1  g494(.A(KEYINPUT12), .B1(new_n407_), .B2(new_n452_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n694_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n465_), .A2(new_n697_), .A3(KEYINPUT55), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT55), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n462_), .A2(new_n699_), .A3(new_n442_), .A4(new_n464_), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n698_), .A2(KEYINPUT118), .A3(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(KEYINPUT118), .B1(new_n698_), .B2(new_n700_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n471_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT56), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  OAI211_X1 g504(.A(KEYINPUT56), .B(new_n471_), .C1(new_n701_), .C2(new_n702_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NOR3_X1   g506(.A1(new_n459_), .A2(new_n466_), .A3(new_n471_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n709_), .B1(new_n513_), .B2(new_n515_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n707_), .A2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT119), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n710_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT119), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n505_), .B1(new_n490_), .B2(new_n416_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n509_), .B1(new_n504_), .B2(new_n717_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n495_), .A2(new_n498_), .A3(new_n505_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  OR2_X1    g519(.A1(new_n510_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n480_), .A2(new_n476_), .A3(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n713_), .A2(new_n716_), .A3(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT57), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n439_), .A2(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n693_), .B1(new_n724_), .B2(new_n726_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n723_), .B1(new_n714_), .B2(new_n715_), .ZN(new_n728_));
  AOI211_X1 g527(.A(KEYINPUT119), .B(new_n710_), .C1(new_n705_), .C2(new_n706_), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n693_), .B(new_n726_), .C1(new_n728_), .C2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n727_), .A2(new_n731_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n551_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n733_));
  AOI211_X1 g532(.A(new_n708_), .B(new_n721_), .C1(new_n705_), .C2(new_n706_), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n734_), .A2(KEYINPUT58), .ZN(new_n735_));
  INV_X1    g534(.A(new_n592_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n736_), .B1(new_n734_), .B2(KEYINPUT58), .ZN(new_n737_));
  AOI22_X1  g536(.A1(new_n733_), .A2(new_n725_), .B1(new_n735_), .B2(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n537_), .B1(new_n732_), .B2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT54), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT117), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n741_), .B1(new_n554_), .B2(new_n516_), .ZN(new_n742_));
  AND3_X1   g541(.A1(new_n549_), .A2(new_n552_), .A3(new_n537_), .ZN(new_n743_));
  AND4_X1   g542(.A1(new_n741_), .A2(new_n482_), .A3(new_n743_), .A4(new_n516_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n740_), .B1(new_n742_), .B2(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n554_), .A2(new_n741_), .A3(new_n516_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n482_), .A2(new_n743_), .A3(new_n516_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(KEYINPUT117), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n746_), .A2(new_n748_), .A3(KEYINPUT54), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n745_), .A2(new_n749_), .ZN(new_n750_));
  OAI211_X1 g549(.A(new_n690_), .B(new_n692_), .C1(new_n739_), .C2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n733_), .A2(new_n725_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n726_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(KEYINPUT120), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n735_), .A2(new_n737_), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n752_), .A2(new_n754_), .A3(new_n755_), .A4(new_n730_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n750_), .B1(new_n756_), .B2(new_n538_), .ZN(new_n757_));
  OAI21_X1  g556(.A(KEYINPUT121), .B1(new_n757_), .B2(new_n691_), .ZN(new_n758_));
  INV_X1    g557(.A(G113gat), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n751_), .A2(new_n758_), .A3(new_n759_), .A4(new_n545_), .ZN(new_n760_));
  OAI211_X1 g559(.A(KEYINPUT59), .B(new_n692_), .C1(new_n739_), .C2(new_n750_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT59), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n762_), .B1(new_n757_), .B2(new_n691_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n516_), .B1(new_n761_), .B2(new_n763_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n760_), .B1(new_n764_), .B2(new_n759_), .ZN(G1340gat));
  INV_X1    g564(.A(G120gat), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n766_), .B1(new_n482_), .B2(KEYINPUT60), .ZN(new_n767_));
  OR2_X1    g566(.A1(new_n766_), .A2(KEYINPUT60), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n751_), .A2(new_n758_), .A3(new_n767_), .A4(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n482_), .B1(new_n761_), .B2(new_n763_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n769_), .B1(new_n770_), .B2(new_n766_), .ZN(G1341gat));
  INV_X1    g570(.A(KEYINPUT122), .ZN(new_n772_));
  INV_X1    g571(.A(G127gat), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n761_), .A2(new_n763_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n773_), .B1(new_n774_), .B2(new_n537_), .ZN(new_n775_));
  AND4_X1   g574(.A1(new_n773_), .A2(new_n751_), .A3(new_n758_), .A4(new_n537_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n772_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n751_), .A2(new_n758_), .A3(new_n773_), .A4(new_n537_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n538_), .B1(new_n761_), .B2(new_n763_), .ZN(new_n779_));
  OAI211_X1 g578(.A(KEYINPUT122), .B(new_n778_), .C1(new_n779_), .C2(new_n773_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n777_), .A2(new_n780_), .ZN(G1342gat));
  INV_X1    g580(.A(G134gat), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n751_), .A2(new_n758_), .A3(new_n782_), .A4(new_n439_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n736_), .B1(new_n761_), .B2(new_n763_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n783_), .B1(new_n784_), .B2(new_n782_), .ZN(G1343gat));
  INV_X1    g584(.A(new_n757_), .ZN(new_n786_));
  NOR3_X1   g585(.A1(new_n329_), .A2(new_n356_), .A3(new_n242_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n786_), .A2(new_n612_), .A3(new_n787_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n788_), .A2(new_n516_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(KEYINPUT123), .B(G141gat), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n789_), .B(new_n790_), .ZN(G1344gat));
  NOR2_X1   g590(.A1(new_n788_), .A2(new_n482_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(KEYINPUT124), .B(G148gat), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n792_), .B(new_n793_), .ZN(G1345gat));
  NOR2_X1   g593(.A1(new_n788_), .A2(new_n538_), .ZN(new_n795_));
  XOR2_X1   g594(.A(KEYINPUT61), .B(G155gat), .Z(new_n796_));
  XNOR2_X1  g595(.A(new_n795_), .B(new_n796_), .ZN(G1346gat));
  OAI21_X1  g596(.A(G162gat), .B1(new_n788_), .B2(new_n736_), .ZN(new_n798_));
  OR2_X1    g597(.A1(new_n551_), .A2(G162gat), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n798_), .B1(new_n788_), .B2(new_n799_), .ZN(G1347gat));
  INV_X1    g599(.A(KEYINPUT62), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n366_), .A2(new_n369_), .ZN(new_n802_));
  NOR3_X1   g601(.A1(new_n757_), .A2(new_n581_), .A3(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n804_), .A2(new_n516_), .ZN(new_n805_));
  INV_X1    g604(.A(G169gat), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n801_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n805_), .A2(new_n202_), .ZN(new_n808_));
  OAI211_X1 g607(.A(KEYINPUT62), .B(G169gat), .C1(new_n804_), .C2(new_n516_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n807_), .A2(new_n808_), .A3(new_n809_), .ZN(G1348gat));
  AOI21_X1  g609(.A(G176gat), .B1(new_n803_), .B2(new_n483_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n757_), .A2(new_n359_), .ZN(new_n812_));
  NOR3_X1   g611(.A1(new_n482_), .A2(new_n802_), .A3(new_n203_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n811_), .B1(new_n812_), .B2(new_n813_), .ZN(G1349gat));
  NAND4_X1  g613(.A1(new_n812_), .A2(new_n366_), .A3(new_n369_), .A4(new_n537_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n538_), .A2(new_n286_), .ZN(new_n816_));
  AOI22_X1  g615(.A1(new_n815_), .A2(new_n209_), .B1(new_n803_), .B2(new_n816_), .ZN(G1350gat));
  OAI21_X1  g616(.A(G190gat), .B1(new_n804_), .B2(new_n736_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n803_), .A2(new_n225_), .A3(new_n439_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(G1351gat));
  NAND3_X1  g619(.A1(new_n329_), .A2(new_n359_), .A3(new_n368_), .ZN(new_n821_));
  NOR3_X1   g620(.A1(new_n757_), .A2(new_n612_), .A3(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n545_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n823_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g623(.A1(new_n822_), .A2(new_n483_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n825_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g625(.A(new_n538_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n822_), .A2(new_n827_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(KEYINPUT125), .B(KEYINPUT126), .ZN(new_n829_));
  NOR2_X1   g628(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n829_), .B(new_n830_), .ZN(new_n831_));
  XOR2_X1   g630(.A(new_n828_), .B(new_n831_), .Z(G1354gat));
  AOI21_X1  g631(.A(G218gat), .B1(new_n822_), .B2(new_n439_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n592_), .A2(G218gat), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(KEYINPUT127), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n833_), .B1(new_n822_), .B2(new_n835_), .ZN(G1355gat));
endmodule


