//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 1 0 1 1 0 1 0 0 0 0 0 1 0 1 1 0 1 0 1 1 1 0 0 0 1 1 1 1 1 1 1 0 0 1 0 0 1 1 0 0 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n769_, new_n770_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n791_, new_n792_, new_n793_,
    new_n795_, new_n796_, new_n797_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n808_,
    new_n809_, new_n811_, new_n812_, new_n813_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n915_, new_n917_, new_n918_, new_n920_,
    new_n921_, new_n922_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n949_, new_n950_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n957_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n966_, new_n967_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G57gat), .B(G64gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT11), .ZN(new_n204_));
  XOR2_X1   g003(.A(G71gat), .B(G78gat), .Z(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n203_), .A2(KEYINPUT11), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n204_), .A2(new_n205_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n211_));
  OR3_X1    g010(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G99gat), .A2(G106gat), .ZN(new_n213_));
  AND2_X1   g012(.A1(new_n213_), .A2(KEYINPUT6), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n213_), .A2(KEYINPUT6), .ZN(new_n215_));
  OAI211_X1 g014(.A(new_n211_), .B(new_n212_), .C1(new_n214_), .C2(new_n215_), .ZN(new_n216_));
  XOR2_X1   g015(.A(G85gat), .B(G92gat), .Z(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT8), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT8), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n216_), .A2(new_n220_), .A3(new_n217_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n219_), .A2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n213_), .B(KEYINPUT6), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT10), .B(G99gat), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n223_), .B1(G106gat), .B2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(G85gat), .ZN(new_n227_));
  INV_X1    g026(.A(G92gat), .ZN(new_n228_));
  OR3_X1    g027(.A1(new_n227_), .A2(new_n228_), .A3(KEYINPUT9), .ZN(new_n229_));
  XOR2_X1   g028(.A(KEYINPUT64), .B(KEYINPUT9), .Z(new_n230_));
  XNOR2_X1  g029(.A(G85gat), .B(G92gat), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n229_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n232_), .A2(KEYINPUT65), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT65), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n217_), .A2(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n234_), .B1(new_n236_), .B2(new_n229_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n226_), .B1(new_n233_), .B2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n222_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n232_), .A2(KEYINPUT65), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n236_), .A2(new_n234_), .A3(new_n229_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n225_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n243_), .A2(KEYINPUT66), .ZN(new_n244_));
  OAI211_X1 g043(.A(KEYINPUT12), .B(new_n210_), .C1(new_n240_), .C2(new_n244_), .ZN(new_n245_));
  AND2_X1   g044(.A1(G230gat), .A2(G233gat), .ZN(new_n246_));
  AND3_X1   g045(.A1(new_n216_), .A2(new_n220_), .A3(new_n217_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n220_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n249_), .A2(new_n243_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n209_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n251_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n246_), .B1(new_n250_), .B2(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n252_), .B1(new_n238_), .B2(new_n222_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT67), .ZN(new_n255_));
  NOR3_X1   g054(.A1(new_n254_), .A2(new_n255_), .A3(KEYINPUT12), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n210_), .B1(new_n249_), .B2(new_n243_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT12), .ZN(new_n258_));
  AOI21_X1  g057(.A(KEYINPUT67), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  OAI211_X1 g058(.A(new_n245_), .B(new_n253_), .C1(new_n256_), .C2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n250_), .A2(new_n252_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(new_n257_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(new_n246_), .ZN(new_n263_));
  AND2_X1   g062(.A1(new_n260_), .A2(new_n263_), .ZN(new_n264_));
  XOR2_X1   g063(.A(G120gat), .B(G148gat), .Z(new_n265_));
  XNOR2_X1  g064(.A(G176gat), .B(G204gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n268_));
  XOR2_X1   g067(.A(new_n267_), .B(new_n268_), .Z(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  AND2_X1   g069(.A1(new_n264_), .A2(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n264_), .A2(new_n270_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT13), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT13), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n275_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n274_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G29gat), .B(G36gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT71), .ZN(new_n280_));
  XOR2_X1   g079(.A(G43gat), .B(G50gat), .Z(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT15), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G15gat), .B(G22gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(KEYINPUT72), .ZN(new_n286_));
  INV_X1    g085(.A(G8gat), .ZN(new_n287_));
  OAI21_X1  g086(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT73), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n286_), .A2(new_n289_), .ZN(new_n290_));
  XOR2_X1   g089(.A(G1gat), .B(G8gat), .Z(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  OR2_X1    g091(.A1(new_n284_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n282_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G229gat), .A2(G233gat), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n293_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n292_), .B(new_n282_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n295_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G113gat), .B(G141gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT77), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G169gat), .B(G197gat), .ZN(new_n302_));
  XOR2_X1   g101(.A(new_n301_), .B(new_n302_), .Z(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n296_), .A2(new_n299_), .A3(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n304_), .B1(new_n296_), .B2(new_n299_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n278_), .A2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G127gat), .B(G155gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G183gat), .B(G211gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  XOR2_X1   g112(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT75), .B(KEYINPUT17), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n317_), .B(KEYINPUT76), .Z(new_n318_));
  XNOR2_X1  g117(.A(new_n292_), .B(new_n252_), .ZN(new_n319_));
  AND2_X1   g118(.A1(G231gat), .A2(G233gat), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  OR2_X1    g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n319_), .A2(new_n321_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n318_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  AND2_X1   g123(.A1(new_n322_), .A2(new_n323_), .ZN(new_n325_));
  XOR2_X1   g124(.A(new_n315_), .B(KEYINPUT17), .Z(new_n326_));
  AOI21_X1  g125(.A(new_n324_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n310_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G183gat), .A2(G190gat), .ZN(new_n330_));
  AND2_X1   g129(.A1(KEYINPUT83), .A2(KEYINPUT23), .ZN(new_n331_));
  NOR2_X1   g130(.A1(KEYINPUT83), .A2(KEYINPUT23), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n330_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n330_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT23), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n333_), .A2(new_n336_), .ZN(new_n337_));
  NOR3_X1   g136(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G169gat), .A2(G176gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT82), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT82), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n341_), .A2(G169gat), .A3(G176gat), .ZN(new_n342_));
  AND2_X1   g141(.A1(new_n340_), .A2(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n338_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n346_));
  AND2_X1   g145(.A1(KEYINPUT79), .A2(KEYINPUT25), .ZN(new_n347_));
  NOR2_X1   g146(.A1(KEYINPUT79), .A2(KEYINPUT25), .ZN(new_n348_));
  OAI21_X1  g147(.A(G183gat), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT80), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT80), .ZN(new_n351_));
  OAI211_X1 g150(.A(new_n351_), .B(G183gat), .C1(new_n347_), .C2(new_n348_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(G183gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(KEYINPUT25), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT26), .ZN(new_n356_));
  OR2_X1    g155(.A1(KEYINPUT81), .A2(G190gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(KEYINPUT81), .A2(G190gat), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n356_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n355_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  OAI211_X1 g160(.A(new_n337_), .B(new_n346_), .C1(new_n353_), .C2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT83), .B(KEYINPUT23), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(new_n334_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n330_), .A2(new_n335_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n357_), .A2(new_n354_), .A3(new_n358_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n364_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(G169gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT22), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT22), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(G169gat), .ZN(new_n371_));
  INV_X1    g170(.A(G176gat), .ZN(new_n372_));
  AND3_X1   g171(.A1(new_n369_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n367_), .A2(new_n343_), .A3(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n362_), .A2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT30), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G227gat), .A2(G233gat), .ZN(new_n378_));
  XOR2_X1   g177(.A(new_n378_), .B(G15gat), .Z(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(G71gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(G99gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n377_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT30), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n376_), .B(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n381_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n382_), .A2(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G127gat), .B(G134gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G113gat), .B(G120gat), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n388_), .A2(new_n389_), .A3(KEYINPUT85), .ZN(new_n390_));
  OR2_X1    g189(.A1(new_n388_), .A2(new_n389_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT85), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n388_), .A2(new_n389_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n391_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n387_), .A2(new_n390_), .A3(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(KEYINPUT84), .B(G43gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT31), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n394_), .A2(new_n390_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n382_), .A2(new_n386_), .A3(new_n398_), .ZN(new_n399_));
  AND3_X1   g198(.A1(new_n395_), .A2(new_n397_), .A3(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n397_), .B1(new_n395_), .B2(new_n399_), .ZN(new_n401_));
  OR2_X1    g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G78gat), .B(G106gat), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT93), .ZN(new_n404_));
  AND2_X1   g203(.A1(G228gat), .A2(G233gat), .ZN(new_n405_));
  INV_X1    g204(.A(G218gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(G211gat), .ZN(new_n407_));
  INV_X1    g206(.A(G211gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(G218gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(G197gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(G204gat), .ZN(new_n412_));
  INV_X1    g211(.A(G204gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(G197gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n410_), .B1(KEYINPUT21), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT90), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n412_), .A2(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n411_), .A2(KEYINPUT90), .A3(G204gat), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT21), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n418_), .A2(new_n419_), .A3(new_n420_), .A4(new_n414_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n418_), .A2(new_n414_), .A3(new_n419_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n420_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n423_));
  AOI22_X1  g222(.A1(new_n416_), .A2(new_n421_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT29), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G155gat), .A2(G162gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT1), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT1), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n429_), .A2(G155gat), .A3(G162gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n428_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT87), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT86), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT86), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT87), .ZN(new_n436_));
  NOR2_X1   g235(.A1(G155gat), .A2(G162gat), .ZN(new_n437_));
  AND3_X1   g236(.A1(new_n434_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n437_), .B1(new_n434_), .B2(new_n436_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n432_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G141gat), .A2(G148gat), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(G141gat), .A2(G148gat), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n440_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT3), .ZN(new_n446_));
  INV_X1    g245(.A(G141gat), .ZN(new_n447_));
  INV_X1    g246(.A(G148gat), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n446_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT2), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n441_), .A2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n449_), .A2(new_n451_), .A3(new_n452_), .A4(new_n453_), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n454_), .B(new_n427_), .C1(new_n438_), .C2(new_n439_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n426_), .B1(new_n445_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT92), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n425_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n437_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n435_), .A2(KEYINPUT87), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n433_), .A2(KEYINPUT86), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n459_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n434_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n431_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n444_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n455_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT29), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n467_), .A2(KEYINPUT92), .ZN(new_n468_));
  OAI211_X1 g267(.A(new_n404_), .B(new_n405_), .C1(new_n458_), .C2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT88), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n466_), .A2(new_n470_), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n455_), .B(KEYINPUT88), .C1(new_n464_), .C2(new_n465_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n471_), .A2(KEYINPUT29), .A3(new_n472_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n424_), .A2(new_n405_), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n473_), .A2(KEYINPUT91), .A3(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(KEYINPUT91), .B1(new_n473_), .B2(new_n474_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n469_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n424_), .B1(new_n467_), .B2(KEYINPUT92), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n478_), .B1(KEYINPUT92), .B2(new_n467_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n404_), .B1(new_n479_), .B2(new_n405_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n403_), .B1(new_n477_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n473_), .A2(new_n474_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT91), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n473_), .A2(KEYINPUT91), .A3(new_n474_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n405_), .B1(new_n458_), .B2(new_n468_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT93), .ZN(new_n488_));
  INV_X1    g287(.A(new_n403_), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n486_), .A2(new_n488_), .A3(new_n489_), .A4(new_n469_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n481_), .A2(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n486_), .A2(new_n488_), .A3(new_n469_), .ZN(new_n492_));
  AOI21_X1  g291(.A(KEYINPUT94), .B1(new_n492_), .B2(new_n403_), .ZN(new_n493_));
  XOR2_X1   g292(.A(G22gat), .B(G50gat), .Z(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT89), .B(KEYINPUT28), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n471_), .A2(new_n472_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n496_), .B1(new_n497_), .B2(new_n426_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n497_), .A2(new_n426_), .A3(new_n496_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n494_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n500_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n494_), .ZN(new_n503_));
  NOR3_X1   g302(.A1(new_n502_), .A2(new_n498_), .A3(new_n503_), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n501_), .A2(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n491_), .B1(new_n493_), .B2(new_n505_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n501_), .A2(new_n504_), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n507_), .A2(new_n481_), .A3(KEYINPUT94), .A4(new_n490_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G225gat), .A2(G233gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT101), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n471_), .A2(new_n472_), .A3(new_n398_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT4), .ZN(new_n512_));
  AND2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n391_), .A2(new_n393_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n445_), .A2(new_n455_), .A3(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n512_), .B1(new_n511_), .B2(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n510_), .B1(new_n513_), .B2(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n511_), .A2(new_n515_), .A3(new_n509_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G1gat), .B(G29gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(G85gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(KEYINPUT0), .B(G57gat), .ZN(new_n521_));
  XOR2_X1   g320(.A(new_n520_), .B(new_n521_), .Z(new_n522_));
  AND3_X1   g321(.A1(new_n517_), .A2(new_n518_), .A3(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n522_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n524_));
  OAI21_X1  g323(.A(KEYINPUT103), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n524_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT103), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n517_), .A2(new_n518_), .A3(new_n522_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n526_), .A2(new_n527_), .A3(new_n528_), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n506_), .A2(new_n508_), .A3(new_n525_), .A4(new_n529_), .ZN(new_n530_));
  XOR2_X1   g329(.A(G8gat), .B(G36gat), .Z(new_n531_));
  XNOR2_X1  g330(.A(KEYINPUT100), .B(KEYINPUT18), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G64gat), .B(G92gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n330_), .A2(KEYINPUT23), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n537_), .B1(new_n363_), .B2(new_n330_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(G183gat), .A2(G190gat), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n374_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n340_), .A2(new_n342_), .A3(KEYINPUT97), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(KEYINPUT97), .B1(new_n340_), .B2(new_n342_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(KEYINPUT98), .B1(new_n540_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n539_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n373_), .B1(new_n337_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT98), .ZN(new_n548_));
  INV_X1    g347(.A(new_n543_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(new_n541_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n547_), .A2(new_n548_), .A3(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n545_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n338_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n364_), .A2(new_n553_), .A3(new_n365_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(KEYINPUT96), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT96), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n364_), .A2(new_n556_), .A3(new_n553_), .A4(new_n365_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n345_), .A2(new_n339_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(KEYINPUT26), .B(G190gat), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT25), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(G183gat), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n355_), .A2(new_n561_), .A3(KEYINPUT95), .ZN(new_n562_));
  AOI21_X1  g361(.A(KEYINPUT95), .B1(new_n355_), .B2(new_n561_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n559_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n555_), .A2(new_n557_), .A3(new_n558_), .A4(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n424_), .B1(new_n552_), .B2(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(KEYINPUT20), .B1(new_n376_), .B2(new_n425_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G226gat), .A2(G233gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT19), .ZN(new_n569_));
  NOR3_X1   g368(.A1(new_n566_), .A2(new_n567_), .A3(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n569_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n424_), .B1(new_n362_), .B2(new_n375_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT20), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  OAI211_X1 g373(.A(new_n565_), .B(new_n424_), .C1(new_n544_), .C2(new_n540_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n571_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n536_), .B1(new_n570_), .B2(new_n576_), .ZN(new_n577_));
  NOR3_X1   g376(.A1(new_n540_), .A2(new_n544_), .A3(KEYINPUT98), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n548_), .B1(new_n547_), .B2(new_n550_), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n565_), .B(new_n424_), .C1(new_n578_), .C2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT99), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NOR3_X1   g381(.A1(new_n572_), .A2(new_n573_), .A3(new_n569_), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n552_), .A2(KEYINPUT99), .A3(new_n424_), .A4(new_n565_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n582_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n569_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n585_), .A2(new_n586_), .A3(new_n535_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n577_), .A2(new_n587_), .A3(KEYINPUT27), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n585_), .A2(new_n586_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(new_n536_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(new_n587_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT27), .ZN(new_n592_));
  AOI21_X1  g391(.A(KEYINPUT104), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  AND3_X1   g392(.A1(new_n585_), .A2(new_n586_), .A3(new_n535_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n535_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n595_));
  OAI211_X1 g394(.A(KEYINPUT104), .B(new_n592_), .C1(new_n594_), .C2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n588_), .B1(new_n593_), .B2(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n530_), .A2(new_n598_), .ZN(new_n599_));
  OAI21_X1  g398(.A(KEYINPUT102), .B1(new_n523_), .B2(KEYINPUT33), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n509_), .B1(new_n513_), .B2(new_n516_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n522_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n511_), .A2(new_n515_), .A3(new_n510_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n601_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  AND3_X1   g403(.A1(new_n604_), .A2(new_n590_), .A3(new_n587_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n523_), .A2(KEYINPUT33), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT102), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT33), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n528_), .A2(new_n607_), .A3(new_n608_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n600_), .A2(new_n605_), .A3(new_n606_), .A4(new_n609_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n535_), .A2(KEYINPUT32), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n611_), .B1(new_n570_), .B2(new_n576_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n612_), .B1(new_n589_), .B2(new_n611_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n613_), .B1(new_n526_), .B2(new_n528_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  AOI22_X1  g414(.A1(new_n610_), .A2(new_n615_), .B1(new_n508_), .B2(new_n506_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n402_), .B1(new_n599_), .B2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n529_), .A2(new_n525_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n402_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT94), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n481_), .A2(new_n620_), .ZN(new_n621_));
  AOI22_X1  g420(.A1(new_n621_), .A2(new_n507_), .B1(new_n481_), .B2(new_n490_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n508_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n588_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n592_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT104), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n626_), .B1(new_n629_), .B2(new_n596_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT105), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  AOI211_X1 g431(.A(KEYINPUT105), .B(new_n626_), .C1(new_n629_), .C2(new_n596_), .ZN(new_n633_));
  OAI211_X1 g432(.A(new_n619_), .B(new_n625_), .C1(new_n632_), .C2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n617_), .A2(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n240_), .A2(new_n244_), .ZN(new_n636_));
  OR2_X1    g435(.A1(new_n284_), .A2(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n638_));
  NAND2_X1  g437(.A1(G232gat), .A2(G233gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n638_), .B(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT35), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n642_), .B(KEYINPUT70), .Z(new_n643_));
  AOI22_X1  g442(.A1(new_n250_), .A2(new_n282_), .B1(new_n641_), .B2(new_n640_), .ZN(new_n644_));
  AND3_X1   g443(.A1(new_n637_), .A2(new_n643_), .A3(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n643_), .B1(new_n637_), .B2(new_n644_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(G190gat), .B(G218gat), .ZN(new_n647_));
  XNOR2_X1  g446(.A(G134gat), .B(G162gat), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n647_), .B(new_n648_), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n649_), .A2(KEYINPUT36), .ZN(new_n650_));
  OR3_X1    g449(.A1(new_n645_), .A2(new_n646_), .A3(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n649_), .A2(KEYINPUT36), .ZN(new_n652_));
  OAI211_X1 g451(.A(new_n650_), .B(new_n652_), .C1(new_n645_), .C2(new_n646_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n329_), .A2(new_n635_), .A3(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n202_), .B1(new_n655_), .B2(new_n618_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT78), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n657_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n307_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n659_), .A2(KEYINPUT78), .A3(new_n305_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n635_), .A2(new_n661_), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n651_), .A2(KEYINPUT37), .A3(new_n653_), .ZN(new_n663_));
  AOI21_X1  g462(.A(KEYINPUT37), .B1(new_n651_), .B2(new_n653_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(new_n327_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n666_), .A2(new_n277_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n662_), .A2(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT106), .ZN(new_n669_));
  INV_X1    g468(.A(new_n618_), .ZN(new_n670_));
  NOR3_X1   g469(.A1(new_n669_), .A2(G1gat), .A3(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n656_), .B1(new_n671_), .B2(KEYINPUT38), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT107), .ZN(new_n673_));
  INV_X1    g472(.A(new_n669_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n674_), .A2(new_n202_), .A3(new_n618_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT38), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n673_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n671_), .A2(KEYINPUT107), .A3(KEYINPUT38), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n672_), .B1(new_n677_), .B2(new_n678_), .ZN(G1324gat));
  INV_X1    g478(.A(KEYINPUT40), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT109), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT108), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n632_), .A2(new_n633_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n655_), .A2(new_n682_), .A3(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(G8gat), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n682_), .B1(new_n655_), .B2(new_n683_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n681_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n686_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n688_), .A2(KEYINPUT109), .A3(G8gat), .A4(new_n684_), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n687_), .A2(new_n689_), .A3(KEYINPUT39), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n683_), .A2(new_n287_), .ZN(new_n691_));
  OAI22_X1  g490(.A1(new_n687_), .A2(KEYINPUT39), .B1(new_n669_), .B2(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n680_), .B1(new_n690_), .B2(new_n692_), .ZN(new_n693_));
  OR2_X1    g492(.A1(new_n687_), .A2(KEYINPUT39), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n687_), .A2(new_n689_), .A3(KEYINPUT39), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n669_), .A2(new_n691_), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n694_), .A2(KEYINPUT40), .A3(new_n695_), .A4(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n693_), .A2(new_n697_), .ZN(G1325gat));
  NAND2_X1  g497(.A1(new_n598_), .A2(KEYINPUT105), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n630_), .A2(new_n631_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n624_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  AND3_X1   g500(.A1(new_n528_), .A2(new_n607_), .A3(new_n608_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n607_), .B1(new_n528_), .B2(new_n608_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n604_), .A2(new_n590_), .A3(new_n587_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n528_), .A2(new_n608_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n614_), .B1(new_n704_), .B2(new_n707_), .ZN(new_n708_));
  OAI22_X1  g507(.A1(new_n708_), .A2(new_n624_), .B1(new_n530_), .B2(new_n598_), .ZN(new_n709_));
  AOI22_X1  g508(.A1(new_n701_), .A2(new_n619_), .B1(new_n709_), .B2(new_n402_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n654_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(new_n329_), .ZN(new_n713_));
  OAI21_X1  g512(.A(G15gat), .B1(new_n713_), .B2(new_n402_), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT41), .Z(new_n715_));
  OR2_X1    g514(.A1(new_n402_), .A2(G15gat), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n715_), .B1(new_n669_), .B2(new_n716_), .ZN(G1326gat));
  OAI21_X1  g516(.A(G22gat), .B1(new_n713_), .B2(new_n625_), .ZN(new_n718_));
  XOR2_X1   g517(.A(new_n718_), .B(KEYINPUT110), .Z(new_n719_));
  OR2_X1    g518(.A1(new_n719_), .A2(KEYINPUT42), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(KEYINPUT42), .ZN(new_n721_));
  OR3_X1    g520(.A1(new_n669_), .A2(G22gat), .A3(new_n625_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n720_), .A2(new_n721_), .A3(new_n722_), .ZN(G1327gat));
  NOR3_X1   g522(.A1(new_n277_), .A2(new_n654_), .A3(new_n327_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n662_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(G29gat), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n726_), .A2(new_n727_), .A3(new_n618_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT112), .ZN(new_n729_));
  OAI21_X1  g528(.A(KEYINPUT43), .B1(new_n710_), .B2(new_n665_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT43), .ZN(new_n731_));
  INV_X1    g530(.A(new_n665_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n635_), .A2(new_n731_), .A3(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n730_), .A2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT44), .ZN(new_n735_));
  AOI211_X1 g534(.A(new_n327_), .B(new_n310_), .C1(KEYINPUT111), .C2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n735_), .A2(KEYINPUT111), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  OAI211_X1 g538(.A(new_n734_), .B(new_n736_), .C1(KEYINPUT111), .C2(new_n735_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(new_n618_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n729_), .B1(new_n742_), .B2(G29gat), .ZN(new_n743_));
  AOI211_X1 g542(.A(KEYINPUT112), .B(new_n727_), .C1(new_n741_), .C2(new_n618_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n728_), .B1(new_n743_), .B2(new_n744_), .ZN(G1328gat));
  INV_X1    g544(.A(new_n683_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n746_), .A2(G36gat), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n662_), .A2(new_n724_), .A3(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(KEYINPUT113), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT113), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n662_), .A2(new_n750_), .A3(new_n724_), .A4(new_n747_), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n749_), .A2(KEYINPUT45), .A3(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(KEYINPUT45), .B1(new_n749_), .B2(new_n751_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n746_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n755_));
  INV_X1    g554(.A(G36gat), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n754_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT46), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n754_), .B(KEYINPUT46), .C1(new_n755_), .C2(new_n756_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(G1329gat));
  AOI21_X1  g560(.A(new_n402_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n762_));
  INV_X1    g561(.A(G43gat), .ZN(new_n763_));
  INV_X1    g562(.A(new_n402_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(new_n763_), .ZN(new_n765_));
  OAI22_X1  g564(.A1(new_n762_), .A2(new_n763_), .B1(new_n725_), .B2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT47), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n766_), .B(new_n767_), .ZN(G1330gat));
  AOI21_X1  g567(.A(G50gat), .B1(new_n726_), .B2(new_n624_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n624_), .A2(G50gat), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n741_), .B2(new_n770_), .ZN(G1331gat));
  NOR2_X1   g570(.A1(new_n710_), .A2(new_n309_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n666_), .A2(new_n278_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(G57gat), .B1(new_n775_), .B2(new_n618_), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n658_), .A2(new_n660_), .A3(new_n327_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n778_), .A2(new_n278_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n712_), .A2(G57gat), .A3(new_n618_), .A4(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT114), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n780_), .A2(new_n781_), .ZN(new_n783_));
  NOR3_X1   g582(.A1(new_n776_), .A2(new_n782_), .A3(new_n783_), .ZN(G1332gat));
  NAND2_X1  g583(.A1(new_n712_), .A2(new_n779_), .ZN(new_n785_));
  OAI21_X1  g584(.A(G64gat), .B1(new_n785_), .B2(new_n746_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(KEYINPUT115), .B(KEYINPUT48), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n786_), .B(new_n787_), .ZN(new_n788_));
  OR2_X1    g587(.A1(new_n746_), .A2(G64gat), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n788_), .B1(new_n774_), .B2(new_n789_), .ZN(G1333gat));
  OAI21_X1  g589(.A(G71gat), .B1(new_n785_), .B2(new_n402_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n791_), .B(KEYINPUT49), .ZN(new_n792_));
  OR2_X1    g591(.A1(new_n402_), .A2(G71gat), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n792_), .B1(new_n774_), .B2(new_n793_), .ZN(G1334gat));
  OAI21_X1  g593(.A(G78gat), .B1(new_n785_), .B2(new_n625_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT50), .ZN(new_n796_));
  OR2_X1    g595(.A1(new_n625_), .A2(G78gat), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n796_), .B1(new_n774_), .B2(new_n797_), .ZN(G1335gat));
  NAND3_X1  g597(.A1(new_n277_), .A2(new_n308_), .A3(new_n328_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n799_), .B1(new_n730_), .B2(new_n733_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(G85gat), .B1(new_n801_), .B2(new_n670_), .ZN(new_n802_));
  NOR3_X1   g601(.A1(new_n278_), .A2(new_n654_), .A3(new_n327_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n772_), .A2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n805_), .A2(new_n227_), .A3(new_n618_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n802_), .A2(new_n806_), .ZN(G1336gat));
  OAI21_X1  g606(.A(G92gat), .B1(new_n801_), .B2(new_n746_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n805_), .A2(new_n228_), .A3(new_n683_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(G1337gat));
  NOR3_X1   g609(.A1(new_n804_), .A2(new_n402_), .A3(new_n224_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n800_), .A2(new_n764_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n811_), .B1(G99gat), .B2(new_n812_), .ZN(new_n813_));
  XOR2_X1   g612(.A(new_n813_), .B(KEYINPUT51), .Z(G1338gat));
  INV_X1    g613(.A(new_n799_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n731_), .B1(new_n635_), .B2(new_n732_), .ZN(new_n816_));
  AOI211_X1 g615(.A(KEYINPUT43), .B(new_n665_), .C1(new_n617_), .C2(new_n634_), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n624_), .B(new_n815_), .C1(new_n816_), .C2(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(G106gat), .B1(new_n818_), .B2(KEYINPUT116), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT116), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n820_), .B1(new_n800_), .B2(new_n624_), .ZN(new_n821_));
  OAI21_X1  g620(.A(KEYINPUT52), .B1(new_n819_), .B2(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n800_), .A2(new_n820_), .A3(new_n624_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n818_), .A2(KEYINPUT116), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n823_), .A2(new_n824_), .A3(new_n825_), .A4(G106gat), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n822_), .A2(new_n826_), .ZN(new_n827_));
  OR3_X1    g626(.A1(new_n804_), .A2(G106gat), .A3(new_n625_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT53), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n827_), .A2(new_n831_), .A3(new_n828_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(G1339gat));
  NAND3_X1  g632(.A1(new_n701_), .A2(new_n618_), .A3(new_n764_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n293_), .A2(new_n294_), .A3(new_n298_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n304_), .B1(new_n297_), .B2(new_n295_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n305_), .A2(new_n837_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n838_), .A2(new_n271_), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n261_), .B(new_n245_), .C1(new_n256_), .C2(new_n259_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n246_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT55), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n260_), .A2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n255_), .B1(new_n254_), .B2(KEYINPUT12), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n257_), .A2(KEYINPUT67), .A3(new_n258_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n846_), .A2(KEYINPUT55), .A3(new_n245_), .A4(new_n253_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n841_), .A2(new_n843_), .A3(new_n847_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n848_), .A2(KEYINPUT56), .A3(new_n269_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(KEYINPUT56), .B1(new_n848_), .B2(new_n269_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n839_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT58), .ZN(new_n853_));
  OR2_X1    g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n852_), .A2(new_n853_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n854_), .A2(new_n732_), .A3(new_n855_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n308_), .A2(new_n271_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n849_), .B1(new_n851_), .B2(KEYINPUT118), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n848_), .A2(new_n269_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT56), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n859_), .A2(KEYINPUT118), .A3(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n857_), .B1(new_n858_), .B2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT119), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT119), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n857_), .B(new_n864_), .C1(new_n858_), .C2(new_n861_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n273_), .A2(new_n838_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n863_), .A2(new_n865_), .A3(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n654_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT120), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n870_), .A2(KEYINPUT57), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n856_), .B1(new_n869_), .B2(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n866_), .B1(new_n862_), .B2(KEYINPUT119), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n711_), .B1(new_n873_), .B2(new_n865_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n871_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n328_), .B1(new_n872_), .B2(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(KEYINPUT117), .B1(new_n778_), .B2(new_n277_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT117), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n278_), .A2(new_n777_), .A3(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n732_), .B1(new_n878_), .B2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT54), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n881_), .B(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n834_), .B1(new_n877_), .B2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  XOR2_X1   g685(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n887_));
  OAI211_X1 g686(.A(new_n886_), .B(new_n661_), .C1(new_n884_), .C2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(G113gat), .ZN(new_n889_));
  INV_X1    g688(.A(G113gat), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n884_), .A2(new_n890_), .A3(new_n309_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n891_), .ZN(G1340gat));
  OAI211_X1 g691(.A(new_n886_), .B(new_n277_), .C1(new_n884_), .C2(new_n887_), .ZN(new_n893_));
  XOR2_X1   g692(.A(KEYINPUT122), .B(G120gat), .Z(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n893_), .A2(new_n895_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n894_), .B1(new_n278_), .B2(KEYINPUT60), .ZN(new_n897_));
  OAI211_X1 g696(.A(new_n884_), .B(new_n897_), .C1(KEYINPUT60), .C2(new_n894_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n896_), .A2(new_n898_), .ZN(G1341gat));
  OAI211_X1 g698(.A(new_n886_), .B(new_n327_), .C1(new_n884_), .C2(new_n887_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(G127gat), .ZN(new_n901_));
  INV_X1    g700(.A(G127gat), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n884_), .A2(new_n902_), .A3(new_n327_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n901_), .A2(new_n903_), .ZN(G1342gat));
  OAI211_X1 g703(.A(new_n886_), .B(new_n732_), .C1(new_n884_), .C2(new_n887_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(G134gat), .ZN(new_n906_));
  INV_X1    g705(.A(G134gat), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n884_), .A2(new_n907_), .A3(new_n711_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n906_), .A2(new_n908_), .ZN(G1343gat));
  NAND3_X1  g708(.A1(new_n624_), .A2(new_n618_), .A3(new_n402_), .ZN(new_n910_));
  AOI211_X1 g709(.A(new_n683_), .B(new_n910_), .C1(new_n877_), .C2(new_n883_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n309_), .ZN(new_n912_));
  XOR2_X1   g711(.A(KEYINPUT123), .B(G141gat), .Z(new_n913_));
  XNOR2_X1  g712(.A(new_n912_), .B(new_n913_), .ZN(G1344gat));
  NAND2_X1  g713(.A1(new_n911_), .A2(new_n277_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g715(.A1(new_n911_), .A2(new_n327_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(KEYINPUT61), .B(G155gat), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n917_), .B(new_n918_), .ZN(G1346gat));
  INV_X1    g718(.A(G162gat), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n911_), .A2(new_n920_), .A3(new_n711_), .ZN(new_n921_));
  AND2_X1   g720(.A1(new_n911_), .A2(new_n732_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n921_), .B1(new_n922_), .B2(new_n920_), .ZN(G1347gat));
  INV_X1    g722(.A(KEYINPUT62), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n746_), .B1(new_n877_), .B2(new_n883_), .ZN(new_n925_));
  NOR3_X1   g724(.A1(new_n624_), .A2(new_n402_), .A3(new_n618_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n925_), .A2(new_n309_), .A3(new_n926_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n924_), .B1(new_n927_), .B2(G169gat), .ZN(new_n928_));
  INV_X1    g727(.A(new_n856_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n929_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n869_), .A2(new_n871_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n327_), .B1(new_n930_), .B2(new_n931_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n881_), .A2(new_n882_), .ZN(new_n933_));
  AOI211_X1 g732(.A(KEYINPUT54), .B(new_n732_), .C1(new_n878_), .C2(new_n880_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n933_), .A2(new_n934_), .ZN(new_n935_));
  OAI211_X1 g734(.A(new_n683_), .B(new_n926_), .C1(new_n932_), .C2(new_n935_), .ZN(new_n936_));
  OAI211_X1 g735(.A(new_n924_), .B(G169gat), .C1(new_n936_), .C2(new_n308_), .ZN(new_n937_));
  INV_X1    g736(.A(new_n937_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n309_), .A2(new_n369_), .A3(new_n371_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n939_), .B(KEYINPUT124), .ZN(new_n940_));
  OAI22_X1  g739(.A1(new_n928_), .A2(new_n938_), .B1(new_n936_), .B2(new_n940_), .ZN(G1348gat));
  NOR2_X1   g740(.A1(new_n936_), .A2(new_n278_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n942_), .B(new_n372_), .ZN(G1349gat));
  NOR2_X1   g742(.A1(new_n936_), .A2(new_n328_), .ZN(new_n944_));
  OAI221_X1 g743(.A(new_n944_), .B1(KEYINPUT125), .B2(G183gat), .C1(new_n562_), .C2(new_n563_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n354_), .A2(KEYINPUT125), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n946_), .B1(new_n936_), .B2(new_n328_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n945_), .A2(new_n947_), .ZN(G1350gat));
  OAI21_X1  g747(.A(G190gat), .B1(new_n936_), .B2(new_n665_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n711_), .A2(new_n559_), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n949_), .B1(new_n936_), .B2(new_n950_), .ZN(G1351gat));
  NOR2_X1   g750(.A1(new_n764_), .A2(new_n530_), .ZN(new_n952_));
  XNOR2_X1  g751(.A(new_n952_), .B(KEYINPUT126), .ZN(new_n953_));
  OAI211_X1 g752(.A(new_n683_), .B(new_n953_), .C1(new_n932_), .C2(new_n935_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n954_), .A2(new_n308_), .ZN(new_n955_));
  XNOR2_X1  g754(.A(new_n955_), .B(new_n411_), .ZN(G1352gat));
  NOR2_X1   g755(.A1(new_n954_), .A2(new_n278_), .ZN(new_n957_));
  XNOR2_X1  g756(.A(new_n957_), .B(new_n413_), .ZN(G1353gat));
  OAI22_X1  g757(.A1(new_n954_), .A2(new_n328_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n959_));
  XNOR2_X1  g758(.A(KEYINPUT63), .B(G211gat), .ZN(new_n960_));
  NAND4_X1  g759(.A1(new_n925_), .A2(new_n327_), .A3(new_n953_), .A4(new_n960_), .ZN(new_n961_));
  INV_X1    g760(.A(KEYINPUT127), .ZN(new_n962_));
  AND3_X1   g761(.A1(new_n959_), .A2(new_n961_), .A3(new_n962_), .ZN(new_n963_));
  AOI21_X1  g762(.A(new_n962_), .B1(new_n959_), .B2(new_n961_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n963_), .A2(new_n964_), .ZN(G1354gat));
  OAI21_X1  g764(.A(G218gat), .B1(new_n954_), .B2(new_n665_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n711_), .A2(new_n406_), .ZN(new_n967_));
  OAI21_X1  g766(.A(new_n966_), .B1(new_n954_), .B2(new_n967_), .ZN(G1355gat));
endmodule


