//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 0 1 1 1 0 1 0 1 1 0 0 1 0 1 1 0 1 0 0 0 1 0 1 1 1 0 1 1 0 0 0 1 1 1 1 0 0 1 0 1 1 0 1 0 1 0 1 1 1 0 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n932_, new_n933_, new_n934_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n942_, new_n943_, new_n944_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n959_,
    new_n960_, new_n962_, new_n963_, new_n964_, new_n966_, new_n967_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n980_, new_n981_, new_n982_;
  XNOR2_X1  g000(.A(G71gat), .B(G99gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G43gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G227gat), .A2(G233gat), .ZN(new_n204_));
  INV_X1    g003(.A(G15gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n203_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT84), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  AND2_X1   g009(.A1(KEYINPUT81), .A2(KEYINPUT23), .ZN(new_n211_));
  NOR2_X1   g010(.A1(KEYINPUT81), .A2(KEYINPUT23), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n210_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G183gat), .ZN(new_n214_));
  INV_X1    g013(.A(G190gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT23), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n209_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n213_), .A2(new_n216_), .A3(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220_));
  INV_X1    g019(.A(G176gat), .ZN(new_n221_));
  INV_X1    g020(.A(G169gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT22), .B1(new_n222_), .B2(KEYINPUT82), .ZN(new_n223_));
  OR2_X1    g022(.A1(new_n222_), .A2(KEYINPUT22), .ZN(new_n224_));
  OAI211_X1 g023(.A(new_n221_), .B(new_n223_), .C1(new_n224_), .C2(KEYINPUT82), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n219_), .A2(new_n220_), .A3(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT24), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n227_), .B1(G169gat), .B2(G176gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT79), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n229_), .A2(new_n222_), .A3(new_n221_), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT79), .B1(G169gat), .B2(G176gat), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n228_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT80), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT80), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n228_), .A2(new_n230_), .A3(new_n234_), .A4(new_n231_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n230_), .A2(new_n231_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(new_n227_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n209_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n210_), .A2(new_n217_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT25), .B(G183gat), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT26), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n243_), .A2(KEYINPUT78), .A3(G190gat), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT78), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT26), .B1(new_n245_), .B2(new_n215_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n242_), .A2(new_n244_), .A3(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n238_), .A2(new_n241_), .A3(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n226_), .B1(new_n236_), .B2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT83), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT83), .ZN(new_n251_));
  OAI211_X1 g050(.A(new_n226_), .B(new_n251_), .C1(new_n236_), .C2(new_n248_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT30), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n250_), .A2(KEYINPUT30), .A3(new_n252_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n208_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n255_), .A2(new_n208_), .A3(new_n256_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n207_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n207_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n257_), .A2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G127gat), .B(G134gat), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  XOR2_X1   g063(.A(G113gat), .B(G120gat), .Z(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G113gat), .B(G120gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n263_), .A2(new_n267_), .ZN(new_n268_));
  AND2_X1   g067(.A1(new_n266_), .A2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(KEYINPUT31), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  OR3_X1    g070(.A1(new_n260_), .A2(new_n262_), .A3(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n271_), .B1(new_n260_), .B2(new_n262_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT91), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT89), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G228gat), .A2(G233gat), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G197gat), .B(G204gat), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT21), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G211gat), .B(G218gat), .ZN(new_n282_));
  INV_X1    g081(.A(G197gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(G204gat), .ZN(new_n284_));
  INV_X1    g083(.A(G204gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(G197gat), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT88), .ZN(new_n287_));
  AND3_X1   g086(.A1(new_n284_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n288_));
  OAI21_X1  g087(.A(KEYINPUT21), .B1(new_n284_), .B2(new_n287_), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n281_), .B(new_n282_), .C1(new_n288_), .C2(new_n289_), .ZN(new_n290_));
  OR3_X1    g089(.A1(new_n279_), .A2(new_n282_), .A3(new_n280_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n278_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT29), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G155gat), .A2(G162gat), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(G155gat), .A2(G162gat), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(G141gat), .ZN(new_n299_));
  INV_X1    g098(.A(G148gat), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n299_), .A2(new_n300_), .A3(KEYINPUT85), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT85), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n302_), .B1(G141gat), .B2(G148gat), .ZN(new_n303_));
  OR2_X1    g102(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n304_));
  NAND2_X1  g103(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n305_));
  AND4_X1   g104(.A1(new_n301_), .A2(new_n303_), .A3(new_n304_), .A4(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G141gat), .A2(G148gat), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT87), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT2), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n307_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  OAI21_X1  g109(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n311_));
  AOI21_X1  g110(.A(KEYINPUT87), .B1(G141gat), .B2(G148gat), .ZN(new_n312_));
  OAI211_X1 g111(.A(new_n310_), .B(new_n311_), .C1(new_n309_), .C2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n298_), .B1(new_n306_), .B2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n299_), .A2(new_n300_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(new_n307_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n297_), .B1(KEYINPUT1), .B2(new_n295_), .ZN(new_n317_));
  OR2_X1    g116(.A1(new_n295_), .A2(KEYINPUT1), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n316_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n294_), .B1(new_n314_), .B2(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n276_), .B1(new_n293_), .B2(new_n321_), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n301_), .A2(new_n303_), .A3(new_n304_), .A4(new_n305_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n312_), .A2(new_n309_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND4_X1  g124(.A1(new_n323_), .A2(new_n325_), .A3(new_n311_), .A4(new_n310_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n319_), .B1(new_n326_), .B2(new_n298_), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n292_), .B(KEYINPUT89), .C1(new_n327_), .C2(new_n294_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT90), .ZN(new_n329_));
  AND3_X1   g128(.A1(new_n290_), .A2(new_n291_), .A3(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n329_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n331_));
  OAI22_X1  g130(.A1(new_n330_), .A2(new_n331_), .B1(new_n327_), .B2(new_n294_), .ZN(new_n332_));
  AOI22_X1  g131(.A1(new_n322_), .A2(new_n328_), .B1(new_n332_), .B2(new_n278_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G78gat), .B(G106gat), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n275_), .B1(new_n333_), .B2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n327_), .A2(new_n294_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G22gat), .B(G50gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT28), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n337_), .B(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n322_), .A2(new_n328_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n332_), .A2(new_n278_), .ZN(new_n343_));
  AND3_X1   g142(.A1(new_n342_), .A2(new_n343_), .A3(new_n335_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n335_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n345_));
  OAI22_X1  g144(.A1(new_n336_), .A2(new_n341_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n342_), .A2(new_n343_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(new_n334_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n333_), .A2(new_n335_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n348_), .A2(new_n349_), .A3(new_n275_), .A4(new_n340_), .ZN(new_n350_));
  AND2_X1   g149(.A1(new_n346_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n298_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n310_), .A2(new_n311_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n353_), .A2(new_n324_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n352_), .B1(new_n354_), .B2(new_n323_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n269_), .B1(new_n355_), .B2(new_n319_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n266_), .A2(new_n268_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n314_), .A2(new_n320_), .A3(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n356_), .A2(KEYINPUT4), .A3(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G225gat), .A2(G233gat), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n357_), .B1(new_n314_), .B2(new_n320_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT95), .B(KEYINPUT4), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n360_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n359_), .A2(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n356_), .A2(new_n358_), .A3(new_n360_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G1gat), .B(G29gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G57gat), .B(G85gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n366_), .A2(new_n371_), .ZN(new_n372_));
  AND2_X1   g171(.A1(new_n359_), .A2(new_n363_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT99), .ZN(new_n374_));
  XOR2_X1   g173(.A(new_n369_), .B(new_n370_), .Z(new_n375_));
  NAND2_X1  g174(.A1(new_n365_), .A2(new_n375_), .ZN(new_n376_));
  NOR3_X1   g175(.A1(new_n373_), .A2(new_n374_), .A3(new_n376_), .ZN(new_n377_));
  AND3_X1   g176(.A1(new_n314_), .A2(new_n320_), .A3(new_n357_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n378_), .A2(new_n361_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n371_), .B1(new_n379_), .B2(new_n360_), .ZN(new_n380_));
  AOI21_X1  g179(.A(KEYINPUT99), .B1(new_n380_), .B2(new_n364_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n372_), .B1(new_n377_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G226gat), .A2(G233gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(KEYINPUT19), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n290_), .A2(new_n291_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n250_), .A2(new_n387_), .A3(new_n252_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT20), .ZN(new_n389_));
  INV_X1    g188(.A(new_n242_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT26), .B(G190gat), .ZN(new_n391_));
  OR2_X1    g190(.A1(new_n391_), .A2(KEYINPUT92), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(KEYINPUT92), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n390_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n238_), .A2(new_n213_), .A3(new_n218_), .A4(new_n232_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n241_), .A2(new_n216_), .ZN(new_n396_));
  XOR2_X1   g195(.A(KEYINPUT22), .B(G169gat), .Z(new_n397_));
  OAI21_X1  g196(.A(new_n220_), .B1(new_n397_), .B2(G176gat), .ZN(new_n398_));
  OAI22_X1  g197(.A1(new_n394_), .A2(new_n395_), .B1(new_n396_), .B2(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n389_), .B1(new_n399_), .B2(new_n386_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n385_), .B1(new_n388_), .B2(new_n400_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n384_), .A2(new_n389_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n402_), .B1(new_n399_), .B2(new_n386_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n403_), .B1(new_n253_), .B2(new_n386_), .ZN(new_n404_));
  XOR2_X1   g203(.A(G8gat), .B(G36gat), .Z(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G64gat), .B(G92gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n409_), .A2(KEYINPUT32), .ZN(new_n410_));
  OR3_X1    g209(.A1(new_n401_), .A2(new_n404_), .A3(new_n410_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n330_), .A2(new_n331_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n399_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n389_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n252_), .ZN(new_n415_));
  AOI22_X1  g214(.A1(new_n227_), .A2(new_n237_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n416_), .A2(new_n247_), .A3(new_n233_), .A4(new_n235_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n251_), .B1(new_n417_), .B2(new_n226_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n386_), .B1(new_n415_), .B2(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n385_), .B1(new_n414_), .B2(new_n419_), .ZN(new_n420_));
  AND3_X1   g219(.A1(new_n388_), .A2(new_n385_), .A3(new_n400_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n410_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n382_), .A2(new_n411_), .A3(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT100), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT100), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n382_), .A2(new_n411_), .A3(new_n425_), .A4(new_n422_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n380_), .A2(KEYINPUT33), .A3(new_n364_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(KEYINPUT97), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT97), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n380_), .A2(new_n430_), .A3(KEYINPUT33), .A4(new_n364_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n429_), .A2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT98), .B1(new_n373_), .B2(new_n376_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT33), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT98), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n380_), .A2(new_n435_), .A3(new_n364_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n433_), .A2(new_n434_), .A3(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n361_), .A2(new_n362_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n359_), .A2(new_n360_), .A3(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n379_), .A2(G225gat), .A3(G233gat), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n439_), .A2(new_n440_), .A3(new_n371_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n432_), .A2(new_n437_), .A3(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT94), .ZN(new_n443_));
  INV_X1    g242(.A(new_n409_), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n443_), .B(new_n444_), .C1(new_n401_), .C2(new_n404_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n388_), .A2(new_n400_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(new_n384_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n413_), .A2(new_n387_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n419_), .A2(new_n448_), .A3(new_n402_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n447_), .A2(new_n409_), .A3(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n444_), .B1(new_n401_), .B2(new_n404_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n450_), .A2(new_n451_), .A3(KEYINPUT94), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n442_), .B1(new_n445_), .B2(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n351_), .B1(new_n427_), .B2(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n382_), .B1(new_n346_), .B2(new_n350_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT27), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n452_), .A2(new_n456_), .A3(new_n445_), .ZN(new_n457_));
  XOR2_X1   g256(.A(new_n409_), .B(KEYINPUT101), .Z(new_n458_));
  OAI21_X1  g257(.A(new_n458_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n459_), .A2(KEYINPUT27), .A3(new_n450_), .ZN(new_n460_));
  AND3_X1   g259(.A1(new_n455_), .A2(new_n457_), .A3(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n274_), .B1(new_n454_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n457_), .A2(new_n460_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n382_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n274_), .A2(new_n465_), .A3(new_n466_), .A4(new_n351_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n463_), .A2(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G1gat), .B(G8gat), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT75), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n470_), .B(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G15gat), .B(G22gat), .ZN(new_n473_));
  INV_X1    g272(.A(G1gat), .ZN(new_n474_));
  INV_X1    g273(.A(G8gat), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT14), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n473_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n472_), .B(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G29gat), .B(G36gat), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  XOR2_X1   g280(.A(G43gat), .B(G50gat), .Z(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G43gat), .B(G50gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n480_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n479_), .A2(new_n487_), .ZN(new_n488_));
  OR2_X1    g287(.A1(new_n472_), .A2(new_n478_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n472_), .A2(new_n478_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n489_), .A2(new_n490_), .A3(new_n486_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n488_), .A2(KEYINPUT77), .A3(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G229gat), .A2(G233gat), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT77), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n479_), .A2(new_n495_), .A3(new_n487_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n492_), .A2(new_n494_), .A3(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT15), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n486_), .A2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n483_), .A2(KEYINPUT15), .A3(new_n485_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(new_n479_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n503_), .A2(new_n493_), .A3(new_n491_), .ZN(new_n504_));
  AND2_X1   g303(.A1(new_n497_), .A2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G113gat), .B(G141gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G169gat), .B(G197gat), .ZN(new_n507_));
  XOR2_X1   g306(.A(new_n506_), .B(new_n507_), .Z(new_n508_));
  XNOR2_X1  g307(.A(new_n505_), .B(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n469_), .A2(new_n510_), .ZN(new_n511_));
  XOR2_X1   g310(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n512_));
  NAND2_X1  g311(.A1(G232gat), .A2(G233gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n514_), .A2(KEYINPUT35), .ZN(new_n515_));
  XNOR2_X1  g314(.A(KEYINPUT10), .B(G99gat), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(KEYINPUT64), .B(G106gat), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  XOR2_X1   g318(.A(KEYINPUT65), .B(G92gat), .Z(new_n520_));
  INV_X1    g319(.A(G85gat), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n521_), .A2(KEYINPUT9), .ZN(new_n522_));
  AOI22_X1  g321(.A1(new_n517_), .A2(new_n519_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G85gat), .B(G92gat), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G99gat), .A2(G106gat), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT6), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT6), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n528_), .A2(G99gat), .A3(G106gat), .ZN(new_n529_));
  AOI22_X1  g328(.A1(new_n525_), .A2(KEYINPUT9), .B1(new_n527_), .B2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n523_), .A2(new_n530_), .A3(KEYINPUT66), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT66), .ZN(new_n532_));
  XNOR2_X1  g331(.A(KEYINPUT65), .B(G92gat), .ZN(new_n533_));
  INV_X1    g332(.A(new_n522_), .ZN(new_n534_));
  OAI22_X1  g333(.A1(new_n516_), .A2(new_n518_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT9), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n528_), .B1(G99gat), .B2(G106gat), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n526_), .A2(KEYINPUT6), .ZN(new_n538_));
  OAI22_X1  g337(.A1(new_n524_), .A2(new_n536_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n532_), .B1(new_n535_), .B2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n531_), .A2(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(G99gat), .A2(G106gat), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT7), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n537_), .A2(new_n538_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n525_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT8), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT8), .ZN(new_n548_));
  OAI211_X1 g347(.A(new_n548_), .B(new_n525_), .C1(new_n544_), .C2(new_n545_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n501_), .B1(new_n541_), .B2(new_n550_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n515_), .B1(new_n551_), .B2(KEYINPUT71), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n541_), .A2(new_n550_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(new_n502_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n541_), .A2(new_n550_), .A3(new_n486_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n514_), .A2(KEYINPUT35), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n552_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n554_), .A2(KEYINPUT71), .A3(new_n515_), .A4(new_n555_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G190gat), .B(G218gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G134gat), .B(G162gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n563_), .A2(KEYINPUT36), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n560_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(KEYINPUT72), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT72), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n560_), .A2(new_n567_), .A3(new_n564_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n566_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n564_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n563_), .A2(KEYINPUT36), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n558_), .A2(new_n570_), .A3(new_n559_), .A4(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n569_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(KEYINPUT74), .B(KEYINPUT37), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n566_), .A2(KEYINPUT73), .A3(new_n568_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT73), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n567_), .B1(new_n560_), .B2(new_n564_), .ZN(new_n578_));
  AOI211_X1 g377(.A(KEYINPUT72), .B(new_n570_), .C1(new_n558_), .C2(new_n559_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n577_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n576_), .A2(new_n580_), .A3(new_n572_), .ZN(new_n581_));
  AOI22_X1  g380(.A1(new_n574_), .A2(new_n575_), .B1(new_n581_), .B2(KEYINPUT37), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G57gat), .B(G64gat), .ZN(new_n583_));
  OR2_X1    g382(.A1(new_n583_), .A2(KEYINPUT11), .ZN(new_n584_));
  XOR2_X1   g383(.A(G71gat), .B(G78gat), .Z(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT67), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n583_), .A2(new_n587_), .A3(KEYINPUT11), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n587_), .B1(new_n583_), .B2(KEYINPUT11), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n586_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n590_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n592_), .A2(new_n584_), .A3(new_n585_), .A4(new_n588_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G231gat), .A2(G233gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n472_), .B(new_n477_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  XOR2_X1   g397(.A(G127gat), .B(G155gat), .Z(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT16), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G183gat), .B(G211gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT17), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n602_), .A2(new_n603_), .ZN(new_n605_));
  OR3_X1    g404(.A1(new_n598_), .A2(new_n604_), .A3(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n598_), .A2(new_n604_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT76), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n606_), .A2(KEYINPUT76), .A3(new_n607_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(G230gat), .A2(G233gat), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n591_), .A2(new_n593_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n553_), .A2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n594_), .A2(new_n550_), .A3(new_n541_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n617_), .A2(KEYINPUT12), .A3(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT12), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n553_), .A2(new_n620_), .A3(new_n616_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n615_), .B1(new_n619_), .B2(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n614_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G120gat), .B(G148gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT5), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G176gat), .B(G204gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n624_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT69), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n628_), .B(KEYINPUT68), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  OAI211_X1 g431(.A(new_n630_), .B(new_n632_), .C1(new_n622_), .C2(new_n623_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n629_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(KEYINPUT69), .B1(new_n624_), .B2(new_n631_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n635_), .A2(KEYINPUT13), .A3(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT13), .ZN(new_n638_));
  INV_X1    g437(.A(new_n636_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n638_), .B1(new_n639_), .B2(new_n634_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n637_), .A2(new_n640_), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n582_), .A2(new_n613_), .A3(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n511_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n644_), .A2(new_n474_), .A3(new_n382_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT38), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n452_), .A2(new_n445_), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n424_), .B(new_n426_), .C1(new_n647_), .C2(new_n442_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n461_), .B1(new_n648_), .B2(new_n351_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n467_), .B1(new_n649_), .B2(new_n274_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n650_), .A2(KEYINPUT103), .A3(new_n573_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(KEYINPUT103), .B1(new_n650_), .B2(new_n573_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n608_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n637_), .A2(new_n640_), .A3(new_n509_), .A4(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT102), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n657_), .A2(new_n658_), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n655_), .A2(new_n382_), .A3(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n646_), .B1(new_n474_), .B2(new_n663_), .ZN(G1324gat));
  INV_X1    g463(.A(KEYINPUT40), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n464_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT103), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n667_), .B1(new_n469_), .B2(new_n574_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n666_), .B1(new_n668_), .B2(new_n651_), .ZN(new_n669_));
  OAI21_X1  g468(.A(KEYINPUT104), .B1(new_n669_), .B2(new_n475_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT104), .ZN(new_n671_));
  OAI211_X1 g470(.A(new_n671_), .B(G8gat), .C1(new_n654_), .C2(new_n666_), .ZN(new_n672_));
  AND3_X1   g471(.A1(new_n670_), .A2(new_n672_), .A3(KEYINPUT39), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT39), .ZN(new_n674_));
  OAI211_X1 g473(.A(KEYINPUT104), .B(new_n674_), .C1(new_n669_), .C2(new_n475_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n644_), .A2(new_n475_), .A3(new_n464_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n665_), .B1(new_n673_), .B2(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n670_), .A2(new_n672_), .A3(KEYINPUT39), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n679_), .A2(KEYINPUT40), .A3(new_n675_), .A4(new_n676_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(G1325gat));
  NAND3_X1  g480(.A1(new_n644_), .A2(new_n205_), .A3(new_n274_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n655_), .A2(new_n662_), .A3(new_n274_), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n683_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n684_));
  AOI21_X1  g483(.A(KEYINPUT41), .B1(new_n683_), .B2(G15gat), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n682_), .B1(new_n684_), .B2(new_n685_), .ZN(G1326gat));
  OR3_X1    g485(.A1(new_n643_), .A2(G22gat), .A3(new_n351_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n351_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n655_), .A2(new_n662_), .A3(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT42), .ZN(new_n690_));
  AND3_X1   g489(.A1(new_n689_), .A2(new_n690_), .A3(G22gat), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n690_), .B1(new_n689_), .B2(G22gat), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n687_), .B1(new_n691_), .B2(new_n692_), .ZN(G1327gat));
  NOR3_X1   g492(.A1(new_n612_), .A2(new_n641_), .A3(new_n510_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n695_));
  OAI211_X1 g494(.A(new_n695_), .B(new_n582_), .C1(new_n463_), .C2(new_n468_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n695_), .B1(new_n650_), .B2(new_n582_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n694_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  OAI211_X1 g500(.A(KEYINPUT44), .B(new_n694_), .C1(new_n697_), .C2(new_n698_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(G29gat), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n466_), .A2(new_n704_), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n612_), .A2(new_n641_), .A3(new_n573_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n511_), .A2(KEYINPUT105), .A3(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n706_), .A2(new_n650_), .A3(new_n509_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT105), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n707_), .A2(new_n382_), .A3(new_n710_), .ZN(new_n711_));
  AOI22_X1  g510(.A1(new_n703_), .A2(new_n705_), .B1(new_n704_), .B2(new_n711_), .ZN(G1328gat));
  NAND3_X1  g511(.A1(new_n701_), .A2(new_n464_), .A3(new_n702_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(G36gat), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n465_), .A2(G36gat), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n707_), .A2(new_n710_), .A3(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(KEYINPUT45), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT45), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n707_), .A2(new_n718_), .A3(new_n710_), .A4(new_n715_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n714_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT46), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n714_), .A2(KEYINPUT46), .A3(new_n720_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1329gat));
  NAND4_X1  g524(.A1(new_n701_), .A2(G43gat), .A3(new_n274_), .A4(new_n702_), .ZN(new_n726_));
  INV_X1    g525(.A(G43gat), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n707_), .A2(new_n710_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n274_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n727_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n726_), .A2(new_n730_), .ZN(new_n731_));
  XOR2_X1   g530(.A(KEYINPUT106), .B(KEYINPUT47), .Z(new_n732_));
  XNOR2_X1  g531(.A(new_n731_), .B(new_n732_), .ZN(G1330gat));
  OR3_X1    g532(.A1(new_n728_), .A2(G50gat), .A3(new_n351_), .ZN(new_n734_));
  AOI21_X1  g533(.A(KEYINPUT107), .B1(new_n703_), .B2(new_n688_), .ZN(new_n735_));
  NAND4_X1  g534(.A1(new_n701_), .A2(KEYINPUT107), .A3(new_n688_), .A4(new_n702_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(G50gat), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n734_), .B1(new_n735_), .B2(new_n737_), .ZN(G1331gat));
  NAND2_X1  g537(.A1(new_n641_), .A2(new_n510_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n739_), .A2(new_n613_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n655_), .A2(new_n382_), .A3(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(G57gat), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n469_), .A2(new_n739_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n582_), .A2(new_n613_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  OR2_X1    g544(.A1(new_n466_), .A2(G57gat), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n742_), .B1(new_n745_), .B2(new_n746_), .ZN(G1332gat));
  OR3_X1    g546(.A1(new_n745_), .A2(G64gat), .A3(new_n465_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n655_), .A2(new_n464_), .A3(new_n740_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT48), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n749_), .A2(new_n750_), .A3(G64gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(new_n749_), .B2(G64gat), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n748_), .B1(new_n751_), .B2(new_n752_), .ZN(G1333gat));
  OR3_X1    g552(.A1(new_n745_), .A2(G71gat), .A3(new_n729_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n655_), .A2(new_n274_), .A3(new_n740_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT49), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n755_), .A2(new_n756_), .A3(G71gat), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n755_), .B2(G71gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n754_), .B1(new_n757_), .B2(new_n758_), .ZN(G1334gat));
  OR3_X1    g558(.A1(new_n745_), .A2(G78gat), .A3(new_n351_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n655_), .A2(new_n688_), .A3(new_n740_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT50), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n761_), .A2(new_n762_), .A3(G78gat), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n762_), .B1(new_n761_), .B2(G78gat), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n760_), .B1(new_n763_), .B2(new_n764_), .ZN(G1335gat));
  NAND3_X1  g564(.A1(new_n743_), .A2(new_n574_), .A3(new_n613_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n521_), .B1(new_n766_), .B2(new_n466_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT108), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n768_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n697_), .A2(new_n698_), .ZN(new_n771_));
  NOR3_X1   g570(.A1(new_n771_), .A2(new_n612_), .A3(new_n739_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n466_), .A2(new_n521_), .ZN(new_n773_));
  AOI22_X1  g572(.A1(new_n769_), .A2(new_n770_), .B1(new_n772_), .B2(new_n773_), .ZN(G1336gat));
  NAND3_X1  g573(.A1(new_n772_), .A2(new_n520_), .A3(new_n464_), .ZN(new_n775_));
  INV_X1    g574(.A(G92gat), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n776_), .B1(new_n766_), .B2(new_n465_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT109), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n778_), .B(new_n779_), .ZN(G1337gat));
  INV_X1    g579(.A(G99gat), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n781_), .B1(new_n772_), .B2(new_n274_), .ZN(new_n782_));
  NOR3_X1   g581(.A1(new_n766_), .A2(new_n516_), .A3(new_n729_), .ZN(new_n783_));
  OR3_X1    g582(.A1(new_n782_), .A2(KEYINPUT51), .A3(new_n783_), .ZN(new_n784_));
  OAI21_X1  g583(.A(KEYINPUT51), .B1(new_n782_), .B2(new_n783_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(G1338gat));
  OR3_X1    g585(.A1(new_n766_), .A2(new_n518_), .A3(new_n351_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n739_), .A2(new_n612_), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n688_), .B(new_n788_), .C1(new_n697_), .C2(new_n698_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT52), .ZN(new_n790_));
  AND4_X1   g589(.A1(KEYINPUT110), .A2(new_n789_), .A3(new_n790_), .A4(G106gat), .ZN(new_n791_));
  INV_X1    g590(.A(G106gat), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT110), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n792_), .B1(new_n793_), .B2(KEYINPUT52), .ZN(new_n794_));
  AOI22_X1  g593(.A1(new_n789_), .A2(new_n794_), .B1(KEYINPUT110), .B2(new_n790_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n787_), .B1(new_n791_), .B2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(KEYINPUT53), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n798_));
  OAI211_X1 g597(.A(new_n798_), .B(new_n787_), .C1(new_n791_), .C2(new_n795_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n797_), .A2(new_n799_), .ZN(G1339gat));
  XNOR2_X1  g599(.A(KEYINPUT114), .B(KEYINPUT57), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n497_), .A2(new_n504_), .A3(new_n508_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n492_), .A2(new_n493_), .A3(new_n496_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT113), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n493_), .B1(new_n597_), .B2(new_n486_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n508_), .B1(new_n806_), .B2(new_n503_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n804_), .A2(new_n805_), .A3(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n803_), .A2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n805_), .B1(new_n804_), .B2(new_n807_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n811_), .B1(new_n639_), .B2(new_n634_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  AND3_X1   g612(.A1(new_n617_), .A2(KEYINPUT12), .A3(new_n618_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n621_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n614_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n619_), .A2(new_n615_), .A3(new_n621_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n816_), .A2(new_n817_), .A3(KEYINPUT55), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n631_), .B1(new_n622_), .B2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n820_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(KEYINPUT111), .B(KEYINPUT56), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT112), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n818_), .A2(new_n820_), .A3(KEYINPUT56), .ZN(new_n826_));
  AND3_X1   g625(.A1(new_n619_), .A2(new_n615_), .A3(new_n621_), .ZN(new_n827_));
  NOR3_X1   g626(.A1(new_n827_), .A2(new_n622_), .A3(new_n819_), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n819_), .B(new_n614_), .C1(new_n814_), .C2(new_n815_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n632_), .ZN(new_n830_));
  OAI211_X1 g629(.A(KEYINPUT112), .B(new_n822_), .C1(new_n828_), .C2(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n825_), .A2(new_n826_), .A3(new_n831_), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n509_), .A2(new_n629_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n813_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n802_), .B1(new_n834_), .B2(new_n574_), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n811_), .A2(new_n629_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n826_), .ZN(new_n837_));
  AOI21_X1  g636(.A(KEYINPUT56), .B1(new_n818_), .B2(new_n820_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n836_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT58), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n581_), .A2(KEYINPUT37), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n569_), .A2(new_n572_), .A3(new_n575_), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n836_), .B(KEYINPUT58), .C1(new_n837_), .C2(new_n838_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n841_), .A2(new_n842_), .A3(new_n843_), .A4(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n831_), .A2(new_n826_), .ZN(new_n846_));
  AOI21_X1  g645(.A(KEYINPUT112), .B1(new_n821_), .B2(new_n822_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n833_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n812_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n573_), .A2(KEYINPUT57), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(KEYINPUT115), .B1(new_n849_), .B2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT115), .ZN(new_n853_));
  AOI211_X1 g652(.A(new_n853_), .B(new_n850_), .C1(new_n848_), .C2(new_n812_), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n835_), .B(new_n845_), .C1(new_n852_), .C2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n842_), .A2(new_n843_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n641_), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n856_), .A2(new_n857_), .A3(new_n510_), .A4(new_n612_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(KEYINPUT54), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT54), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n744_), .A2(new_n860_), .A3(new_n510_), .A4(new_n857_), .ZN(new_n861_));
  AOI22_X1  g660(.A1(new_n855_), .A2(new_n608_), .B1(new_n859_), .B2(new_n861_), .ZN(new_n862_));
  NOR4_X1   g661(.A1(new_n729_), .A2(new_n466_), .A3(new_n688_), .A4(new_n464_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT116), .ZN(new_n864_));
  OR2_X1    g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n863_), .A2(new_n864_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n862_), .A2(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(G113gat), .B1(new_n868_), .B2(new_n509_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n855_), .A2(new_n613_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n861_), .A2(new_n859_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  AND2_X1   g671(.A1(new_n865_), .A2(new_n866_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT117), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(KEYINPUT59), .B1(new_n867_), .B2(KEYINPUT117), .ZN(new_n876_));
  AND2_X1   g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n852_), .A2(new_n854_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n574_), .B1(new_n848_), .B2(new_n812_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n845_), .B1(new_n879_), .B2(new_n801_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n608_), .B1(new_n878_), .B2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n871_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(new_n873_), .ZN(new_n883_));
  AOI22_X1  g682(.A1(new_n872_), .A2(new_n877_), .B1(new_n883_), .B2(KEYINPUT59), .ZN(new_n884_));
  INV_X1    g683(.A(G113gat), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n885_), .B1(new_n509_), .B2(KEYINPUT118), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n886_), .B1(KEYINPUT118), .B2(new_n885_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n869_), .B1(new_n884_), .B2(new_n887_), .ZN(G1340gat));
  NAND3_X1  g687(.A1(new_n872_), .A2(new_n875_), .A3(new_n876_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT59), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n889_), .B(new_n641_), .C1(new_n890_), .C2(new_n868_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(G120gat), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n857_), .A2(KEYINPUT60), .ZN(new_n893_));
  MUX2_X1   g692(.A(new_n893_), .B(KEYINPUT60), .S(G120gat), .Z(new_n894_));
  NAND2_X1  g693(.A1(new_n868_), .A2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT119), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n868_), .A2(KEYINPUT119), .A3(new_n894_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n892_), .A2(new_n899_), .ZN(G1341gat));
  OAI211_X1 g699(.A(new_n889_), .B(new_n656_), .C1(new_n890_), .C2(new_n868_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(G127gat), .ZN(new_n902_));
  OR3_X1    g701(.A1(new_n883_), .A2(G127gat), .A3(new_n613_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(G1342gat));
  NAND3_X1  g703(.A1(new_n882_), .A2(new_n574_), .A3(new_n873_), .ZN(new_n905_));
  INV_X1    g704(.A(G134gat), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(KEYINPUT120), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT120), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n905_), .A2(new_n909_), .A3(new_n906_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n856_), .A2(new_n906_), .ZN(new_n911_));
  AOI22_X1  g710(.A1(new_n908_), .A2(new_n910_), .B1(new_n884_), .B2(new_n911_), .ZN(G1343gat));
  INV_X1    g711(.A(KEYINPUT122), .ZN(new_n913_));
  NOR4_X1   g712(.A1(new_n274_), .A2(new_n464_), .A3(new_n466_), .A4(new_n351_), .ZN(new_n914_));
  XOR2_X1   g713(.A(new_n914_), .B(KEYINPUT121), .Z(new_n915_));
  AOI21_X1  g714(.A(new_n913_), .B1(new_n882_), .B2(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n915_), .ZN(new_n917_));
  AOI211_X1 g716(.A(KEYINPUT122), .B(new_n917_), .C1(new_n881_), .C2(new_n871_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n509_), .B1(new_n916_), .B2(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(G141gat), .ZN(new_n920_));
  OAI21_X1  g719(.A(KEYINPUT122), .B1(new_n862_), .B2(new_n917_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n880_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n853_), .B1(new_n834_), .B2(new_n850_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n849_), .A2(new_n851_), .A3(KEYINPUT115), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(new_n924_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n656_), .B1(new_n922_), .B2(new_n925_), .ZN(new_n926_));
  AND2_X1   g725(.A1(new_n861_), .A2(new_n859_), .ZN(new_n927_));
  OAI211_X1 g726(.A(new_n913_), .B(new_n915_), .C1(new_n926_), .C2(new_n927_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n921_), .A2(new_n928_), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n929_), .A2(new_n299_), .A3(new_n509_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n920_), .A2(new_n930_), .ZN(G1344gat));
  OAI21_X1  g730(.A(new_n641_), .B1(new_n916_), .B2(new_n918_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(G148gat), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n929_), .A2(new_n300_), .A3(new_n641_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n933_), .A2(new_n934_), .ZN(G1345gat));
  XNOR2_X1  g734(.A(KEYINPUT61), .B(G155gat), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n936_), .B(KEYINPUT123), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n937_), .B1(new_n929_), .B2(new_n612_), .ZN(new_n938_));
  INV_X1    g737(.A(new_n937_), .ZN(new_n939_));
  AOI211_X1 g738(.A(new_n613_), .B(new_n939_), .C1(new_n921_), .C2(new_n928_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n938_), .A2(new_n940_), .ZN(G1346gat));
  INV_X1    g740(.A(G162gat), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n929_), .A2(new_n942_), .A3(new_n574_), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n856_), .B1(new_n921_), .B2(new_n928_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n943_), .B1(new_n942_), .B2(new_n944_), .ZN(G1347gat));
  NOR4_X1   g744(.A1(new_n729_), .A2(new_n465_), .A3(new_n382_), .A4(new_n688_), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n872_), .A2(new_n509_), .A3(new_n946_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n947_), .A2(G169gat), .ZN(new_n948_));
  INV_X1    g747(.A(KEYINPUT62), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n948_), .A2(new_n949_), .ZN(new_n950_));
  NAND3_X1  g749(.A1(new_n947_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n951_));
  OAI211_X1 g750(.A(new_n950_), .B(new_n951_), .C1(new_n397_), .C2(new_n947_), .ZN(G1348gat));
  AND2_X1   g751(.A1(new_n872_), .A2(new_n946_), .ZN(new_n953_));
  AOI21_X1  g752(.A(G176gat), .B1(new_n953_), .B2(new_n641_), .ZN(new_n954_));
  NAND4_X1  g753(.A1(new_n882_), .A2(G176gat), .A3(new_n641_), .A4(new_n946_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n955_), .A2(KEYINPUT124), .ZN(new_n956_));
  OR2_X1    g755(.A1(new_n955_), .A2(KEYINPUT124), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n954_), .B1(new_n956_), .B2(new_n957_), .ZN(G1349gat));
  NOR2_X1   g757(.A1(new_n608_), .A2(new_n242_), .ZN(new_n959_));
  NAND3_X1  g758(.A1(new_n882_), .A2(new_n612_), .A3(new_n946_), .ZN(new_n960_));
  AOI22_X1  g759(.A1(new_n953_), .A2(new_n959_), .B1(new_n960_), .B2(new_n214_), .ZN(G1350gat));
  NAND2_X1  g760(.A1(new_n392_), .A2(new_n393_), .ZN(new_n962_));
  NAND3_X1  g761(.A1(new_n953_), .A2(new_n962_), .A3(new_n574_), .ZN(new_n963_));
  AND2_X1   g762(.A1(new_n953_), .A2(new_n582_), .ZN(new_n964_));
  OAI21_X1  g763(.A(new_n963_), .B1(new_n964_), .B2(new_n215_), .ZN(G1351gat));
  AND3_X1   g764(.A1(new_n729_), .A2(new_n455_), .A3(new_n464_), .ZN(new_n966_));
  NAND3_X1  g765(.A1(new_n882_), .A2(new_n509_), .A3(new_n966_), .ZN(new_n967_));
  XNOR2_X1  g766(.A(new_n967_), .B(G197gat), .ZN(G1352gat));
  AND2_X1   g767(.A1(new_n882_), .A2(new_n966_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n969_), .A2(new_n641_), .ZN(new_n970_));
  XNOR2_X1  g769(.A(KEYINPUT125), .B(G204gat), .ZN(new_n971_));
  NAND2_X1  g770(.A1(new_n970_), .A2(new_n971_), .ZN(new_n972_));
  AND2_X1   g771(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n973_));
  OAI21_X1  g772(.A(new_n972_), .B1(new_n970_), .B2(new_n973_), .ZN(G1353gat));
  AOI21_X1  g773(.A(new_n608_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n975_));
  XNOR2_X1  g774(.A(new_n975_), .B(KEYINPUT126), .ZN(new_n976_));
  NAND3_X1  g775(.A1(new_n882_), .A2(new_n966_), .A3(new_n976_), .ZN(new_n977_));
  NOR2_X1   g776(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n978_));
  XOR2_X1   g777(.A(new_n977_), .B(new_n978_), .Z(G1354gat));
  NAND2_X1  g778(.A1(new_n969_), .A2(new_n574_), .ZN(new_n980_));
  XOR2_X1   g779(.A(KEYINPUT127), .B(G218gat), .Z(new_n981_));
  NOR2_X1   g780(.A1(new_n856_), .A2(new_n981_), .ZN(new_n982_));
  AOI22_X1  g781(.A1(new_n980_), .A2(new_n981_), .B1(new_n969_), .B2(new_n982_), .ZN(G1355gat));
endmodule


