//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 1 0 0 0 0 1 1 1 1 1 0 1 1 1 0 1 0 0 1 0 0 0 0 1 0 0 1 0 0 0 1 0 0 0 1 1 1 1 0 1 0 1 1 1 1 0 0 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n737_, new_n738_, new_n739_, new_n740_, new_n742_,
    new_n743_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n786_, new_n787_, new_n788_, new_n789_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n909_, new_n911_, new_n912_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n936_, new_n938_, new_n939_, new_n940_, new_n942_, new_n943_,
    new_n944_, new_n946_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n954_, new_n955_;
  INV_X1    g000(.A(KEYINPUT104), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G57gat), .B(G64gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT11), .ZN(new_n204_));
  XOR2_X1   g003(.A(G71gat), .B(G78gat), .Z(new_n205_));
  OR2_X1    g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n205_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n203_), .A2(KEYINPUT11), .ZN(new_n208_));
  OR2_X1    g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  XOR2_X1   g008(.A(G85gat), .B(G92gat), .Z(new_n210_));
  XOR2_X1   g009(.A(KEYINPUT10), .B(G99gat), .Z(new_n211_));
  INV_X1    g010(.A(G106gat), .ZN(new_n212_));
  AOI22_X1  g011(.A1(KEYINPUT9), .A2(new_n210_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G99gat), .A2(G106gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n214_), .B(KEYINPUT6), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G85gat), .A2(G92gat), .ZN(new_n216_));
  OAI211_X1 g015(.A(new_n213_), .B(new_n215_), .C1(KEYINPUT9), .C2(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n218_));
  OR3_X1    g017(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n215_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(new_n210_), .ZN(new_n221_));
  AOI21_X1  g020(.A(KEYINPUT8), .B1(new_n210_), .B2(KEYINPUT65), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n217_), .A2(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n221_), .A2(new_n222_), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n206_), .B(new_n209_), .C1(new_n224_), .C2(new_n225_), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n226_), .A2(KEYINPUT12), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n217_), .A2(new_n223_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n206_), .B1(new_n208_), .B2(new_n207_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n225_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n228_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n231_), .A2(new_n226_), .A3(KEYINPUT12), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n227_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G230gat), .A2(G233gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT64), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n233_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n231_), .A2(new_n226_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(new_n235_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n238_), .A2(KEYINPUT66), .A3(new_n235_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n237_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G120gat), .B(G148gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT5), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G176gat), .B(G204gat), .ZN(new_n246_));
  XOR2_X1   g045(.A(new_n245_), .B(new_n246_), .Z(new_n247_));
  NAND2_X1  g046(.A1(new_n243_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n247_), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n237_), .A2(new_n241_), .A3(new_n242_), .A4(new_n249_), .ZN(new_n250_));
  XOR2_X1   g049(.A(KEYINPUT67), .B(KEYINPUT13), .Z(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n248_), .A2(new_n250_), .A3(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(KEYINPUT67), .A2(KEYINPUT13), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n255_), .B1(new_n248_), .B2(new_n250_), .ZN(new_n256_));
  OR3_X1    g055(.A1(new_n254_), .A2(new_n256_), .A3(KEYINPUT68), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n248_), .A2(new_n250_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n255_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(new_n253_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT68), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n257_), .A2(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G29gat), .B(G36gat), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  XOR2_X1   g064(.A(G43gat), .B(G50gat), .Z(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G43gat), .B(G50gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n264_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT15), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G15gat), .B(G22gat), .ZN(new_n272_));
  INV_X1    g071(.A(G1gat), .ZN(new_n273_));
  INV_X1    g072(.A(G8gat), .ZN(new_n274_));
  OAI21_X1  g073(.A(KEYINPUT14), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n272_), .A2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G1gat), .B(G8gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n271_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n278_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(new_n270_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G229gat), .A2(G233gat), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n279_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n278_), .A2(new_n269_), .A3(new_n267_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n281_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n282_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n283_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT74), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(KEYINPUT75), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT75), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n288_), .A2(new_n289_), .A3(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G113gat), .B(G141gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G169gat), .B(G197gat), .ZN(new_n295_));
  XOR2_X1   g094(.A(new_n294_), .B(new_n295_), .Z(new_n296_));
  NAND3_X1  g095(.A1(new_n291_), .A2(new_n293_), .A3(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n296_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n202_), .B1(new_n263_), .B2(new_n300_), .ZN(new_n301_));
  XOR2_X1   g100(.A(G127gat), .B(G155gat), .Z(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT16), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G183gat), .B(G211gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(KEYINPUT17), .ZN(new_n306_));
  AND2_X1   g105(.A1(G231gat), .A2(G233gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n229_), .B(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT73), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(new_n278_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n309_), .A2(new_n278_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n306_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n312_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT17), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n305_), .A2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n314_), .A2(new_n316_), .A3(new_n310_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n313_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n300_), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n257_), .A2(new_n262_), .A3(KEYINPUT104), .A4(new_n320_), .ZN(new_n321_));
  AND3_X1   g120(.A1(new_n301_), .A2(new_n319_), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G225gat), .A2(G233gat), .ZN(new_n323_));
  INV_X1    g122(.A(G141gat), .ZN(new_n324_));
  INV_X1    g123(.A(G148gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT2), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G141gat), .A2(G148gat), .ZN(new_n328_));
  AOI22_X1  g127(.A1(new_n326_), .A2(KEYINPUT3), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT83), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT83), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n332_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(KEYINPUT82), .B1(new_n326_), .B2(KEYINPUT3), .ZN(new_n335_));
  NOR2_X1   g134(.A1(G141gat), .A2(G148gat), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT82), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT3), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n336_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n329_), .A2(new_n334_), .A3(new_n335_), .A4(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT81), .ZN(new_n341_));
  INV_X1    g140(.A(G155gat), .ZN(new_n342_));
  INV_X1    g141(.A(G162gat), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n341_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(KEYINPUT81), .B1(G155gat), .B2(G162gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G155gat), .A2(G162gat), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n340_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n347_), .A2(KEYINPUT1), .ZN(new_n350_));
  OR2_X1    g149(.A1(new_n347_), .A2(KEYINPUT1), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n346_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  AND2_X1   g151(.A1(new_n326_), .A2(new_n328_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G113gat), .B(G120gat), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G127gat), .B(G134gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(KEYINPUT79), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n357_), .A2(KEYINPUT79), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n356_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  OR2_X1    g160(.A1(new_n357_), .A2(KEYINPUT79), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n362_), .A2(new_n358_), .A3(new_n355_), .ZN(new_n363_));
  AOI22_X1  g162(.A1(new_n349_), .A2(new_n354_), .B1(new_n361_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT4), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n323_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n349_), .A2(new_n354_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n361_), .A2(new_n363_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  AOI22_X1  g168(.A1(new_n340_), .A2(new_n348_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n370_), .A2(new_n363_), .A3(new_n361_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n369_), .A2(new_n371_), .A3(KEYINPUT4), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n366_), .A2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n369_), .A2(new_n371_), .A3(new_n323_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G1gat), .B(G29gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT99), .B(G85gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(KEYINPUT0), .B(G57gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n375_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT103), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n373_), .A2(new_n374_), .A3(new_n380_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n382_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n375_), .A2(KEYINPUT103), .A3(new_n381_), .ZN(new_n386_));
  AND2_X1   g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  AND2_X1   g186(.A1(G183gat), .A2(G190gat), .ZN(new_n388_));
  AND2_X1   g187(.A1(KEYINPUT77), .A2(KEYINPUT23), .ZN(new_n389_));
  NOR2_X1   g188(.A1(KEYINPUT77), .A2(KEYINPUT23), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n388_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(G183gat), .A2(G190gat), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n391_), .A2(new_n393_), .A3(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT22), .ZN(new_n397_));
  INV_X1    g196(.A(G169gat), .ZN(new_n398_));
  INV_X1    g197(.A(G176gat), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n397_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n396_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(G183gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(KEYINPUT25), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT25), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(G183gat), .ZN(new_n408_));
  INV_X1    g207(.A(G190gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT26), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT26), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(G190gat), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n406_), .A2(new_n408_), .A3(new_n410_), .A4(new_n412_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(G169gat), .A2(G176gat), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT24), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  OR2_X1    g215(.A1(KEYINPUT77), .A2(KEYINPUT23), .ZN(new_n417_));
  NAND2_X1  g216(.A1(KEYINPUT77), .A2(KEYINPUT23), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n388_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G183gat), .A2(G190gat), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n420_), .A2(KEYINPUT23), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n413_), .B(new_n416_), .C1(new_n419_), .C2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G169gat), .A2(G176gat), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT76), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n398_), .A2(new_n399_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT76), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n427_), .A2(new_n428_), .A3(KEYINPUT24), .A4(new_n423_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n426_), .A2(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n404_), .B1(new_n422_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G71gat), .B(G99gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(G43gat), .ZN(new_n434_));
  OR2_X1    g233(.A1(new_n432_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n432_), .A2(new_n434_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G227gat), .A2(G233gat), .ZN(new_n438_));
  INV_X1    g237(.A(G15gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n438_), .B(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n437_), .A2(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(KEYINPUT78), .B(KEYINPUT30), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n435_), .A2(new_n440_), .A3(new_n436_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n442_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT80), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n443_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n447_));
  OAI21_X1  g246(.A(KEYINPUT31), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n447_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT31), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n449_), .A2(KEYINPUT80), .A3(new_n450_), .A4(new_n445_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n448_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(new_n368_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n448_), .A2(new_n451_), .A3(new_n363_), .A4(new_n361_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n385_), .A2(new_n386_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G22gat), .B(G50gat), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(KEYINPUT85), .B(KEYINPUT28), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(KEYINPUT86), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT29), .ZN(new_n462_));
  AOI21_X1  g261(.A(KEYINPUT84), .B1(new_n370_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n370_), .A2(KEYINPUT84), .A3(new_n462_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n461_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n465_), .ZN(new_n467_));
  NOR3_X1   g266(.A1(new_n467_), .A2(new_n463_), .A3(new_n460_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n458_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n460_), .B1(new_n467_), .B2(new_n463_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n464_), .A2(new_n465_), .A3(new_n461_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n470_), .A2(new_n471_), .A3(new_n457_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n469_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(G233gat), .ZN(new_n474_));
  INV_X1    g273(.A(G228gat), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n474_), .B1(KEYINPUT87), .B2(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n476_), .B1(KEYINPUT87), .B2(new_n475_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G197gat), .B(G204gat), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT21), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(G218gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(G211gat), .ZN(new_n482_));
  INV_X1    g281(.A(G211gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(G218gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n482_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(G197gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(G204gat), .ZN(new_n488_));
  INV_X1    g287(.A(G204gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(G197gat), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT88), .ZN(new_n491_));
  AND3_X1   g290(.A1(new_n488_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n487_), .A2(KEYINPUT88), .A3(G204gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(KEYINPUT21), .ZN(new_n494_));
  OAI211_X1 g293(.A(new_n480_), .B(new_n486_), .C1(new_n492_), .C2(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n479_), .B1(new_n488_), .B2(new_n490_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n496_), .A2(KEYINPUT89), .A3(new_n485_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(KEYINPUT89), .B1(new_n496_), .B2(new_n485_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n495_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT90), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n477_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n500_), .B1(new_n370_), .B2(new_n462_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  OAI221_X1 g303(.A(new_n500_), .B1(new_n501_), .B2(new_n477_), .C1(new_n370_), .C2(new_n462_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G78gat), .B(G106gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT91), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n506_), .A2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n504_), .A2(new_n505_), .A3(new_n508_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n473_), .A2(new_n512_), .ZN(new_n513_));
  OR2_X1    g312(.A1(new_n511_), .A2(KEYINPUT92), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n506_), .A2(new_n507_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n511_), .A2(KEYINPUT92), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n514_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n513_), .B1(new_n473_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G226gat), .A2(G233gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT19), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n488_), .A2(new_n490_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n522_), .A2(new_n485_), .A3(KEYINPUT21), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT89), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  OAI211_X1 g324(.A(KEYINPUT21), .B(new_n493_), .C1(new_n522_), .C2(KEYINPUT88), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n485_), .B1(new_n479_), .B2(new_n478_), .ZN(new_n527_));
  AOI22_X1  g326(.A1(new_n525_), .A2(new_n497_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT93), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n413_), .A2(new_n416_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n427_), .A2(KEYINPUT24), .A3(new_n423_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n391_), .A2(new_n531_), .A3(new_n395_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n529_), .B1(new_n530_), .B2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT25), .B(G183gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(KEYINPUT26), .B(G190gat), .ZN(new_n535_));
  AOI22_X1  g334(.A1(new_n534_), .A2(new_n535_), .B1(new_n415_), .B2(new_n414_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(KEYINPUT77), .B(KEYINPUT23), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n394_), .B1(new_n537_), .B2(new_n388_), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n536_), .A2(KEYINPUT93), .A3(new_n538_), .A4(new_n531_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n533_), .A2(new_n539_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n393_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT94), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n402_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n403_), .A2(KEYINPUT94), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n541_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n528_), .B1(new_n540_), .B2(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(KEYINPUT20), .B1(new_n500_), .B2(new_n431_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n521_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n500_), .A2(new_n431_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT95), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n500_), .A2(new_n431_), .A3(KEYINPUT95), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n551_), .A2(KEYINPUT20), .A3(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n540_), .A2(new_n528_), .A3(new_n545_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n521_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n548_), .B1(new_n553_), .B2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G64gat), .B(G92gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT97), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G8gat), .B(G36gat), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  OR2_X1    g360(.A1(new_n559_), .A2(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n559_), .A2(new_n561_), .ZN(new_n564_));
  AND3_X1   g363(.A1(new_n562_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n563_), .B1(new_n562_), .B2(new_n564_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n557_), .A2(new_n568_), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n548_), .B(new_n567_), .C1(new_n553_), .C2(new_n556_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n569_), .A2(KEYINPUT98), .A3(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT27), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT98), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n557_), .A2(new_n573_), .A3(new_n568_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n571_), .A2(new_n572_), .A3(new_n574_), .ZN(new_n575_));
  NOR3_X1   g374(.A1(new_n546_), .A2(new_n547_), .A3(new_n521_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n536_), .A2(new_n538_), .A3(new_n531_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n545_), .A2(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n500_), .B1(new_n578_), .B2(KEYINPUT102), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n579_), .B1(KEYINPUT102), .B2(new_n578_), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n552_), .A2(KEYINPUT20), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n580_), .A2(new_n551_), .A3(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n576_), .B1(new_n582_), .B2(new_n521_), .ZN(new_n583_));
  OAI211_X1 g382(.A(KEYINPUT27), .B(new_n570_), .C1(new_n583_), .C2(new_n567_), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n575_), .A2(new_n584_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n455_), .A2(new_n456_), .A3(new_n519_), .A4(new_n585_), .ZN(new_n586_));
  AND4_X1   g385(.A1(new_n456_), .A2(new_n518_), .A3(new_n575_), .A4(new_n584_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n570_), .A2(KEYINPUT98), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n581_), .A2(new_n555_), .A3(new_n551_), .A4(new_n554_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n567_), .B1(new_n589_), .B2(new_n548_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n574_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT33), .ZN(new_n594_));
  OAI211_X1 g393(.A(new_n372_), .B(new_n323_), .C1(KEYINPUT4), .C2(new_n369_), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n369_), .A2(new_n371_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n323_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n380_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  AOI22_X1  g397(.A1(new_n384_), .A2(new_n594_), .B1(new_n595_), .B2(new_n598_), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n373_), .A2(KEYINPUT33), .A3(new_n374_), .A4(new_n380_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT100), .ZN(new_n601_));
  AND2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n600_), .A2(new_n601_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n599_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(KEYINPUT101), .B1(new_n593_), .B2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n571_), .A2(new_n574_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n600_), .B(new_n601_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT101), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n606_), .A2(new_n607_), .A3(new_n608_), .A4(new_n599_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n567_), .A2(KEYINPUT32), .ZN(new_n610_));
  MUX2_X1   g409(.A(new_n583_), .B(new_n557_), .S(new_n610_), .Z(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(new_n387_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n605_), .A2(new_n609_), .A3(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n587_), .B1(new_n613_), .B2(new_n519_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n586_), .B1(new_n614_), .B2(new_n455_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G190gat), .B(G218gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G134gat), .B(G162gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n619_), .B(KEYINPUT36), .Z(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n228_), .A2(new_n270_), .A3(new_n230_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n271_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n624_));
  NAND2_X1  g423(.A1(G232gat), .A2(G233gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n627_), .A2(KEYINPUT35), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n622_), .A2(new_n623_), .A3(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n629_), .A2(KEYINPUT35), .A3(new_n627_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n627_), .A2(KEYINPUT35), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n622_), .A2(new_n623_), .A3(new_n631_), .A4(new_n628_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT72), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n621_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n635_), .B1(new_n634_), .B2(new_n633_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n619_), .A2(KEYINPUT36), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n630_), .A2(new_n637_), .A3(new_n632_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n636_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n616_), .A2(new_n640_), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n322_), .A2(new_n387_), .A3(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n642_), .A2(new_n273_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT38), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT69), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n263_), .A2(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n257_), .A2(new_n262_), .A3(KEYINPUT69), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n455_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n606_), .A2(new_n607_), .A3(new_n599_), .ZN(new_n650_));
  AOI22_X1  g449(.A1(new_n650_), .A2(KEYINPUT101), .B1(new_n611_), .B2(new_n387_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n518_), .B1(new_n651_), .B2(new_n609_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n649_), .B1(new_n652_), .B2(new_n587_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n300_), .B1(new_n653_), .B2(new_n586_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT37), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n636_), .A2(new_n655_), .A3(new_n638_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n620_), .B(KEYINPUT71), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n633_), .A2(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n655_), .B1(new_n658_), .B2(new_n638_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n656_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n662_), .A2(new_n318_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n648_), .A2(new_n654_), .A3(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n665_), .A2(new_n273_), .A3(new_n387_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n643_), .B1(new_n644_), .B2(new_n666_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n667_), .B1(new_n644_), .B2(new_n666_), .ZN(G1324gat));
  INV_X1    g467(.A(new_n585_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n322_), .A2(new_n669_), .A3(new_n641_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT39), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n670_), .A2(new_n671_), .A3(G8gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n671_), .B1(new_n670_), .B2(G8gat), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n669_), .A2(new_n274_), .ZN(new_n674_));
  OAI22_X1  g473(.A1(new_n672_), .A2(new_n673_), .B1(new_n664_), .B2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT40), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  OAI221_X1 g476(.A(KEYINPUT40), .B1(new_n664_), .B2(new_n674_), .C1(new_n672_), .C2(new_n673_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1325gat));
  NAND3_X1  g478(.A1(new_n665_), .A2(new_n439_), .A3(new_n455_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n322_), .A2(new_n455_), .A3(new_n641_), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n681_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(KEYINPUT41), .B1(new_n681_), .B2(G15gat), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n680_), .B1(new_n682_), .B2(new_n683_), .ZN(G1326gat));
  NAND3_X1  g483(.A1(new_n322_), .A2(new_n518_), .A3(new_n641_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT42), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n685_), .A2(new_n686_), .A3(G22gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n686_), .B1(new_n685_), .B2(G22gat), .ZN(new_n688_));
  OR2_X1    g487(.A1(new_n519_), .A2(G22gat), .ZN(new_n689_));
  OAI22_X1  g488(.A1(new_n687_), .A2(new_n688_), .B1(new_n664_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT105), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  OAI221_X1 g491(.A(KEYINPUT105), .B1(new_n664_), .B2(new_n689_), .C1(new_n687_), .C2(new_n688_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1327gat));
  NAND2_X1  g493(.A1(new_n640_), .A2(new_n318_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n263_), .A2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n654_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(G29gat), .B1(new_n698_), .B2(new_n387_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n661_), .A2(KEYINPUT43), .ZN(new_n701_));
  AND3_X1   g500(.A1(new_n615_), .A2(KEYINPUT107), .A3(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT43), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT106), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n656_), .A2(new_n704_), .A3(new_n660_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n704_), .B1(new_n656_), .B2(new_n660_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n703_), .B1(new_n615_), .B2(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(KEYINPUT107), .B1(new_n615_), .B2(new_n701_), .ZN(new_n710_));
  NOR3_X1   g509(.A1(new_n702_), .A2(new_n709_), .A3(new_n710_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n301_), .A2(new_n318_), .A3(new_n321_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n700_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  AND3_X1   g512(.A1(new_n301_), .A2(new_n318_), .A3(new_n321_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n707_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(new_n705_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n716_), .B1(new_n653_), .B2(new_n586_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n701_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n718_), .B1(new_n653_), .B2(new_n586_), .ZN(new_n719_));
  OAI22_X1  g518(.A1(new_n717_), .A2(new_n703_), .B1(new_n719_), .B2(KEYINPUT107), .ZN(new_n720_));
  OAI211_X1 g519(.A(new_n714_), .B(KEYINPUT44), .C1(new_n720_), .C2(new_n702_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n713_), .A2(new_n721_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n387_), .A2(G29gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n699_), .B1(new_n722_), .B2(new_n723_), .ZN(G1328gat));
  NAND3_X1  g523(.A1(new_n713_), .A2(new_n669_), .A3(new_n721_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(G36gat), .ZN(new_n726_));
  OR2_X1    g525(.A1(new_n669_), .A2(KEYINPUT108), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n669_), .A2(KEYINPUT108), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  NOR3_X1   g528(.A1(new_n697_), .A2(G36gat), .A3(new_n729_), .ZN(new_n730_));
  XOR2_X1   g529(.A(new_n730_), .B(KEYINPUT45), .Z(new_n731_));
  NAND2_X1  g530(.A1(new_n726_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT46), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n726_), .A2(KEYINPUT46), .A3(new_n731_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(G1329gat));
  NAND4_X1  g535(.A1(new_n713_), .A2(new_n721_), .A3(G43gat), .A4(new_n455_), .ZN(new_n737_));
  INV_X1    g536(.A(G43gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n738_), .B1(new_n697_), .B2(new_n649_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g540(.A(G50gat), .B1(new_n698_), .B2(new_n518_), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n518_), .A2(G50gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n722_), .B2(new_n743_), .ZN(G1331gat));
  INV_X1    g543(.A(new_n648_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n299_), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n746_), .A2(new_n317_), .A3(new_n313_), .A4(new_n297_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n745_), .A2(new_n641_), .A3(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(G57gat), .B1(new_n749_), .B2(new_n456_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n616_), .A2(new_n320_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n751_), .A2(new_n263_), .A3(new_n663_), .ZN(new_n752_));
  OR2_X1    g551(.A1(new_n456_), .A2(G57gat), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n750_), .B1(new_n752_), .B2(new_n753_), .ZN(G1332gat));
  OR3_X1    g553(.A1(new_n752_), .A2(G64gat), .A3(new_n729_), .ZN(new_n755_));
  OR2_X1    g554(.A1(new_n749_), .A2(new_n729_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT48), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n756_), .A2(new_n757_), .A3(G64gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n757_), .B1(new_n756_), .B2(G64gat), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n755_), .B1(new_n758_), .B2(new_n759_), .ZN(G1333gat));
  OR3_X1    g559(.A1(new_n752_), .A2(G71gat), .A3(new_n649_), .ZN(new_n761_));
  OR2_X1    g560(.A1(new_n749_), .A2(new_n649_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT49), .ZN(new_n763_));
  AND3_X1   g562(.A1(new_n762_), .A2(new_n763_), .A3(G71gat), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n762_), .B2(G71gat), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n761_), .B1(new_n764_), .B2(new_n765_), .ZN(G1334gat));
  OR3_X1    g565(.A1(new_n752_), .A2(G78gat), .A3(new_n519_), .ZN(new_n767_));
  OR2_X1    g566(.A1(new_n749_), .A2(new_n519_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT50), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n768_), .A2(new_n769_), .A3(G78gat), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n768_), .B2(G78gat), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n767_), .B1(new_n770_), .B2(new_n771_), .ZN(G1335gat));
  INV_X1    g571(.A(G85gat), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n320_), .A2(new_n319_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n263_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT109), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n263_), .A2(KEYINPUT109), .A3(new_n774_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n711_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n773_), .B1(new_n779_), .B2(new_n387_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n695_), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n646_), .A2(new_n647_), .A3(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(new_n751_), .ZN(new_n783_));
  NOR3_X1   g582(.A1(new_n783_), .A2(G85gat), .A3(new_n456_), .ZN(new_n784_));
  OR2_X1    g583(.A1(new_n780_), .A2(new_n784_), .ZN(G1336gat));
  INV_X1    g584(.A(G92gat), .ZN(new_n786_));
  INV_X1    g585(.A(new_n729_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n779_), .B2(new_n787_), .ZN(new_n788_));
  NOR3_X1   g587(.A1(new_n783_), .A2(G92gat), .A3(new_n585_), .ZN(new_n789_));
  OR2_X1    g588(.A1(new_n788_), .A2(new_n789_), .ZN(G1337gat));
  NAND4_X1  g589(.A1(new_n782_), .A2(new_n751_), .A3(new_n455_), .A4(new_n211_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT110), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n791_), .B(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT111), .ZN(new_n794_));
  INV_X1    g593(.A(G99gat), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n795_), .B1(new_n779_), .B2(new_n455_), .ZN(new_n796_));
  OAI21_X1  g595(.A(KEYINPUT51), .B1(new_n794_), .B2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n796_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT51), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n798_), .A2(KEYINPUT111), .A3(new_n799_), .A4(new_n793_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n797_), .A2(new_n800_), .ZN(G1338gat));
  NAND4_X1  g600(.A1(new_n782_), .A2(new_n751_), .A3(new_n212_), .A4(new_n518_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n777_), .A2(new_n778_), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n518_), .B(new_n803_), .C1(new_n720_), .C2(new_n702_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n212_), .B1(KEYINPUT112), .B2(KEYINPUT52), .ZN(new_n805_));
  NOR2_X1   g604(.A1(KEYINPUT112), .A2(KEYINPUT52), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n804_), .A2(new_n805_), .A3(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n806_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n802_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT53), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n811_), .B(new_n802_), .C1(new_n807_), .C2(new_n808_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n812_), .ZN(G1339gat));
  INV_X1    g612(.A(G113gat), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT59), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n250_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT56), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n227_), .A2(new_n235_), .A3(new_n232_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n235_), .B1(new_n227_), .B2(new_n232_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n818_), .B1(new_n819_), .B2(KEYINPUT55), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n821_));
  OAI21_X1  g620(.A(KEYINPUT114), .B1(new_n237_), .B2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT114), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n819_), .A2(new_n823_), .A3(KEYINPUT55), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n820_), .B1(new_n822_), .B2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n817_), .B1(new_n825_), .B2(new_n249_), .ZN(new_n826_));
  AND3_X1   g625(.A1(new_n227_), .A2(new_n235_), .A3(new_n232_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n827_), .B1(new_n237_), .B2(new_n821_), .ZN(new_n828_));
  AND3_X1   g627(.A1(new_n819_), .A2(new_n823_), .A3(KEYINPUT55), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n823_), .B1(new_n819_), .B2(KEYINPUT55), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n828_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n831_), .A2(KEYINPUT56), .A3(new_n247_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n816_), .B1(new_n826_), .B2(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n279_), .A2(new_n281_), .A3(new_n286_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n285_), .A2(new_n282_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n296_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n836_), .B1(new_n288_), .B2(new_n296_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n837_), .B1(new_n248_), .B2(new_n250_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n639_), .B1(new_n833_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT57), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n250_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n842_), .A2(new_n837_), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n825_), .A2(new_n817_), .A3(new_n249_), .ZN(new_n844_));
  AOI21_X1  g643(.A(KEYINPUT56), .B1(new_n831_), .B2(new_n247_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n843_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT58), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  OAI211_X1 g647(.A(KEYINPUT58), .B(new_n843_), .C1(new_n844_), .C2(new_n845_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n848_), .A2(new_n662_), .A3(new_n849_), .ZN(new_n850_));
  OAI211_X1 g649(.A(KEYINPUT57), .B(new_n639_), .C1(new_n833_), .C2(new_n838_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n841_), .A2(new_n850_), .A3(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(KEYINPUT113), .B1(new_n261_), .B2(new_n748_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT113), .ZN(new_n854_));
  AOI211_X1 g653(.A(new_n854_), .B(new_n747_), .C1(new_n260_), .C2(new_n253_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n661_), .B1(new_n853_), .B2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(KEYINPUT54), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n254_), .A2(new_n256_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n854_), .B1(new_n858_), .B2(new_n747_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n261_), .A2(new_n748_), .A3(KEYINPUT113), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT54), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n861_), .A2(new_n862_), .A3(new_n661_), .ZN(new_n863_));
  AOI22_X1  g662(.A1(new_n852_), .A2(new_n318_), .B1(new_n857_), .B2(new_n863_), .ZN(new_n864_));
  NOR4_X1   g663(.A1(new_n649_), .A2(new_n456_), .A3(new_n518_), .A4(new_n669_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(KEYINPUT115), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n815_), .B1(new_n864_), .B2(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n661_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n869_));
  AOI22_X1  g668(.A1(new_n849_), .A2(new_n869_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n319_), .B1(new_n870_), .B2(new_n851_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n862_), .B1(new_n861_), .B2(new_n661_), .ZN(new_n872_));
  AOI211_X1 g671(.A(KEYINPUT54), .B(new_n662_), .C1(new_n859_), .C2(new_n860_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  OAI211_X1 g673(.A(KEYINPUT59), .B(new_n866_), .C1(new_n871_), .C2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n868_), .A2(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n814_), .B1(new_n876_), .B2(new_n320_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n864_), .A2(new_n867_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n320_), .A2(new_n814_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  OAI21_X1  g680(.A(KEYINPUT116), .B1(new_n877_), .B2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT116), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n300_), .B1(new_n868_), .B2(new_n875_), .ZN(new_n884_));
  OAI221_X1 g683(.A(new_n883_), .B1(new_n879_), .B2(new_n880_), .C1(new_n884_), .C2(new_n814_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n882_), .A2(new_n885_), .ZN(G1340gat));
  INV_X1    g685(.A(G120gat), .ZN(new_n887_));
  INV_X1    g686(.A(new_n263_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n888_), .B2(KEYINPUT60), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n878_), .B(new_n889_), .C1(KEYINPUT60), .C2(new_n887_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n648_), .B1(new_n868_), .B2(new_n875_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n891_), .B2(new_n887_), .ZN(G1341gat));
  AOI21_X1  g691(.A(G127gat), .B1(new_n878_), .B2(new_n319_), .ZN(new_n893_));
  OR2_X1    g692(.A1(new_n893_), .A2(KEYINPUT117), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(KEYINPUT117), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n319_), .A2(G127gat), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(KEYINPUT118), .ZN(new_n897_));
  AOI22_X1  g696(.A1(new_n894_), .A2(new_n895_), .B1(new_n876_), .B2(new_n897_), .ZN(G1342gat));
  AOI21_X1  g697(.A(G134gat), .B1(new_n878_), .B2(new_n640_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n662_), .A2(G134gat), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(KEYINPUT119), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n899_), .B1(new_n876_), .B2(new_n901_), .ZN(G1343gat));
  INV_X1    g701(.A(new_n864_), .ZN(new_n903_));
  NAND4_X1  g702(.A1(new_n729_), .A2(new_n387_), .A3(new_n518_), .A4(new_n649_), .ZN(new_n904_));
  XOR2_X1   g703(.A(new_n904_), .B(KEYINPUT120), .Z(new_n905_));
  NAND2_X1  g704(.A1(new_n903_), .A2(new_n905_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n906_), .A2(new_n300_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(new_n324_), .ZN(G1344gat));
  NOR2_X1   g707(.A1(new_n906_), .A2(new_n648_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(new_n325_), .ZN(G1345gat));
  NOR2_X1   g709(.A1(new_n906_), .A2(new_n318_), .ZN(new_n911_));
  XOR2_X1   g710(.A(KEYINPUT61), .B(G155gat), .Z(new_n912_));
  XNOR2_X1  g711(.A(new_n911_), .B(new_n912_), .ZN(G1346gat));
  NOR3_X1   g712(.A1(new_n906_), .A2(new_n343_), .A3(new_n716_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n343_), .B1(new_n906_), .B2(new_n639_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(KEYINPUT121), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT121), .ZN(new_n917_));
  OAI211_X1 g716(.A(new_n917_), .B(new_n343_), .C1(new_n906_), .C2(new_n639_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n914_), .B1(new_n916_), .B2(new_n918_), .ZN(G1347gat));
  NOR4_X1   g718(.A1(new_n729_), .A2(new_n387_), .A3(new_n518_), .A4(new_n649_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n903_), .A2(new_n320_), .A3(new_n920_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(KEYINPUT122), .B(KEYINPUT62), .ZN(new_n922_));
  AND3_X1   g721(.A1(new_n921_), .A2(G169gat), .A3(new_n922_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n922_), .B1(new_n921_), .B2(G169gat), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n903_), .A2(new_n920_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(KEYINPUT22), .B(G169gat), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n320_), .A2(new_n926_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(KEYINPUT123), .ZN(new_n928_));
  OAI22_X1  g727(.A1(new_n923_), .A2(new_n924_), .B1(new_n925_), .B2(new_n928_), .ZN(G1348gat));
  INV_X1    g728(.A(new_n925_), .ZN(new_n930_));
  AOI21_X1  g729(.A(G176gat), .B1(new_n930_), .B2(new_n263_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n745_), .A2(G176gat), .ZN(new_n932_));
  OR3_X1    g731(.A1(new_n925_), .A2(KEYINPUT124), .A3(new_n932_), .ZN(new_n933_));
  OAI21_X1  g732(.A(KEYINPUT124), .B1(new_n925_), .B2(new_n932_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n931_), .B1(new_n933_), .B2(new_n934_), .ZN(G1349gat));
  NOR2_X1   g734(.A1(new_n925_), .A2(new_n318_), .ZN(new_n936_));
  MUX2_X1   g735(.A(G183gat), .B(new_n534_), .S(new_n936_), .Z(G1350gat));
  OAI21_X1  g736(.A(G190gat), .B1(new_n925_), .B2(new_n661_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n640_), .A2(new_n535_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n939_), .B(KEYINPUT125), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n938_), .B1(new_n925_), .B2(new_n940_), .ZN(G1351gat));
  NOR4_X1   g740(.A1(new_n729_), .A2(new_n387_), .A3(new_n519_), .A4(new_n455_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n903_), .A2(new_n942_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n943_), .A2(new_n300_), .ZN(new_n944_));
  XNOR2_X1  g743(.A(new_n944_), .B(new_n487_), .ZN(G1352gat));
  NOR2_X1   g744(.A1(new_n943_), .A2(new_n648_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(new_n489_), .ZN(G1353gat));
  INV_X1    g746(.A(new_n943_), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n318_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n949_));
  XNOR2_X1  g748(.A(new_n949_), .B(KEYINPUT126), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n948_), .A2(new_n950_), .ZN(new_n951_));
  OR2_X1    g750(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n952_));
  XNOR2_X1  g751(.A(new_n951_), .B(new_n952_), .ZN(G1354gat));
  OAI21_X1  g752(.A(G218gat), .B1(new_n943_), .B2(new_n661_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n640_), .A2(new_n481_), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n954_), .B1(new_n943_), .B2(new_n955_), .ZN(G1355gat));
endmodule


