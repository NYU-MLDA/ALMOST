//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 1 0 1 1 1 0 0 0 1 1 0 1 0 0 0 0 0 1 0 0 0 1 0 0 1 1 0 0 1 1 1 0 1 1 1 0 1 0 0 0 1 0 1 1 0 1 1 0 0 1 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n707_, new_n708_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n721_, new_n722_, new_n723_, new_n725_, new_n726_, new_n727_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n859_, new_n860_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n867_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n890_, new_n892_, new_n893_, new_n894_,
    new_n896_, new_n897_, new_n898_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G85gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT0), .B(G57gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  NAND2_X1  g004(.A1(G225gat), .A2(G233gat), .ZN(new_n206_));
  XOR2_X1   g005(.A(G155gat), .B(G162gat), .Z(new_n207_));
  INV_X1    g006(.A(KEYINPUT1), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT87), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G141gat), .A2(G148gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n209_), .A2(new_n212_), .A3(new_n213_), .A4(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT3), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n210_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT2), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n213_), .A2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n217_), .A2(new_n219_), .A3(new_n220_), .A4(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(new_n207_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n215_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  XOR2_X1   g024(.A(G127gat), .B(G134gat), .Z(new_n226_));
  XOR2_X1   g025(.A(G113gat), .B(G120gat), .Z(new_n227_));
  XOR2_X1   g026(.A(new_n226_), .B(new_n227_), .Z(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n225_), .A2(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT102), .B1(new_n224_), .B2(new_n228_), .ZN(new_n231_));
  OR2_X1    g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n230_), .A2(new_n231_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT4), .ZN(new_n235_));
  NOR3_X1   g034(.A1(new_n225_), .A2(new_n229_), .A3(KEYINPUT4), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n206_), .B1(new_n235_), .B2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n206_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n234_), .A2(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n205_), .B1(new_n238_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT4), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n242_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n239_), .B1(new_n243_), .B2(new_n236_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n205_), .ZN(new_n245_));
  OAI211_X1 g044(.A(new_n244_), .B(new_n245_), .C1(new_n239_), .C2(new_n234_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n241_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G226gat), .A2(G233gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT19), .ZN(new_n250_));
  NOR2_X1   g049(.A1(G183gat), .A2(G190gat), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT23), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G183gat), .A2(G190gat), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n251_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n254_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT22), .B(G169gat), .ZN(new_n256_));
  INV_X1    g055(.A(G176gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G169gat), .A2(G176gat), .ZN(new_n259_));
  AND3_X1   g058(.A1(new_n258_), .A2(KEYINPUT100), .A3(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(KEYINPUT100), .B1(new_n258_), .B2(new_n259_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n255_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT101), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  OAI211_X1 g063(.A(KEYINPUT101), .B(new_n255_), .C1(new_n260_), .C2(new_n261_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n253_), .B(KEYINPUT23), .ZN(new_n266_));
  NOR2_X1   g065(.A1(G169gat), .A2(G176gat), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT24), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  AND3_X1   g068(.A1(new_n266_), .A2(KEYINPUT99), .A3(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(KEYINPUT99), .B1(new_n266_), .B2(new_n269_), .ZN(new_n271_));
  OR2_X1    g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT81), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n267_), .B(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n259_), .A2(KEYINPUT24), .ZN(new_n275_));
  OR2_X1    g074(.A1(new_n275_), .A2(KEYINPUT98), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(KEYINPUT98), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n274_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT25), .B(G183gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT26), .B(G190gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n278_), .A2(new_n281_), .ZN(new_n282_));
  AOI22_X1  g081(.A1(new_n264_), .A2(new_n265_), .B1(new_n272_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(G197gat), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT90), .B1(new_n284_), .B2(G204gat), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT90), .ZN(new_n286_));
  INV_X1    g085(.A(G204gat), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n286_), .A2(new_n287_), .A3(G197gat), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n285_), .B(new_n288_), .C1(G197gat), .C2(new_n287_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT21), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G211gat), .B(G218gat), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT91), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n292_), .B1(new_n284_), .B2(G204gat), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n287_), .A2(KEYINPUT91), .A3(G197gat), .ZN(new_n294_));
  OAI211_X1 g093(.A(new_n293_), .B(new_n294_), .C1(G197gat), .C2(new_n287_), .ZN(new_n295_));
  OAI211_X1 g094(.A(new_n290_), .B(new_n291_), .C1(KEYINPUT21), .C2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT21), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n291_), .A2(new_n297_), .ZN(new_n298_));
  AND3_X1   g097(.A1(new_n298_), .A2(new_n295_), .A3(KEYINPUT92), .ZN(new_n299_));
  AOI21_X1  g098(.A(KEYINPUT92), .B1(new_n298_), .B2(new_n295_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n296_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(KEYINPUT20), .B1(new_n283_), .B2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT82), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n258_), .B(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n305_), .A2(new_n259_), .A3(new_n255_), .ZN(new_n306_));
  AND2_X1   g105(.A1(new_n281_), .A2(new_n266_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n274_), .A2(KEYINPUT24), .A3(new_n259_), .ZN(new_n308_));
  OAI211_X1 g107(.A(new_n307_), .B(new_n308_), .C1(KEYINPUT24), .C2(new_n274_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n306_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n301_), .A2(KEYINPUT93), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT93), .ZN(new_n312_));
  OAI211_X1 g111(.A(new_n296_), .B(new_n312_), .C1(new_n299_), .C2(new_n300_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n310_), .B1(new_n311_), .B2(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n250_), .B1(new_n303_), .B2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n283_), .A2(new_n302_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n250_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n311_), .A2(new_n310_), .A3(new_n313_), .ZN(new_n318_));
  NAND4_X1  g117(.A1(new_n316_), .A2(KEYINPUT20), .A3(new_n317_), .A4(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n315_), .A2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G8gat), .B(G36gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT18), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G64gat), .B(G92gat), .ZN(new_n323_));
  XOR2_X1   g122(.A(new_n322_), .B(new_n323_), .Z(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n320_), .A2(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n315_), .A2(new_n324_), .A3(new_n319_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT27), .ZN(new_n329_));
  AND2_X1   g128(.A1(new_n327_), .A2(KEYINPUT27), .ZN(new_n330_));
  OAI211_X1 g129(.A(new_n281_), .B(new_n278_), .C1(new_n270_), .C2(new_n271_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(new_n262_), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT20), .B1(new_n332_), .B2(new_n301_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n318_), .B1(new_n333_), .B2(KEYINPUT104), .ZN(new_n334_));
  AND2_X1   g133(.A1(new_n333_), .A2(KEYINPUT104), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n250_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n311_), .A2(new_n313_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n310_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  OAI211_X1 g138(.A(new_n339_), .B(KEYINPUT20), .C1(new_n302_), .C2(new_n283_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n336_), .B1(new_n250_), .B2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(new_n325_), .ZN(new_n342_));
  AOI22_X1  g141(.A1(new_n328_), .A2(new_n329_), .B1(new_n330_), .B2(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n224_), .A2(KEYINPUT29), .ZN(new_n344_));
  XOR2_X1   g143(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(KEYINPUT89), .ZN(new_n346_));
  AND2_X1   g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n344_), .A2(new_n346_), .ZN(new_n348_));
  XOR2_X1   g147(.A(G22gat), .B(G50gat), .Z(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  OR3_X1    g149(.A1(new_n347_), .A2(new_n348_), .A3(new_n350_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n350_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n224_), .A2(KEYINPUT29), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G228gat), .A2(G233gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(KEYINPUT94), .B1(new_n337_), .B2(new_n356_), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n354_), .A2(new_n355_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT94), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n358_), .A2(new_n359_), .A3(new_n311_), .A4(new_n313_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n357_), .A2(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n355_), .B1(new_n301_), .B2(new_n354_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n361_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT96), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G78gat), .B(G106gat), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n364_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n362_), .B1(new_n357_), .B2(new_n360_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n366_), .ZN(new_n369_));
  OAI21_X1  g168(.A(KEYINPUT96), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  AND2_X1   g169(.A1(new_n367_), .A2(new_n370_), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n368_), .A2(KEYINPUT95), .A3(new_n369_), .ZN(new_n372_));
  AOI21_X1  g171(.A(KEYINPUT95), .B1(new_n368_), .B2(new_n369_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n353_), .B1(new_n371_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT97), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n353_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n377_));
  AOI211_X1 g176(.A(new_n366_), .B(new_n362_), .C1(new_n357_), .C2(new_n360_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n376_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n364_), .A2(new_n366_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n368_), .A2(new_n369_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n380_), .A2(KEYINPUT97), .A3(new_n353_), .A4(new_n381_), .ZN(new_n382_));
  AND2_X1   g181(.A1(new_n379_), .A2(new_n382_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n248_), .B(new_n343_), .C1(new_n375_), .C2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(KEYINPUT105), .ZN(new_n385_));
  INV_X1    g184(.A(new_n373_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n378_), .A2(KEYINPUT95), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n386_), .A2(new_n387_), .A3(new_n367_), .A4(new_n370_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n353_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n379_), .A2(new_n382_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT105), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n392_), .A2(new_n393_), .A3(new_n248_), .A4(new_n343_), .ZN(new_n394_));
  NOR3_X1   g193(.A1(new_n243_), .A2(new_n239_), .A3(new_n236_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n234_), .A2(new_n239_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(new_n245_), .ZN(new_n397_));
  OAI21_X1  g196(.A(KEYINPUT33), .B1(new_n395_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n241_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n328_), .ZN(new_n400_));
  OAI211_X1 g199(.A(KEYINPUT33), .B(new_n205_), .C1(new_n238_), .C2(new_n240_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n399_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n324_), .A2(KEYINPUT32), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n320_), .A2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(KEYINPUT103), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n341_), .A2(new_n403_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n247_), .A2(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n402_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n375_), .A2(new_n383_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n385_), .A2(new_n394_), .A3(new_n410_), .ZN(new_n411_));
  XOR2_X1   g210(.A(G15gat), .B(G43gat), .Z(new_n412_));
  XNOR2_X1  g211(.A(new_n412_), .B(KEYINPUT84), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n310_), .B(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G227gat), .A2(G233gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT85), .ZN(new_n416_));
  XOR2_X1   g215(.A(G71gat), .B(G99gat), .Z(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  XOR2_X1   g217(.A(KEYINPUT83), .B(KEYINPUT30), .Z(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n414_), .B(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT86), .ZN(new_n422_));
  AND2_X1   g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n228_), .B(KEYINPUT31), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n423_), .A2(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n424_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n426_), .B1(new_n423_), .B2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n411_), .A2(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n428_), .A2(new_n247_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n409_), .A2(new_n430_), .A3(new_n343_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT106), .ZN(new_n432_));
  INV_X1    g231(.A(new_n343_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n392_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT106), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n434_), .A2(new_n435_), .A3(new_n430_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n432_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n429_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT8), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT67), .ZN(new_n440_));
  NOR2_X1   g239(.A1(G99gat), .A2(G106gat), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT65), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT7), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n441_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(G99gat), .ZN(new_n447_));
  INV_X1    g246(.A(G106gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  AND2_X1   g248(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n440_), .B1(new_n446_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G99gat), .A2(G106gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT6), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT6), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n455_), .A2(G99gat), .A3(G106gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n454_), .A2(new_n456_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n449_), .B1(new_n450_), .B2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n441_), .A2(new_n445_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n459_), .A2(KEYINPUT67), .A3(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n452_), .A2(new_n457_), .A3(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G85gat), .B(G92gat), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n439_), .B1(new_n462_), .B2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n459_), .A2(new_n457_), .A3(new_n460_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT66), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n463_), .A2(KEYINPUT8), .ZN(new_n468_));
  AND3_X1   g267(.A1(new_n466_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n467_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT70), .B1(new_n465_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n466_), .A2(new_n468_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT66), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n466_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT70), .ZN(new_n477_));
  INV_X1    g276(.A(new_n457_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n459_), .A2(new_n460_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n478_), .B1(new_n479_), .B2(new_n440_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n463_), .B1(new_n480_), .B2(new_n461_), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n476_), .B(new_n477_), .C1(new_n439_), .C2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n472_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n464_), .A2(KEYINPUT9), .ZN(new_n484_));
  XOR2_X1   g283(.A(KEYINPUT10), .B(G99gat), .Z(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(new_n448_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(KEYINPUT64), .B(G92gat), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT9), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n487_), .A2(new_n488_), .A3(G85gat), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n484_), .A2(new_n486_), .A3(new_n457_), .A4(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n483_), .A2(new_n490_), .ZN(new_n491_));
  XOR2_X1   g290(.A(G71gat), .B(G78gat), .Z(new_n492_));
  XNOR2_X1  g291(.A(G57gat), .B(G64gat), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n492_), .B1(KEYINPUT11), .B2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT69), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n493_), .A2(KEYINPUT11), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n495_), .B(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT12), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n491_), .A2(new_n500_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n476_), .B1(new_n481_), .B2(new_n439_), .ZN(new_n502_));
  AOI21_X1  g301(.A(KEYINPUT68), .B1(new_n502_), .B2(new_n490_), .ZN(new_n503_));
  OAI211_X1 g302(.A(KEYINPUT68), .B(new_n490_), .C1(new_n465_), .C2(new_n471_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n498_), .B1(new_n503_), .B2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n501_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT71), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT68), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n462_), .A2(new_n464_), .ZN(new_n510_));
  AOI22_X1  g309(.A1(new_n510_), .A2(KEYINPUT8), .B1(new_n474_), .B2(new_n475_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n490_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n509_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT69), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n494_), .B(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(new_n497_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n513_), .A2(new_n516_), .A3(new_n504_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n508_), .B1(new_n517_), .B2(new_n499_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n507_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G230gat), .A2(G233gat), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n517_), .A2(new_n508_), .A3(new_n499_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n519_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n506_), .A2(new_n517_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n520_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n522_), .A2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G120gat), .B(G148gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT5), .ZN(new_n528_));
  XOR2_X1   g327(.A(G176gat), .B(G204gat), .Z(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  OR2_X1    g329(.A1(new_n526_), .A2(new_n530_), .ZN(new_n531_));
  XOR2_X1   g330(.A(new_n530_), .B(KEYINPUT72), .Z(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n526_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n531_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(KEYINPUT13), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT13), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n531_), .A2(new_n537_), .A3(new_n534_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G29gat), .B(G36gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G43gat), .B(G50gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT78), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G1gat), .B(G8gat), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT76), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(G15gat), .ZN(new_n547_));
  INV_X1    g346(.A(G22gat), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G15gat), .A2(G22gat), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G1gat), .A2(G8gat), .ZN(new_n551_));
  AOI22_X1  g350(.A1(new_n549_), .A2(new_n550_), .B1(KEYINPUT14), .B2(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n546_), .B(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n543_), .A2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT79), .ZN(new_n555_));
  INV_X1    g354(.A(new_n553_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n542_), .B(KEYINPUT15), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n555_), .A2(new_n558_), .ZN(new_n559_));
  AND2_X1   g358(.A1(G229gat), .A2(G233gat), .ZN(new_n560_));
  OR2_X1    g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  OR2_X1    g360(.A1(new_n543_), .A2(new_n553_), .ZN(new_n562_));
  AND2_X1   g361(.A1(new_n555_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(new_n560_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n561_), .A2(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G113gat), .B(G141gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G169gat), .B(G197gat), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n566_), .B(new_n567_), .Z(new_n568_));
  NAND2_X1  g367(.A1(new_n565_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n568_), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n564_), .B(new_n570_), .C1(new_n560_), .C2(new_n559_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n569_), .A2(KEYINPUT80), .A3(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT80), .ZN(new_n573_));
  INV_X1    g372(.A(new_n571_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n570_), .B1(new_n561_), .B2(new_n564_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n573_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n572_), .A2(new_n576_), .ZN(new_n577_));
  AND3_X1   g376(.A1(new_n438_), .A2(new_n539_), .A3(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n491_), .A2(new_n557_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n513_), .A2(new_n504_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(new_n542_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G232gat), .A2(G233gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n584_), .A2(KEYINPUT35), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n579_), .A2(new_n581_), .A3(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n586_), .A2(KEYINPUT35), .A3(new_n584_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G190gat), .B(G218gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT74), .ZN(new_n589_));
  XOR2_X1   g388(.A(G134gat), .B(G162gat), .Z(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n592_), .A2(KEYINPUT36), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n584_), .A2(KEYINPUT35), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n579_), .A2(new_n581_), .A3(new_n594_), .A4(new_n585_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n587_), .A2(new_n593_), .A3(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT75), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n587_), .A2(KEYINPUT75), .A3(new_n593_), .A4(new_n595_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n587_), .A2(new_n595_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n591_), .B(KEYINPUT36), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(KEYINPUT37), .B1(new_n600_), .B2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n600_), .A2(KEYINPUT37), .A3(new_n603_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n498_), .B(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(new_n553_), .ZN(new_n610_));
  XOR2_X1   g409(.A(G127gat), .B(G155gat), .Z(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT16), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G183gat), .B(G211gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT17), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n614_), .A2(new_n615_), .ZN(new_n617_));
  NOR3_X1   g416(.A1(new_n610_), .A2(new_n616_), .A3(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n610_), .A2(new_n616_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT77), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n610_), .A2(KEYINPUT77), .A3(new_n616_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n618_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n607_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n578_), .A2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT107), .ZN(new_n627_));
  INV_X1    g426(.A(G1gat), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n627_), .A2(new_n628_), .A3(new_n247_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT38), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  AOI22_X1  g430(.A1(new_n411_), .A2(new_n428_), .B1(new_n432_), .B2(new_n436_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n600_), .A2(new_n603_), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n633_), .B(KEYINPUT108), .Z(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n632_), .A2(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n574_), .A2(new_n575_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n539_), .A2(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n639_), .A2(new_n624_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n636_), .A2(new_n640_), .ZN(new_n641_));
  OAI21_X1  g440(.A(G1gat), .B1(new_n641_), .B2(new_n248_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n629_), .A2(new_n630_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n631_), .A2(new_n642_), .A3(new_n643_), .ZN(G1324gat));
  INV_X1    g443(.A(G8gat), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n627_), .A2(new_n645_), .A3(new_n433_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n641_), .A2(new_n343_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT109), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n645_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT39), .ZN(new_n650_));
  OAI21_X1  g449(.A(KEYINPUT109), .B1(new_n641_), .B2(new_n343_), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n649_), .A2(new_n650_), .A3(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n650_), .B1(new_n649_), .B2(new_n651_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n646_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT40), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n654_), .B(new_n655_), .ZN(G1325gat));
  INV_X1    g455(.A(new_n428_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n627_), .A2(new_n547_), .A3(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(G15gat), .B1(new_n641_), .B2(new_n428_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(KEYINPUT110), .B(KEYINPUT41), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n659_), .A2(new_n660_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n658_), .A2(new_n661_), .A3(new_n662_), .ZN(G1326gat));
  NAND3_X1  g462(.A1(new_n627_), .A2(new_n548_), .A3(new_n392_), .ZN(new_n664_));
  OAI21_X1  g463(.A(G22gat), .B1(new_n641_), .B2(new_n409_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT42), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(G1327gat));
  NOR2_X1   g466(.A1(new_n633_), .A2(new_n623_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n578_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  OR3_X1    g469(.A1(new_n670_), .A2(G29gat), .A3(new_n248_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n639_), .A2(new_n623_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT43), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n673_), .B1(new_n438_), .B2(new_n607_), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n600_), .A2(KEYINPUT37), .A3(new_n603_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n675_), .A2(new_n604_), .ZN(new_n676_));
  NOR3_X1   g475(.A1(new_n632_), .A2(KEYINPUT43), .A3(new_n676_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n672_), .B1(new_n674_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT44), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  OAI211_X1 g479(.A(KEYINPUT44), .B(new_n672_), .C1(new_n674_), .C2(new_n677_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT111), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n682_), .A2(new_n683_), .A3(new_n247_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(G29gat), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n683_), .B1(new_n682_), .B2(new_n247_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n671_), .B1(new_n685_), .B2(new_n686_), .ZN(G1328gat));
  INV_X1    g486(.A(G36gat), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n669_), .A2(new_n688_), .A3(new_n433_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT45), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n680_), .A2(new_n433_), .A3(new_n681_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT112), .ZN(new_n692_));
  AND3_X1   g491(.A1(new_n691_), .A2(new_n692_), .A3(G36gat), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n692_), .B1(new_n691_), .B2(G36gat), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n690_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT46), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  OAI211_X1 g496(.A(new_n690_), .B(KEYINPUT46), .C1(new_n693_), .C2(new_n694_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(G1329gat));
  INV_X1    g498(.A(G43gat), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n700_), .B1(new_n682_), .B2(new_n657_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT47), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n670_), .A2(G43gat), .A3(new_n428_), .ZN(new_n703_));
  OR3_X1    g502(.A1(new_n701_), .A2(new_n702_), .A3(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n702_), .B1(new_n701_), .B2(new_n703_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1330gat));
  AOI21_X1  g505(.A(G50gat), .B1(new_n669_), .B2(new_n392_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n392_), .A2(G50gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n707_), .B1(new_n682_), .B2(new_n708_), .ZN(G1331gat));
  NOR3_X1   g508(.A1(new_n632_), .A2(new_n539_), .A3(new_n638_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(new_n625_), .ZN(new_n711_));
  AOI211_X1 g510(.A(G57gat), .B(new_n248_), .C1(new_n711_), .C2(KEYINPUT113), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n712_), .B1(KEYINPUT113), .B2(new_n711_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n536_), .A2(new_n538_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n623_), .A2(new_n572_), .A3(new_n576_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n636_), .A2(new_n714_), .A3(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(G57gat), .B1(new_n717_), .B2(new_n248_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n713_), .A2(new_n718_), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT114), .Z(G1332gat));
  OAI21_X1  g519(.A(G64gat), .B1(new_n717_), .B2(new_n343_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT48), .ZN(new_n722_));
  OR2_X1    g521(.A1(new_n343_), .A2(G64gat), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n722_), .B1(new_n711_), .B2(new_n723_), .ZN(G1333gat));
  OAI21_X1  g523(.A(G71gat), .B1(new_n717_), .B2(new_n428_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT49), .ZN(new_n726_));
  OR2_X1    g525(.A1(new_n428_), .A2(G71gat), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n726_), .B1(new_n711_), .B2(new_n727_), .ZN(G1334gat));
  OAI21_X1  g527(.A(G78gat), .B1(new_n717_), .B2(new_n409_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(KEYINPUT115), .B(KEYINPUT50), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n729_), .B(new_n730_), .ZN(new_n731_));
  OR2_X1    g530(.A1(new_n409_), .A2(G78gat), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n731_), .B1(new_n711_), .B2(new_n732_), .ZN(G1335gat));
  NAND2_X1  g532(.A1(new_n710_), .A2(new_n668_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(G85gat), .B1(new_n735_), .B2(new_n247_), .ZN(new_n736_));
  OR2_X1    g535(.A1(new_n674_), .A2(new_n677_), .ZN(new_n737_));
  NOR3_X1   g536(.A1(new_n539_), .A2(new_n623_), .A3(new_n638_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n247_), .A2(G85gat), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n741_), .B(KEYINPUT116), .Z(new_n742_));
  AOI21_X1  g541(.A(new_n736_), .B1(new_n740_), .B2(new_n742_), .ZN(G1336gat));
  AOI21_X1  g542(.A(G92gat), .B1(new_n735_), .B2(new_n433_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n433_), .A2(new_n487_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n740_), .B2(new_n745_), .ZN(G1337gat));
  INV_X1    g545(.A(KEYINPUT118), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n747_), .A2(KEYINPUT51), .ZN(new_n748_));
  AND4_X1   g547(.A1(new_n485_), .A2(new_n710_), .A3(new_n657_), .A4(new_n668_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT117), .ZN(new_n750_));
  OAI21_X1  g549(.A(G99gat), .B1(new_n739_), .B2(new_n428_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n748_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT51), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n752_), .B1(KEYINPUT118), .B2(new_n753_), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n750_), .A2(new_n747_), .A3(KEYINPUT51), .A4(new_n751_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n754_), .A2(new_n755_), .ZN(G1338gat));
  XNOR2_X1  g555(.A(KEYINPUT119), .B(KEYINPUT53), .ZN(new_n757_));
  OAI21_X1  g556(.A(G106gat), .B1(new_n739_), .B2(new_n409_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT52), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT52), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n760_), .B(G106gat), .C1(new_n739_), .C2(new_n409_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n392_), .A2(new_n448_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n734_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n757_), .B1(new_n762_), .B2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n757_), .ZN(new_n767_));
  AOI211_X1 g566(.A(new_n764_), .B(new_n767_), .C1(new_n759_), .C2(new_n761_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n766_), .A2(new_n768_), .ZN(G1339gat));
  INV_X1    g568(.A(KEYINPUT120), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n623_), .A2(new_n572_), .A3(new_n576_), .A4(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n715_), .A2(KEYINPUT120), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n539_), .A2(new_n676_), .A3(new_n771_), .A4(new_n772_), .ZN(new_n773_));
  XOR2_X1   g572(.A(new_n773_), .B(KEYINPUT54), .Z(new_n774_));
  OAI21_X1  g573(.A(new_n570_), .B1(new_n563_), .B2(new_n560_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n775_), .B1(new_n560_), .B2(new_n559_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n776_), .A2(new_n575_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n531_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT55), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n517_), .A2(new_n499_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT71), .ZN(new_n781_));
  AOI22_X1  g580(.A1(new_n491_), .A2(new_n500_), .B1(new_n580_), .B2(new_n498_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n781_), .A2(new_n521_), .A3(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n779_), .B1(new_n783_), .B2(new_n524_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n783_), .A2(new_n524_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NOR3_X1   g585(.A1(new_n783_), .A2(new_n779_), .A3(new_n524_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n533_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT56), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n520_), .B1(new_n519_), .B2(new_n521_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n522_), .B1(new_n791_), .B2(new_n779_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n787_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n794_), .A2(KEYINPUT56), .A3(new_n533_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n778_), .B1(new_n790_), .B2(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n607_), .B1(new_n796_), .B2(KEYINPUT58), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT122), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT58), .ZN(new_n800_));
  AOI211_X1 g599(.A(new_n800_), .B(new_n778_), .C1(new_n790_), .C2(new_n795_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  OAI211_X1 g601(.A(KEYINPUT122), .B(new_n607_), .C1(new_n796_), .C2(KEYINPUT58), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n799_), .A2(new_n802_), .A3(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT57), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n535_), .A2(new_n777_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT121), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n532_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n807_), .B1(new_n808_), .B2(KEYINPUT56), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n788_), .A2(KEYINPUT121), .A3(new_n789_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n809_), .A2(new_n810_), .A3(new_n795_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n638_), .A2(new_n531_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n806_), .B1(new_n811_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n633_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n805_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT123), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n633_), .A2(KEYINPUT57), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  AOI211_X1 g618(.A(new_n789_), .B(new_n532_), .C1(new_n792_), .C2(new_n793_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n820_), .B1(new_n807_), .B2(new_n790_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n812_), .B1(new_n821_), .B2(new_n810_), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n817_), .B(new_n819_), .C1(new_n822_), .C2(new_n806_), .ZN(new_n823_));
  OAI21_X1  g622(.A(KEYINPUT123), .B1(new_n814_), .B2(new_n818_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n804_), .A2(new_n816_), .A3(new_n823_), .A4(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n774_), .B1(new_n825_), .B2(new_n624_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n434_), .A2(new_n657_), .A3(new_n247_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(G113gat), .B1(new_n828_), .B2(new_n638_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n827_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n633_), .B1(new_n822_), .B2(new_n806_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n531_), .A2(new_n777_), .ZN(new_n832_));
  AOI21_X1  g631(.A(KEYINPUT56), .B1(new_n794_), .B2(new_n533_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n832_), .B1(new_n833_), .B2(new_n820_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n676_), .B1(new_n834_), .B2(new_n800_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n801_), .B1(new_n835_), .B2(KEYINPUT122), .ZN(new_n836_));
  AOI22_X1  g635(.A1(new_n805_), .A2(new_n831_), .B1(new_n836_), .B2(new_n799_), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n823_), .A2(new_n824_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n623_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  OAI211_X1 g638(.A(KEYINPUT59), .B(new_n830_), .C1(new_n839_), .C2(new_n774_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT59), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n841_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n842_));
  AND3_X1   g641(.A1(new_n840_), .A2(KEYINPUT124), .A3(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(KEYINPUT124), .B1(new_n840_), .B2(new_n842_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n577_), .A2(G113gat), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n829_), .B1(new_n845_), .B2(new_n846_), .ZN(G1340gat));
  AOI21_X1  g646(.A(new_n539_), .B1(new_n840_), .B2(new_n842_), .ZN(new_n848_));
  INV_X1    g647(.A(G120gat), .ZN(new_n849_));
  INV_X1    g648(.A(new_n828_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n849_), .B1(new_n539_), .B2(KEYINPUT60), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n849_), .A2(KEYINPUT60), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n851_), .B1(KEYINPUT125), .B2(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n853_), .B1(KEYINPUT125), .B2(new_n851_), .ZN(new_n854_));
  OAI22_X1  g653(.A1(new_n848_), .A2(new_n849_), .B1(new_n850_), .B2(new_n854_), .ZN(G1341gat));
  AOI21_X1  g654(.A(G127gat), .B1(new_n828_), .B2(new_n623_), .ZN(new_n856_));
  AND2_X1   g655(.A1(new_n623_), .A2(G127gat), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n856_), .B1(new_n845_), .B2(new_n857_), .ZN(G1342gat));
  AOI21_X1  g657(.A(G134gat), .B1(new_n828_), .B2(new_n635_), .ZN(new_n859_));
  AND2_X1   g658(.A1(new_n607_), .A2(G134gat), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n859_), .B1(new_n845_), .B2(new_n860_), .ZN(G1343gat));
  INV_X1    g660(.A(new_n826_), .ZN(new_n862_));
  NOR4_X1   g661(.A1(new_n409_), .A2(new_n657_), .A3(new_n433_), .A4(new_n248_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n864_), .A2(new_n637_), .ZN(new_n865_));
  XOR2_X1   g664(.A(new_n865_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g665(.A1(new_n864_), .A2(new_n539_), .ZN(new_n867_));
  XOR2_X1   g666(.A(new_n867_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g667(.A1(new_n864_), .A2(new_n624_), .ZN(new_n869_));
  XOR2_X1   g668(.A(KEYINPUT61), .B(G155gat), .Z(new_n870_));
  XNOR2_X1  g669(.A(new_n869_), .B(new_n870_), .ZN(G1346gat));
  OAI21_X1  g670(.A(G162gat), .B1(new_n864_), .B2(new_n676_), .ZN(new_n872_));
  OR2_X1    g671(.A1(new_n634_), .A2(G162gat), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n864_), .B2(new_n873_), .ZN(G1347gat));
  INV_X1    g673(.A(G169gat), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n826_), .A2(new_n392_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n430_), .A2(new_n433_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n638_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(KEYINPUT126), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n875_), .B1(new_n876_), .B2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT62), .ZN(new_n882_));
  AND2_X1   g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n881_), .A2(new_n882_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n876_), .A2(new_n878_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n638_), .A2(new_n256_), .ZN(new_n886_));
  OAI22_X1  g685(.A1(new_n883_), .A2(new_n884_), .B1(new_n885_), .B2(new_n886_), .ZN(G1348gat));
  NOR2_X1   g686(.A1(new_n885_), .A2(new_n539_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(new_n257_), .ZN(G1349gat));
  NAND3_X1  g688(.A1(new_n876_), .A2(new_n623_), .A3(new_n878_), .ZN(new_n890_));
  MUX2_X1   g689(.A(new_n279_), .B(G183gat), .S(new_n890_), .Z(G1350gat));
  OAI21_X1  g690(.A(G190gat), .B1(new_n885_), .B2(new_n676_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n635_), .A2(new_n280_), .ZN(new_n893_));
  XOR2_X1   g692(.A(new_n893_), .B(KEYINPUT127), .Z(new_n894_));
  OAI21_X1  g693(.A(new_n892_), .B1(new_n885_), .B2(new_n894_), .ZN(G1351gat));
  NOR4_X1   g694(.A1(new_n409_), .A2(new_n657_), .A3(new_n343_), .A4(new_n247_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n862_), .A2(new_n896_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n897_), .A2(new_n637_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(new_n284_), .ZN(G1352gat));
  NOR2_X1   g698(.A1(new_n897_), .A2(new_n539_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(new_n287_), .ZN(G1353gat));
  NOR2_X1   g700(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n902_));
  AND2_X1   g701(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n903_));
  NOR4_X1   g702(.A1(new_n897_), .A2(new_n624_), .A3(new_n902_), .A4(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n897_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(new_n623_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n904_), .B1(new_n906_), .B2(new_n902_), .ZN(G1354gat));
  OR3_X1    g706(.A1(new_n897_), .A2(G218gat), .A3(new_n634_), .ZN(new_n908_));
  OAI21_X1  g707(.A(G218gat), .B1(new_n897_), .B2(new_n676_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(G1355gat));
endmodule


