//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 0 0 0 1 1 0 0 1 1 0 0 1 1 1 0 1 0 0 0 1 1 0 0 0 0 1 0 1 1 1 1 0 1 1 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n726_, new_n727_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n833_, new_n834_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n842_, new_n843_, new_n844_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n881_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_, new_n900_;
  XNOR2_X1  g000(.A(G1gat), .B(G8gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT71), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT70), .B(G1gat), .ZN(new_n204_));
  INV_X1    g003(.A(G8gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT14), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G15gat), .B(G22gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  OR2_X1    g007(.A1(new_n203_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n203_), .A2(new_n208_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G231gat), .A2(G233gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT72), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n211_), .B(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G57gat), .B(G64gat), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n215_), .A2(KEYINPUT11), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(KEYINPUT11), .ZN(new_n217_));
  XNOR2_X1  g016(.A(G71gat), .B(G78gat), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n216_), .A2(new_n217_), .A3(new_n219_), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n220_), .B1(new_n217_), .B2(new_n219_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n214_), .B(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT74), .ZN(new_n223_));
  XOR2_X1   g022(.A(G183gat), .B(G211gat), .Z(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G127gat), .B(G155gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n226_), .B(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT17), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  XOR2_X1   g029(.A(new_n223_), .B(new_n230_), .Z(new_n231_));
  NOR2_X1   g030(.A1(new_n222_), .A2(KEYINPUT17), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(new_n228_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n231_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(G230gat), .ZN(new_n235_));
  INV_X1    g034(.A(G233gat), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G99gat), .A2(G106gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT6), .ZN(new_n239_));
  OAI21_X1  g038(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n240_));
  OR3_X1    g039(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n239_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  XOR2_X1   g041(.A(G85gat), .B(G92gat), .Z(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT8), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT10), .B(G99gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT64), .B(G106gat), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT65), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G85gat), .A2(G92gat), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n251_), .A2(KEYINPUT9), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n243_), .A2(KEYINPUT9), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n250_), .A2(new_n252_), .A3(new_n239_), .A4(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n245_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(new_n221_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT12), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n221_), .B1(new_n245_), .B2(new_n254_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT12), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n237_), .B1(new_n257_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n237_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n262_), .B1(new_n263_), .B2(new_n256_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G120gat), .B(G148gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(G204gat), .ZN(new_n266_));
  XOR2_X1   g065(.A(KEYINPUT5), .B(G176gat), .Z(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  OR2_X1    g067(.A1(new_n264_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n264_), .A2(new_n268_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT13), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n269_), .A2(KEYINPUT13), .A3(new_n270_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G29gat), .B(G36gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G43gat), .B(G50gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n211_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT76), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT77), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n211_), .A2(new_n278_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G229gat), .A2(G233gat), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n278_), .B(KEYINPUT15), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n287_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n288_), .A2(new_n284_), .A3(new_n279_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n286_), .A2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G113gat), .B(G141gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G169gat), .B(G197gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n290_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n290_), .A2(new_n293_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n275_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT102), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT102), .B1(new_n275_), .B2(new_n297_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT99), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G8gat), .B(G36gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(G92gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT18), .B(G64gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G197gat), .B(G204gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT21), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G211gat), .B(G218gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT21), .B1(new_n309_), .B2(KEYINPUT89), .ZN(new_n313_));
  INV_X1    g112(.A(G204gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(G197gat), .ZN(new_n315_));
  INV_X1    g114(.A(G197gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(G204gat), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n315_), .A2(new_n317_), .A3(KEYINPUT89), .ZN(new_n318_));
  AND2_X1   g117(.A1(G211gat), .A2(G218gat), .ZN(new_n319_));
  NOR2_X1   g118(.A1(G211gat), .A2(G218gat), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n318_), .A2(new_n321_), .ZN(new_n322_));
  NOR3_X1   g121(.A1(new_n313_), .A2(new_n322_), .A3(KEYINPUT90), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT90), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n311_), .B1(KEYINPUT89), .B2(new_n309_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT21), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n315_), .A2(new_n317_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT89), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n326_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n324_), .B1(new_n325_), .B2(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n312_), .B1(new_n323_), .B2(new_n330_), .ZN(new_n331_));
  AND2_X1   g130(.A1(G183gat), .A2(G190gat), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT23), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(KEYINPUT79), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT79), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT23), .ZN(new_n338_));
  AND2_X1   g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G183gat), .A2(G190gat), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n335_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  OR2_X1    g140(.A1(KEYINPUT92), .A2(KEYINPUT24), .ZN(new_n342_));
  NAND2_X1  g141(.A1(KEYINPUT92), .A2(KEYINPUT24), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(G169gat), .ZN(new_n345_));
  INV_X1    g144(.A(G176gat), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n344_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n346_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G169gat), .A2(G176gat), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n342_), .A2(new_n348_), .A3(new_n349_), .A4(new_n343_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(KEYINPUT25), .B(G183gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT26), .B(G190gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND4_X1  g152(.A1(new_n341_), .A2(new_n347_), .A3(new_n350_), .A4(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n349_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT22), .B(G169gat), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n355_), .B1(new_n356_), .B2(new_n346_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n340_), .A2(KEYINPUT23), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n358_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(G183gat), .A2(G190gat), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n357_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n354_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n331_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G226gat), .A2(G233gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT19), .ZN(new_n365_));
  OAI21_X1  g164(.A(KEYINPUT90), .B1(new_n313_), .B2(new_n322_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n325_), .A2(new_n329_), .A3(new_n324_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n336_), .A2(new_n338_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n334_), .B1(new_n369_), .B2(new_n332_), .ZN(new_n370_));
  AND2_X1   g169(.A1(KEYINPUT78), .A2(G190gat), .ZN(new_n371_));
  NOR2_X1   g170(.A1(KEYINPUT78), .A2(G190gat), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n373_), .A2(G183gat), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n357_), .B1(new_n370_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT26), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(G190gat), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n351_), .B(new_n377_), .C1(new_n373_), .C2(new_n376_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n358_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n379_), .B1(new_n369_), .B2(new_n332_), .ZN(new_n380_));
  OR2_X1    g179(.A1(new_n348_), .A2(KEYINPUT24), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n348_), .A2(KEYINPUT24), .A3(new_n349_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n378_), .A2(new_n380_), .A3(new_n381_), .A4(new_n382_), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n368_), .A2(new_n375_), .A3(new_n383_), .A4(new_n312_), .ZN(new_n384_));
  AND4_X1   g183(.A1(KEYINPUT20), .A2(new_n363_), .A3(new_n365_), .A4(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT20), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n375_), .A2(new_n383_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n386_), .B1(new_n331_), .B2(new_n387_), .ZN(new_n388_));
  AOI22_X1  g187(.A1(new_n366_), .A2(new_n367_), .B1(new_n311_), .B2(new_n310_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n389_), .A2(new_n361_), .A3(new_n354_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n365_), .B1(new_n388_), .B2(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n308_), .B1(new_n385_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n365_), .ZN(new_n393_));
  AND2_X1   g192(.A1(new_n375_), .A2(new_n383_), .ZN(new_n394_));
  OAI21_X1  g193(.A(KEYINPUT20), .B1(new_n394_), .B2(new_n389_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n331_), .A2(new_n362_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n393_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n386_), .B1(new_n331_), .B2(new_n362_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n398_), .A2(new_n365_), .A3(new_n384_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n397_), .A2(new_n307_), .A3(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(KEYINPUT27), .B1(new_n392_), .B2(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n307_), .B1(new_n397_), .B2(new_n399_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n363_), .A2(KEYINPUT20), .A3(new_n384_), .A4(new_n393_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT96), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n365_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT96), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n398_), .A2(new_n406_), .A3(new_n393_), .A4(new_n384_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n404_), .A2(new_n405_), .A3(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n402_), .B1(new_n408_), .B2(new_n307_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n401_), .B1(KEYINPUT27), .B2(new_n409_), .ZN(new_n410_));
  OR2_X1    g209(.A1(G127gat), .A2(G134gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G127gat), .A2(G134gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(G113gat), .ZN(new_n414_));
  INV_X1    g213(.A(G120gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G113gat), .A2(G120gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n413_), .A2(new_n418_), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n411_), .A2(new_n416_), .A3(new_n412_), .A4(new_n417_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT86), .ZN(new_n424_));
  INV_X1    g223(.A(G141gat), .ZN(new_n425_));
  INV_X1    g224(.A(G148gat), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n424_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n423_), .B1(new_n427_), .B2(KEYINPUT3), .ZN(new_n428_));
  NAND3_X1  g227(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n428_), .B(new_n429_), .C1(KEYINPUT3), .C2(new_n427_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT84), .ZN(new_n431_));
  INV_X1    g230(.A(G155gat), .ZN(new_n432_));
  INV_X1    g231(.A(G162gat), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n431_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT84), .B1(G155gat), .B2(G162gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G155gat), .A2(G162gat), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(KEYINPUT1), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n436_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT85), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  OR2_X1    g241(.A1(new_n437_), .A2(KEYINPUT1), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n436_), .A2(KEYINPUT85), .A3(new_n439_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n442_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  OR3_X1    g244(.A1(KEYINPUT83), .A2(G141gat), .A3(G148gat), .ZN(new_n446_));
  OAI21_X1  g245(.A(KEYINPUT83), .B1(G141gat), .B2(G148gat), .ZN(new_n447_));
  AOI22_X1  g246(.A1(new_n446_), .A2(new_n447_), .B1(G141gat), .B2(G148gat), .ZN(new_n448_));
  AOI221_X4 g247(.A(new_n422_), .B1(new_n430_), .B2(new_n438_), .C1(new_n445_), .C2(new_n448_), .ZN(new_n449_));
  AND3_X1   g248(.A1(new_n419_), .A2(KEYINPUT80), .A3(new_n420_), .ZN(new_n450_));
  NOR3_X1   g249(.A1(new_n413_), .A2(new_n418_), .A3(KEYINPUT80), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n445_), .A2(new_n448_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n430_), .A2(new_n438_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n452_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(KEYINPUT93), .B1(new_n449_), .B2(new_n455_), .ZN(new_n456_));
  AOI22_X1  g255(.A1(new_n445_), .A2(new_n448_), .B1(new_n430_), .B2(new_n438_), .ZN(new_n457_));
  AOI21_X1  g256(.A(KEYINPUT93), .B1(new_n457_), .B2(new_n421_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n456_), .A2(KEYINPUT4), .A3(new_n459_), .ZN(new_n460_));
  NOR3_X1   g259(.A1(new_n457_), .A2(KEYINPUT4), .A3(new_n452_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G225gat), .A2(G233gat), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n460_), .A2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n453_), .A2(new_n454_), .A3(new_n421_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n465_), .B1(new_n452_), .B2(new_n457_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n458_), .B1(new_n466_), .B2(KEYINPUT93), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(new_n462_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G1gat), .B(G29gat), .ZN(new_n469_));
  INV_X1    g268(.A(G85gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(KEYINPUT0), .B(G57gat), .ZN(new_n472_));
  XOR2_X1   g271(.A(new_n471_), .B(new_n472_), .Z(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n464_), .A2(new_n468_), .A3(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT98), .ZN(new_n476_));
  AOI22_X1  g275(.A1(new_n460_), .A2(new_n463_), .B1(new_n467_), .B2(new_n462_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n476_), .B1(new_n477_), .B2(new_n474_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n462_), .ZN(new_n479_));
  OR2_X1    g278(.A1(new_n457_), .A2(new_n452_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n479_), .B1(new_n480_), .B2(KEYINPUT4), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n481_), .B1(new_n467_), .B2(KEYINPUT4), .ZN(new_n482_));
  AND3_X1   g281(.A1(new_n456_), .A2(new_n462_), .A3(new_n459_), .ZN(new_n483_));
  OAI211_X1 g282(.A(KEYINPUT98), .B(new_n473_), .C1(new_n482_), .C2(new_n483_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n410_), .A2(new_n475_), .A3(new_n478_), .A4(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT29), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n457_), .A2(new_n486_), .ZN(new_n487_));
  XOR2_X1   g286(.A(new_n487_), .B(KEYINPUT91), .Z(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G78gat), .B(G106gat), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n486_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n490_), .B1(new_n491_), .B2(new_n389_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n490_), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n493_), .B(new_n331_), .C1(new_n457_), .C2(new_n486_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT88), .ZN(new_n496_));
  INV_X1    g295(.A(G228gat), .ZN(new_n497_));
  OAI22_X1  g296(.A1(new_n389_), .A2(new_n496_), .B1(new_n497_), .B2(new_n236_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n499_), .ZN(new_n501_));
  OAI221_X1 g300(.A(new_n501_), .B1(new_n497_), .B2(new_n236_), .C1(new_n389_), .C2(new_n496_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n500_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n495_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G22gat), .B(G50gat), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n492_), .A2(new_n500_), .A3(new_n494_), .A4(new_n502_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n504_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n506_), .B1(new_n504_), .B2(new_n507_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n489_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  AND4_X1   g310(.A1(new_n492_), .A2(new_n494_), .A3(new_n500_), .A4(new_n502_), .ZN(new_n512_));
  AOI22_X1  g311(.A1(new_n492_), .A2(new_n494_), .B1(new_n500_), .B2(new_n502_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n505_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n514_), .A2(new_n488_), .A3(new_n508_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n511_), .A2(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n303_), .B1(new_n485_), .B2(new_n516_), .ZN(new_n517_));
  AND3_X1   g316(.A1(new_n514_), .A2(new_n488_), .A3(new_n508_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n488_), .B1(new_n514_), .B2(new_n508_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  AND3_X1   g319(.A1(new_n478_), .A2(new_n484_), .A3(new_n475_), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n520_), .A2(new_n521_), .A3(KEYINPUT99), .A4(new_n410_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n517_), .A2(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n475_), .A2(KEYINPUT33), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT33), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n525_), .B1(new_n477_), .B2(new_n474_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n524_), .A2(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n461_), .A2(new_n479_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n460_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT94), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n474_), .B1(new_n467_), .B2(new_n479_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n460_), .A2(new_n528_), .A3(KEYINPUT94), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n531_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  AND2_X1   g333(.A1(new_n392_), .A2(new_n400_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(KEYINPUT95), .B1(new_n527_), .B2(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n478_), .A2(new_n484_), .A3(new_n475_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n385_), .A2(new_n391_), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n308_), .A2(KEYINPUT32), .ZN(new_n540_));
  OAI21_X1  g339(.A(KEYINPUT97), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n408_), .A2(new_n540_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT97), .ZN(new_n544_));
  OAI211_X1 g343(.A(new_n538_), .B(new_n543_), .C1(new_n544_), .C2(new_n542_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n475_), .A2(KEYINPUT33), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n477_), .A2(new_n525_), .A3(new_n474_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT95), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n548_), .A2(new_n549_), .A3(new_n535_), .A4(new_n534_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n537_), .A2(new_n545_), .A3(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n523_), .B1(new_n516_), .B2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT30), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n387_), .B(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(G43gat), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G227gat), .A2(G233gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(G15gat), .ZN(new_n557_));
  XOR2_X1   g356(.A(G71gat), .B(G99gat), .Z(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n555_), .B(new_n559_), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n452_), .B(KEYINPUT31), .Z(new_n561_));
  NOR2_X1   g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT81), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n560_), .A2(new_n561_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT82), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n563_), .A2(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(KEYINPUT100), .B1(new_n552_), .B2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n410_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n520_), .A2(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n567_), .A2(new_n521_), .A3(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT100), .ZN(new_n572_));
  INV_X1    g371(.A(new_n567_), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n551_), .A2(new_n516_), .ZN(new_n574_));
  OAI211_X1 g373(.A(new_n572_), .B(new_n573_), .C1(new_n574_), .C2(new_n523_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n568_), .A2(new_n571_), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n255_), .A2(new_n287_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(KEYINPUT67), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G232gat), .A2(G233gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT34), .ZN(new_n581_));
  XNOR2_X1  g380(.A(KEYINPUT66), .B(KEYINPUT35), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n579_), .A2(new_n581_), .A3(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n278_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n578_), .B1(new_n584_), .B2(new_n255_), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n583_), .A2(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n581_), .A2(new_n582_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n583_), .B1(new_n585_), .B2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n586_), .A2(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(G190gat), .B(G218gat), .Z(new_n590_));
  XNOR2_X1  g389(.A(G134gat), .B(G162gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(KEYINPUT68), .B(KEYINPUT36), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n594_), .B(KEYINPUT69), .Z(new_n595_));
  NAND2_X1  g394(.A1(new_n589_), .A2(new_n595_), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n592_), .B(KEYINPUT36), .Z(new_n597_));
  NAND3_X1  g396(.A1(new_n586_), .A2(new_n588_), .A3(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n596_), .A2(new_n598_), .ZN(new_n599_));
  NOR3_X1   g398(.A1(new_n577_), .A2(KEYINPUT103), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT103), .ZN(new_n601_));
  INV_X1    g400(.A(new_n599_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n601_), .B1(new_n576_), .B2(new_n602_), .ZN(new_n603_));
  OAI211_X1 g402(.A(new_n234_), .B(new_n302_), .C1(new_n600_), .C2(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(G1gat), .B1(new_n604_), .B2(new_n521_), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n599_), .B(KEYINPUT37), .Z(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n577_), .A2(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n234_), .B(KEYINPUT75), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n608_), .A2(new_n298_), .A3(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n611_), .A2(new_n538_), .A3(new_n204_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(KEYINPUT38), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n613_), .A2(KEYINPUT101), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(KEYINPUT101), .ZN(new_n615_));
  OAI221_X1 g414(.A(new_n605_), .B1(KEYINPUT38), .B2(new_n612_), .C1(new_n614_), .C2(new_n615_), .ZN(G1324gat));
  NAND3_X1  g415(.A1(new_n611_), .A2(new_n205_), .A3(new_n569_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT39), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n604_), .A2(new_n410_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n618_), .B1(new_n619_), .B2(G8gat), .ZN(new_n620_));
  OAI211_X1 g419(.A(new_n618_), .B(G8gat), .C1(new_n604_), .C2(new_n410_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n617_), .B1(new_n620_), .B2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT40), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  OAI211_X1 g424(.A(KEYINPUT40), .B(new_n617_), .C1(new_n620_), .C2(new_n622_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(G1325gat));
  NOR3_X1   g426(.A1(new_n610_), .A2(G15gat), .A3(new_n573_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT104), .ZN(new_n629_));
  OAI21_X1  g428(.A(G15gat), .B1(new_n604_), .B2(new_n573_), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n630_), .A2(KEYINPUT41), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(KEYINPUT41), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n629_), .A2(new_n631_), .A3(new_n632_), .ZN(G1326gat));
  OR3_X1    g432(.A1(new_n610_), .A2(G22gat), .A3(new_n516_), .ZN(new_n634_));
  OAI21_X1  g433(.A(G22gat), .B1(new_n604_), .B2(new_n516_), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n635_), .A2(KEYINPUT42), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n635_), .A2(KEYINPUT42), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n634_), .B1(new_n637_), .B2(new_n638_), .ZN(G1327gat));
  AOI21_X1  g438(.A(new_n609_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT43), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n576_), .A2(new_n641_), .A3(new_n607_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n641_), .B1(new_n576_), .B2(new_n607_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n640_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT44), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  OAI211_X1 g445(.A(new_n640_), .B(KEYINPUT44), .C1(new_n642_), .C2(new_n643_), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n646_), .A2(G29gat), .A3(new_n538_), .A4(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(G29gat), .ZN(new_n649_));
  INV_X1    g448(.A(new_n609_), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n576_), .A2(new_n298_), .A3(new_n650_), .A4(new_n599_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n649_), .B1(new_n651_), .B2(new_n521_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n648_), .A2(new_n652_), .ZN(G1328gat));
  INV_X1    g452(.A(KEYINPUT45), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n410_), .B(KEYINPUT106), .Z(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n651_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(G36gat), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n654_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  NOR4_X1   g458(.A1(new_n651_), .A2(KEYINPUT45), .A3(G36gat), .A4(new_n656_), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n659_), .A2(KEYINPUT107), .A3(new_n660_), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n646_), .A2(KEYINPUT105), .A3(new_n569_), .A4(new_n647_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT107), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n646_), .A2(new_n569_), .A3(new_n647_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT105), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n658_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  AOI211_X1 g466(.A(KEYINPUT46), .B(new_n661_), .C1(new_n664_), .C2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT46), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n665_), .A2(new_n666_), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n670_), .A2(new_n663_), .A3(G36gat), .A4(new_n662_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n661_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n669_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n668_), .A2(new_n673_), .ZN(G1329gat));
  NAND4_X1  g473(.A1(new_n646_), .A2(G43gat), .A3(new_n567_), .A4(new_n647_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n651_), .A2(new_n573_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n675_), .B1(G43gat), .B2(new_n676_), .ZN(new_n677_));
  XOR2_X1   g476(.A(KEYINPUT108), .B(KEYINPUT47), .Z(new_n678_));
  XNOR2_X1  g477(.A(new_n677_), .B(new_n678_), .ZN(G1330gat));
  OR3_X1    g478(.A1(new_n651_), .A2(G50gat), .A3(new_n516_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n646_), .A2(new_n520_), .A3(new_n647_), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n681_), .A2(KEYINPUT109), .A3(G50gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(KEYINPUT109), .B1(new_n681_), .B2(G50gat), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n680_), .B1(new_n682_), .B2(new_n683_), .ZN(G1331gat));
  NAND2_X1  g483(.A1(new_n275_), .A2(new_n297_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n685_), .A2(new_n650_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n608_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(G57gat), .B1(new_n688_), .B2(new_n538_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n600_), .A2(new_n603_), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n690_), .A2(new_n650_), .A3(new_n685_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n538_), .A2(G57gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n689_), .B1(new_n691_), .B2(new_n692_), .ZN(G1332gat));
  INV_X1    g492(.A(G64gat), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n688_), .A2(new_n694_), .A3(new_n655_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT48), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n691_), .A2(new_n655_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n696_), .B1(new_n697_), .B2(G64gat), .ZN(new_n698_));
  AOI211_X1 g497(.A(KEYINPUT48), .B(new_n694_), .C1(new_n691_), .C2(new_n655_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n695_), .B1(new_n698_), .B2(new_n699_), .ZN(G1333gat));
  INV_X1    g499(.A(KEYINPUT49), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n691_), .A2(new_n567_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n701_), .B1(new_n702_), .B2(G71gat), .ZN(new_n703_));
  INV_X1    g502(.A(G71gat), .ZN(new_n704_));
  AOI211_X1 g503(.A(KEYINPUT49), .B(new_n704_), .C1(new_n691_), .C2(new_n567_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n567_), .A2(new_n704_), .ZN(new_n706_));
  XOR2_X1   g505(.A(new_n706_), .B(KEYINPUT110), .Z(new_n707_));
  OAI22_X1  g506(.A1(new_n703_), .A2(new_n705_), .B1(new_n687_), .B2(new_n707_), .ZN(G1334gat));
  OR3_X1    g507(.A1(new_n687_), .A2(G78gat), .A3(new_n516_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n691_), .A2(new_n520_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT50), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n710_), .A2(new_n711_), .A3(G78gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n711_), .B1(new_n710_), .B2(G78gat), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n709_), .B1(new_n712_), .B2(new_n713_), .ZN(G1335gat));
  NOR2_X1   g513(.A1(new_n577_), .A2(new_n602_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n685_), .A2(new_n609_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(G85gat), .B1(new_n718_), .B2(new_n538_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT111), .ZN(new_n720_));
  OR3_X1    g519(.A1(new_n642_), .A2(new_n643_), .A3(new_n720_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n720_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n721_), .A2(new_n716_), .A3(new_n722_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n521_), .A2(new_n470_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n719_), .B1(new_n723_), .B2(new_n724_), .ZN(G1336gat));
  AOI21_X1  g524(.A(G92gat), .B1(new_n718_), .B2(new_n569_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n655_), .A2(G92gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n723_), .B2(new_n727_), .ZN(G1337gat));
  NAND3_X1  g527(.A1(new_n721_), .A2(new_n716_), .A3(new_n722_), .ZN(new_n729_));
  OAI21_X1  g528(.A(G99gat), .B1(new_n729_), .B2(new_n573_), .ZN(new_n730_));
  OR2_X1    g529(.A1(new_n573_), .A2(new_n246_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n730_), .B1(new_n717_), .B2(new_n731_), .ZN(new_n732_));
  XOR2_X1   g531(.A(KEYINPUT112), .B(KEYINPUT51), .Z(new_n733_));
  XNOR2_X1  g532(.A(new_n732_), .B(new_n733_), .ZN(G1338gat));
  OAI211_X1 g533(.A(new_n520_), .B(new_n716_), .C1(new_n642_), .C2(new_n643_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT52), .ZN(new_n736_));
  OAI211_X1 g535(.A(new_n735_), .B(G106gat), .C1(KEYINPUT113), .C2(new_n736_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n736_), .A2(KEYINPUT113), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  OR3_X1    g538(.A1(new_n717_), .A2(new_n247_), .A3(new_n516_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n737_), .A2(new_n738_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n739_), .A2(new_n740_), .A3(new_n741_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g542(.A1(new_n609_), .A2(new_n297_), .ZN(new_n744_));
  OR2_X1    g543(.A1(new_n744_), .A2(KEYINPUT114), .ZN(new_n745_));
  INV_X1    g544(.A(new_n275_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n607_), .B1(new_n744_), .B2(KEYINPUT114), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n745_), .A2(new_n746_), .A3(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(KEYINPUT54), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT54), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n745_), .A2(new_n747_), .A3(new_n750_), .A4(new_n746_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n749_), .A2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT116), .ZN(new_n754_));
  XNOR2_X1  g553(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n755_));
  OR3_X1    g554(.A1(new_n261_), .A2(new_n754_), .A3(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n257_), .A2(new_n237_), .A3(new_n260_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n754_), .B1(new_n261_), .B2(new_n755_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n261_), .A2(KEYINPUT55), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n756_), .A2(new_n757_), .A3(new_n758_), .A4(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(new_n268_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT56), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n760_), .A2(KEYINPUT56), .A3(new_n268_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n763_), .A2(KEYINPUT118), .A3(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT118), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n761_), .A2(new_n766_), .A3(new_n762_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n765_), .A2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n283_), .A2(new_n284_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n288_), .A2(new_n285_), .A3(new_n279_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n769_), .A2(new_n293_), .A3(new_n770_), .ZN(new_n771_));
  AND3_X1   g570(.A1(new_n294_), .A2(new_n269_), .A3(new_n771_), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n768_), .A2(KEYINPUT119), .A3(KEYINPUT58), .A4(new_n772_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n765_), .A2(new_n772_), .A3(KEYINPUT58), .A4(new_n767_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT119), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n606_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n765_), .A2(new_n772_), .A3(new_n767_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT58), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n773_), .A2(new_n776_), .A3(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT120), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n271_), .A2(new_n294_), .A3(new_n771_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT117), .B1(new_n760_), .B2(new_n268_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT56), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(new_n296_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n269_), .B1(new_n783_), .B2(KEYINPUT56), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n782_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n787_), .A2(KEYINPUT57), .A3(new_n602_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(KEYINPUT57), .B1(new_n787_), .B2(new_n602_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT120), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n773_), .A2(new_n776_), .A3(new_n792_), .A4(new_n779_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n781_), .A2(new_n791_), .A3(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n234_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n753_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n567_), .A2(new_n570_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n797_), .A2(new_n521_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(KEYINPUT59), .B1(new_n796_), .B2(new_n799_), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n773_), .A2(new_n776_), .A3(new_n779_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n787_), .A2(new_n602_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT57), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n788_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n650_), .B1(new_n801_), .B2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n752_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT59), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n799_), .B1(KEYINPUT121), .B2(new_n808_), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n807_), .B(new_n809_), .C1(KEYINPUT121), .C2(new_n808_), .ZN(new_n810_));
  OAI21_X1  g609(.A(KEYINPUT122), .B1(new_n297_), .B2(new_n414_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n800_), .A2(new_n810_), .A3(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n794_), .A2(new_n795_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n752_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n798_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n815_), .A2(new_n297_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n812_), .A2(new_n816_), .ZN(new_n817_));
  AND3_X1   g616(.A1(new_n800_), .A2(new_n810_), .A3(new_n811_), .ZN(new_n818_));
  AOI22_X1  g617(.A1(new_n817_), .A2(new_n414_), .B1(new_n818_), .B2(KEYINPUT122), .ZN(G1340gat));
  INV_X1    g618(.A(new_n815_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n415_), .B1(new_n746_), .B2(KEYINPUT60), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n415_), .A2(KEYINPUT60), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n821_), .B1(KEYINPUT123), .B2(new_n822_), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n820_), .B(new_n823_), .C1(KEYINPUT123), .C2(new_n821_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n800_), .A2(new_n275_), .A3(new_n810_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(G120gat), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n826_), .ZN(G1341gat));
  AOI21_X1  g626(.A(G127gat), .B1(new_n820_), .B2(new_n609_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n800_), .A2(new_n810_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n234_), .A2(G127gat), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n830_), .B(KEYINPUT124), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n828_), .B1(new_n829_), .B2(new_n831_), .ZN(G1342gat));
  AOI21_X1  g631(.A(G134gat), .B1(new_n820_), .B2(new_n599_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n607_), .A2(G134gat), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n833_), .B1(new_n829_), .B2(new_n834_), .ZN(G1343gat));
  NOR3_X1   g634(.A1(new_n567_), .A2(new_n521_), .A3(new_n516_), .ZN(new_n836_));
  AND3_X1   g635(.A1(new_n814_), .A2(new_n656_), .A3(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n296_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(G141gat), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n837_), .A2(new_n425_), .A3(new_n296_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(G1344gat));
  NAND2_X1  g640(.A1(new_n837_), .A2(new_n275_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(G148gat), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n837_), .A2(new_n426_), .A3(new_n275_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(G1345gat));
  NAND4_X1  g644(.A1(new_n814_), .A2(new_n609_), .A3(new_n656_), .A4(new_n836_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(KEYINPUT61), .B(G155gat), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n846_), .B(new_n847_), .ZN(G1346gat));
  NAND2_X1  g647(.A1(new_n837_), .A2(new_n599_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n606_), .A2(new_n433_), .ZN(new_n850_));
  AOI22_X1  g649(.A1(new_n849_), .A2(new_n433_), .B1(new_n837_), .B2(new_n850_), .ZN(G1347gat));
  INV_X1    g650(.A(KEYINPUT62), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT125), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n656_), .A2(new_n538_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n567_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n609_), .B1(new_n791_), .B2(new_n780_), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n516_), .B(new_n856_), .C1(new_n857_), .C2(new_n753_), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n853_), .B(G169gat), .C1(new_n858_), .C2(new_n297_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n807_), .A2(new_n296_), .A3(new_n516_), .A4(new_n856_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n853_), .B1(new_n861_), .B2(G169gat), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n852_), .B1(new_n860_), .B2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n861_), .A2(G169gat), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(KEYINPUT125), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n865_), .A2(KEYINPUT62), .A3(new_n859_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n858_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n867_), .A2(new_n296_), .A3(new_n356_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n863_), .A2(new_n866_), .A3(new_n868_), .ZN(G1348gat));
  OAI21_X1  g668(.A(new_n346_), .B1(new_n858_), .B2(new_n746_), .ZN(new_n870_));
  OR2_X1    g669(.A1(new_n870_), .A2(KEYINPUT126), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(KEYINPUT126), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n796_), .A2(new_n520_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n746_), .A2(new_n855_), .A3(new_n346_), .ZN(new_n874_));
  AOI22_X1  g673(.A1(new_n871_), .A2(new_n872_), .B1(new_n873_), .B2(new_n874_), .ZN(G1349gat));
  NOR3_X1   g674(.A1(new_n858_), .A2(new_n795_), .A3(new_n351_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n873_), .A2(new_n609_), .A3(new_n856_), .ZN(new_n877_));
  INV_X1    g676(.A(G183gat), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n876_), .B1(new_n877_), .B2(new_n878_), .ZN(G1350gat));
  OAI21_X1  g678(.A(G190gat), .B1(new_n858_), .B2(new_n606_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n599_), .A2(new_n352_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n858_), .B2(new_n881_), .ZN(G1351gat));
  NOR2_X1   g681(.A1(new_n567_), .A2(new_n516_), .ZN(new_n883_));
  AND3_X1   g682(.A1(new_n814_), .A2(new_n883_), .A3(new_n854_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n296_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(G197gat), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n884_), .A2(new_n316_), .A3(new_n296_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(G1352gat));
  NAND4_X1  g687(.A1(new_n814_), .A2(new_n275_), .A3(new_n883_), .A4(new_n854_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g689(.A(KEYINPUT63), .ZN(new_n891_));
  INV_X1    g690(.A(G211gat), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n234_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(KEYINPUT127), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n814_), .A2(new_n883_), .A3(new_n854_), .A4(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n891_), .A2(new_n892_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n895_), .B(new_n896_), .ZN(G1354gat));
  NAND2_X1  g696(.A1(new_n884_), .A2(new_n599_), .ZN(new_n898_));
  INV_X1    g697(.A(G218gat), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n606_), .A2(new_n899_), .ZN(new_n900_));
  AOI22_X1  g699(.A1(new_n898_), .A2(new_n899_), .B1(new_n884_), .B2(new_n900_), .ZN(G1355gat));
endmodule


