//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 0 1 0 0 1 1 1 1 0 1 0 0 0 0 1 0 0 1 1 0 1 0 0 1 1 1 1 1 0 1 1 1 1 1 1 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n612_,
    new_n613_, new_n614_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n653_, new_n654_, new_n655_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n676_, new_n677_, new_n678_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n694_,
    new_n695_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n792_, new_n793_, new_n795_, new_n796_,
    new_n797_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n805_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n813_, new_n814_, new_n815_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n861_, new_n862_, new_n863_, new_n864_,
    new_n865_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n885_;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G169gat), .B(G197gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT15), .ZN(new_n206_));
  INV_X1    g005(.A(G36gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(G29gat), .ZN(new_n208_));
  INV_X1    g007(.A(G29gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G36gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT68), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n208_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n211_), .B1(new_n208_), .B2(new_n210_), .ZN(new_n214_));
  XOR2_X1   g013(.A(G43gat), .B(G50gat), .Z(new_n215_));
  NOR3_X1   g014(.A1(new_n213_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(G43gat), .B(G50gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n209_), .A2(G36gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n207_), .A2(G29gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT68), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n217_), .B1(new_n220_), .B2(new_n212_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n206_), .B1(new_n216_), .B2(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n215_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n220_), .A2(new_n212_), .A3(new_n217_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n223_), .A2(new_n224_), .A3(KEYINPUT15), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n222_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G15gat), .B(G22gat), .ZN(new_n227_));
  INV_X1    g026(.A(G1gat), .ZN(new_n228_));
  INV_X1    g027(.A(G8gat), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT14), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n227_), .A2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G1gat), .B(G8gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n231_), .B(new_n232_), .ZN(new_n233_));
  AND2_X1   g032(.A1(new_n226_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n223_), .A2(new_n224_), .ZN(new_n235_));
  OR2_X1    g034(.A1(new_n235_), .A2(new_n233_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G229gat), .A2(G233gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n234_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n235_), .A2(new_n233_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n237_), .B1(new_n236_), .B2(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n205_), .B1(new_n239_), .B2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n241_), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n243_), .B(new_n204_), .C1(new_n234_), .C2(new_n238_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G183gat), .A2(G190gat), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n246_), .A2(KEYINPUT23), .ZN(new_n247_));
  XOR2_X1   g046(.A(KEYINPUT77), .B(KEYINPUT23), .Z(new_n248_));
  AOI21_X1  g047(.A(new_n247_), .B1(new_n248_), .B2(new_n246_), .ZN(new_n249_));
  OR2_X1    g048(.A1(G169gat), .A2(G176gat), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n250_), .A2(KEYINPUT24), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n249_), .A2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT26), .B(G190gat), .ZN(new_n253_));
  INV_X1    g052(.A(G183gat), .ZN(new_n254_));
  OAI21_X1  g053(.A(KEYINPUT25), .B1(new_n254_), .B2(KEYINPUT75), .ZN(new_n255_));
  OR2_X1    g054(.A1(new_n254_), .A2(KEYINPUT25), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n253_), .B(new_n255_), .C1(new_n256_), .C2(KEYINPUT75), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G169gat), .A2(G176gat), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n250_), .A2(KEYINPUT24), .A3(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT76), .ZN(new_n260_));
  OR2_X1    g059(.A1(new_n259_), .A2(KEYINPUT76), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n252_), .A2(new_n257_), .A3(new_n260_), .A4(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n246_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n263_), .A2(KEYINPUT23), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n264_), .B1(new_n248_), .B2(new_n263_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n265_), .B1(G183gat), .B2(G190gat), .ZN(new_n266_));
  NOR2_X1   g065(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(G169gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n266_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n262_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G227gat), .A2(G233gat), .ZN(new_n271_));
  INV_X1    g070(.A(G71gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(G99gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n270_), .B(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G15gat), .B(G43gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT78), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT30), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n275_), .B(new_n278_), .ZN(new_n279_));
  XOR2_X1   g078(.A(G127gat), .B(G134gat), .Z(new_n280_));
  XNOR2_X1  g079(.A(G113gat), .B(G120gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(new_n282_), .B(KEYINPUT31), .Z(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  OR2_X1    g083(.A1(new_n279_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(KEYINPUT79), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n279_), .A2(new_n284_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT80), .ZN(new_n288_));
  OR2_X1    g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G225gat), .A2(G233gat), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT4), .ZN(new_n292_));
  NOR2_X1   g091(.A1(G141gat), .A2(G148gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT3), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G141gat), .A2(G148gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT2), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G155gat), .A2(G162gat), .ZN(new_n298_));
  NOR2_X1   g097(.A1(G155gat), .A2(G162gat), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n297_), .A2(new_n298_), .A3(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n299_), .B1(KEYINPUT1), .B2(new_n298_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n302_), .B1(KEYINPUT1), .B2(new_n298_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n293_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n303_), .A2(new_n304_), .A3(new_n295_), .ZN(new_n305_));
  AND2_X1   g104(.A1(new_n301_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT81), .ZN(new_n307_));
  OR2_X1    g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n307_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n308_), .A2(new_n309_), .A3(new_n282_), .ZN(new_n310_));
  OR2_X1    g109(.A1(new_n282_), .A2(KEYINPUT92), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n282_), .A2(KEYINPUT92), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n306_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n292_), .B1(new_n310_), .B2(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n306_), .B(KEYINPUT81), .ZN(new_n315_));
  AOI21_X1  g114(.A(KEYINPUT4), .B1(new_n315_), .B2(new_n282_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n291_), .B1(new_n314_), .B2(new_n316_), .ZN(new_n317_));
  AND2_X1   g116(.A1(new_n310_), .A2(new_n313_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(new_n290_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  XOR2_X1   g119(.A(G1gat), .B(G29gat), .Z(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT93), .B(G85gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(KEYINPUT0), .B(G57gat), .ZN(new_n324_));
  XOR2_X1   g123(.A(new_n323_), .B(new_n324_), .Z(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n320_), .A2(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n317_), .A2(new_n319_), .A3(new_n325_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n251_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n265_), .A2(new_n330_), .ZN(new_n331_));
  OR2_X1    g130(.A1(new_n331_), .A2(KEYINPUT89), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT25), .B(G183gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n253_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(new_n259_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT88), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n331_), .A2(KEYINPUT89), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n332_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(G183gat), .A2(G190gat), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n268_), .B1(new_n249_), .B2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G211gat), .B(G218gat), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n341_), .A2(KEYINPUT84), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT21), .ZN(new_n343_));
  XOR2_X1   g142(.A(G197gat), .B(G204gat), .Z(new_n344_));
  OR3_X1    g143(.A1(new_n342_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n342_), .A2(new_n343_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n344_), .B1(KEYINPUT21), .B2(new_n341_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n345_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n338_), .A2(new_n340_), .A3(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT90), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT20), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n353_), .B1(new_n270_), .B2(new_n348_), .ZN(new_n354_));
  AND2_X1   g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  OR2_X1    g154(.A1(new_n350_), .A2(new_n351_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G226gat), .A2(G233gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT19), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n357_), .A2(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n349_), .B1(new_n338_), .B2(new_n340_), .ZN(new_n362_));
  OAI21_X1  g161(.A(KEYINPUT20), .B1(new_n270_), .B2(new_n348_), .ZN(new_n363_));
  NOR3_X1   g162(.A1(new_n362_), .A2(new_n363_), .A3(new_n360_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n361_), .A2(new_n365_), .ZN(new_n366_));
  XOR2_X1   g165(.A(G8gat), .B(G36gat), .Z(new_n367_));
  XNOR2_X1  g166(.A(G64gat), .B(G92gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  AND2_X1   g170(.A1(new_n371_), .A2(KEYINPUT32), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT95), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n366_), .A2(new_n373_), .ZN(new_n374_));
  OR3_X1    g173(.A1(new_n362_), .A2(new_n363_), .A3(new_n359_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT96), .ZN(new_n376_));
  OR4_X1    g175(.A1(KEYINPUT96), .A2(new_n362_), .A3(new_n363_), .A4(new_n359_), .ZN(new_n377_));
  AND2_X1   g176(.A1(new_n350_), .A2(new_n354_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n376_), .B(new_n377_), .C1(new_n360_), .C2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(new_n372_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n329_), .A2(new_n374_), .A3(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT94), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT33), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n328_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n382_), .B1(new_n328_), .B2(new_n383_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n371_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n361_), .A2(new_n387_), .A3(new_n365_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n359_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n371_), .B1(new_n389_), .B2(new_n364_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n325_), .B1(new_n318_), .B2(new_n291_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n290_), .B1(new_n314_), .B2(new_n316_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n317_), .A2(KEYINPUT33), .A3(new_n319_), .A4(new_n325_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n388_), .A2(new_n390_), .A3(new_n393_), .A4(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n381_), .B1(new_n386_), .B2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT86), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT29), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n348_), .B1(new_n306_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(G228gat), .ZN(new_n400_));
  INV_X1    g199(.A(G233gat), .ZN(new_n401_));
  OR2_X1    g200(.A1(new_n401_), .A2(KEYINPUT83), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(KEYINPUT83), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n400_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n399_), .A2(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n306_), .B(new_n307_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n406_), .A2(new_n398_), .ZN(new_n407_));
  OR2_X1    g206(.A1(new_n349_), .A2(new_n404_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n405_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  XOR2_X1   g208(.A(G78gat), .B(G106gat), .Z(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(KEYINPUT85), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n397_), .B1(new_n409_), .B2(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n412_), .B1(new_n411_), .B2(new_n409_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n409_), .A2(new_n397_), .A3(new_n411_), .ZN(new_n414_));
  XOR2_X1   g213(.A(KEYINPUT82), .B(KEYINPUT28), .Z(new_n415_));
  OR3_X1    g214(.A1(new_n315_), .A2(KEYINPUT29), .A3(new_n415_), .ZN(new_n416_));
  XOR2_X1   g215(.A(G22gat), .B(G50gat), .Z(new_n417_));
  OAI21_X1  g216(.A(new_n415_), .B1(new_n315_), .B2(KEYINPUT29), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n416_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n417_), .B1(new_n416_), .B2(new_n418_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n413_), .A2(new_n414_), .A3(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT87), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n411_), .A2(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n409_), .B(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n425_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n422_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n396_), .A2(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n329_), .B1(new_n422_), .B2(new_n426_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT27), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n430_), .B1(new_n366_), .B2(new_n371_), .ZN(new_n431_));
  AND3_X1   g230(.A1(new_n379_), .A2(KEYINPUT97), .A3(new_n387_), .ZN(new_n432_));
  AOI21_X1  g231(.A(KEYINPUT97), .B1(new_n379_), .B2(new_n387_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n431_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n388_), .A2(new_n390_), .ZN(new_n435_));
  AOI21_X1  g234(.A(KEYINPUT98), .B1(new_n435_), .B2(new_n430_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT98), .ZN(new_n437_));
  AOI211_X1 g236(.A(new_n437_), .B(KEYINPUT27), .C1(new_n388_), .C2(new_n390_), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n429_), .B(new_n434_), .C1(new_n436_), .C2(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n289_), .B1(new_n428_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n329_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n289_), .A2(new_n441_), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n427_), .B(new_n434_), .C1(new_n436_), .C2(new_n438_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n245_), .B1(new_n440_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT99), .ZN(new_n447_));
  XOR2_X1   g246(.A(G190gat), .B(G218gat), .Z(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(KEYINPUT69), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G134gat), .B(G162gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n449_), .B(new_n450_), .ZN(new_n451_));
  XOR2_X1   g250(.A(new_n451_), .B(KEYINPUT36), .Z(new_n452_));
  NAND2_X1  g251(.A1(G99gat), .A2(G106gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT6), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT6), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n455_), .A2(G99gat), .A3(G106gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n454_), .A2(new_n456_), .ZN(new_n457_));
  OR2_X1    g256(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n458_));
  INV_X1    g257(.A(G106gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n458_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(G85gat), .ZN(new_n462_));
  INV_X1    g261(.A(G92gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G85gat), .A2(G92gat), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n464_), .A2(KEYINPUT9), .A3(new_n465_), .ZN(new_n466_));
  OR2_X1    g265(.A1(new_n465_), .A2(KEYINPUT9), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n457_), .A2(new_n461_), .A3(new_n466_), .A4(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT65), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n464_), .A2(new_n469_), .A3(new_n465_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT7), .ZN(new_n471_));
  INV_X1    g270(.A(G99gat), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n471_), .A2(new_n472_), .A3(new_n459_), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  AOI211_X1 g274(.A(KEYINPUT8), .B(new_n470_), .C1(new_n475_), .C2(new_n457_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT8), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n457_), .A2(new_n474_), .A3(new_n473_), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n464_), .A2(new_n469_), .A3(new_n465_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n477_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  OAI211_X1 g279(.A(new_n235_), .B(new_n468_), .C1(new_n476_), .C2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n468_), .ZN(new_n482_));
  AND2_X1   g281(.A1(new_n454_), .A2(new_n456_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n473_), .A2(new_n474_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n479_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT8), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n478_), .A2(new_n477_), .A3(new_n479_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n482_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n481_), .B1(new_n226_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT71), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G232gat), .A2(G233gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT34), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n492_), .A2(KEYINPUT35), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n492_), .A2(KEYINPUT35), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n489_), .A2(new_n490_), .A3(new_n495_), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n481_), .B(new_n493_), .C1(new_n226_), .C2(new_n488_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n490_), .B1(new_n489_), .B2(new_n495_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n452_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n499_), .ZN(new_n501_));
  XOR2_X1   g300(.A(KEYINPUT70), .B(KEYINPUT36), .Z(new_n502_));
  NOR2_X1   g301(.A1(new_n451_), .A2(new_n502_), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n501_), .A2(new_n497_), .A3(new_n496_), .A4(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n500_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n500_), .A2(KEYINPUT72), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n505_), .A2(new_n506_), .A3(KEYINPUT37), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT37), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n500_), .B(new_n504_), .C1(KEYINPUT72), .C2(new_n508_), .ZN(new_n509_));
  AND2_X1   g308(.A1(new_n507_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(KEYINPUT73), .A2(KEYINPUT17), .ZN(new_n511_));
  XOR2_X1   g310(.A(G127gat), .B(G155gat), .Z(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT16), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G183gat), .B(G211gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  MUX2_X1   g314(.A(new_n511_), .B(KEYINPUT17), .S(new_n515_), .Z(new_n516_));
  NAND2_X1  g315(.A1(G231gat), .A2(G233gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n233_), .B(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n272_), .A2(G78gat), .ZN(new_n519_));
  INV_X1    g318(.A(G78gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(G71gat), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G57gat), .B(G64gat), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n522_), .B1(new_n523_), .B2(KEYINPUT11), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT66), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n525_), .B1(new_n523_), .B2(KEYINPUT11), .ZN(new_n526_));
  INV_X1    g325(.A(G64gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(G57gat), .ZN(new_n528_));
  INV_X1    g327(.A(G57gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(G64gat), .ZN(new_n530_));
  AND4_X1   g329(.A1(new_n525_), .A2(new_n528_), .A3(new_n530_), .A4(KEYINPUT11), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n524_), .B1(new_n526_), .B2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n528_), .A2(new_n530_), .A3(KEYINPUT11), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT66), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n528_), .A2(new_n530_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT11), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n528_), .A2(new_n530_), .A3(new_n525_), .A4(KEYINPUT11), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n534_), .A2(new_n537_), .A3(new_n522_), .A4(new_n538_), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n532_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n518_), .B(new_n540_), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n516_), .A2(new_n541_), .ZN(new_n542_));
  NOR3_X1   g341(.A1(new_n541_), .A2(new_n515_), .A3(new_n511_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n510_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G230gat), .A2(G233gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(KEYINPUT64), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n548_), .B1(new_n488_), .B2(new_n540_), .ZN(new_n549_));
  NOR3_X1   g348(.A1(new_n488_), .A2(new_n540_), .A3(KEYINPUT12), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT12), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n468_), .B1(new_n476_), .B2(new_n480_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n532_), .A2(new_n539_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n551_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n549_), .B1(new_n550_), .B2(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n488_), .A2(new_n540_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n552_), .A2(new_n553_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n548_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n555_), .A2(new_n558_), .ZN(new_n559_));
  XOR2_X1   g358(.A(G120gat), .B(G148gat), .Z(new_n560_));
  XNOR2_X1  g359(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G176gat), .B(G204gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n559_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n559_), .A2(new_n565_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT13), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n566_), .A2(KEYINPUT13), .A3(new_n567_), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n546_), .A2(new_n572_), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n573_), .B(KEYINPUT74), .Z(new_n574_));
  NAND3_X1  g373(.A1(new_n446_), .A2(new_n447_), .A3(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n574_), .ZN(new_n576_));
  OAI21_X1  g375(.A(KEYINPUT99), .B1(new_n445_), .B2(new_n576_), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n575_), .A2(new_n577_), .A3(new_n228_), .A4(new_n329_), .ZN(new_n578_));
  XOR2_X1   g377(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n578_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n578_), .A2(new_n580_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n572_), .A2(new_n245_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n583_), .A2(new_n545_), .ZN(new_n584_));
  OAI211_X1 g383(.A(new_n505_), .B(new_n584_), .C1(new_n440_), .C2(new_n444_), .ZN(new_n585_));
  OAI21_X1  g384(.A(G1gat), .B1(new_n585_), .B2(new_n441_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n581_), .A2(new_n582_), .A3(new_n586_), .ZN(G1324gat));
  OAI21_X1  g386(.A(new_n434_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n575_), .A2(new_n577_), .A3(new_n229_), .A4(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT39), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n440_), .A2(new_n444_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n592_), .A2(new_n588_), .A3(new_n505_), .A4(new_n584_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n590_), .B1(new_n593_), .B2(G8gat), .ZN(new_n594_));
  INV_X1    g393(.A(new_n588_), .ZN(new_n595_));
  OAI211_X1 g394(.A(new_n590_), .B(G8gat), .C1(new_n585_), .C2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n589_), .B1(new_n594_), .B2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(KEYINPUT40), .ZN(new_n599_));
  XNOR2_X1  g398(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT40), .ZN(new_n601_));
  OAI211_X1 g400(.A(new_n589_), .B(new_n601_), .C1(new_n594_), .C2(new_n597_), .ZN(new_n602_));
  AND3_X1   g401(.A1(new_n599_), .A2(new_n600_), .A3(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n600_), .B1(new_n599_), .B2(new_n602_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(G1325gat));
  NOR2_X1   g404(.A1(new_n286_), .A2(new_n288_), .ZN(new_n606_));
  OAI21_X1  g405(.A(G15gat), .B1(new_n585_), .B2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT41), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n446_), .A2(new_n574_), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n609_), .A2(G15gat), .A3(new_n606_), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n608_), .A2(new_n610_), .ZN(G1326gat));
  OAI21_X1  g410(.A(G22gat), .B1(new_n585_), .B2(new_n427_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT42), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n427_), .A2(G22gat), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n613_), .B1(new_n609_), .B2(new_n614_), .ZN(G1327gat));
  NOR2_X1   g414(.A1(new_n544_), .A2(new_n505_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n572_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n446_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(G29gat), .B1(new_n619_), .B2(new_n329_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n510_), .B1(new_n440_), .B2(new_n444_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(KEYINPUT43), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT43), .ZN(new_n623_));
  OAI211_X1 g422(.A(new_n623_), .B(new_n510_), .C1(new_n440_), .C2(new_n444_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n622_), .A2(new_n624_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n583_), .A2(new_n544_), .ZN(new_n626_));
  AOI21_X1  g425(.A(KEYINPUT44), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT44), .ZN(new_n628_));
  INV_X1    g427(.A(new_n626_), .ZN(new_n629_));
  AOI211_X1 g428(.A(new_n628_), .B(new_n629_), .C1(new_n622_), .C2(new_n624_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n627_), .A2(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n441_), .A2(new_n209_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n620_), .B1(new_n631_), .B2(new_n632_), .ZN(G1328gat));
  NOR2_X1   g432(.A1(new_n595_), .A2(G36gat), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n618_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT45), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n627_), .A2(new_n630_), .A3(new_n595_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n638_), .B1(new_n639_), .B2(new_n207_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT46), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  OAI211_X1 g441(.A(new_n638_), .B(KEYINPUT46), .C1(new_n639_), .C2(new_n207_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(G1329gat));
  INV_X1    g443(.A(G43gat), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n606_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n631_), .A2(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n645_), .B1(new_n618_), .B2(new_n606_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(KEYINPUT103), .B(KEYINPUT47), .ZN(new_n649_));
  AND3_X1   g448(.A1(new_n647_), .A2(new_n648_), .A3(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n649_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n650_), .A2(new_n651_), .ZN(G1330gat));
  INV_X1    g451(.A(new_n427_), .ZN(new_n653_));
  AOI21_X1  g452(.A(G50gat), .B1(new_n619_), .B2(new_n653_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n653_), .A2(G50gat), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n654_), .B1(new_n631_), .B2(new_n655_), .ZN(G1331gat));
  NOR3_X1   g455(.A1(new_n572_), .A2(new_n245_), .A3(new_n545_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n592_), .A2(new_n505_), .A3(new_n657_), .ZN(new_n658_));
  NOR3_X1   g457(.A1(new_n658_), .A2(new_n529_), .A3(new_n441_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT105), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n572_), .A2(new_n245_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n591_), .A2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(new_n546_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(KEYINPUT104), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT104), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n441_), .B1(new_n664_), .B2(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(G57gat), .B1(new_n666_), .B2(new_n668_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n660_), .A2(new_n669_), .ZN(G1332gat));
  OAI21_X1  g469(.A(G64gat), .B1(new_n658_), .B2(new_n595_), .ZN(new_n671_));
  XOR2_X1   g470(.A(KEYINPUT106), .B(KEYINPUT48), .Z(new_n672_));
  XNOR2_X1  g471(.A(new_n671_), .B(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n665_), .A2(new_n527_), .A3(new_n588_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(G1333gat));
  OAI21_X1  g474(.A(G71gat), .B1(new_n658_), .B2(new_n606_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT49), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n665_), .A2(new_n272_), .A3(new_n289_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1334gat));
  OAI21_X1  g478(.A(G78gat), .B1(new_n658_), .B2(new_n427_), .ZN(new_n680_));
  XOR2_X1   g479(.A(KEYINPUT107), .B(KEYINPUT50), .Z(new_n681_));
  XNOR2_X1  g480(.A(new_n680_), .B(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n665_), .A2(new_n520_), .A3(new_n653_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(G1335gat));
  INV_X1    g483(.A(new_n572_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n245_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n685_), .A2(new_n686_), .A3(new_n545_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n687_), .B1(new_n622_), .B2(new_n624_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(G85gat), .B1(new_n689_), .B2(new_n441_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n663_), .A2(new_n616_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n329_), .A2(new_n462_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n690_), .B1(new_n691_), .B2(new_n692_), .ZN(G1336gat));
  OAI21_X1  g492(.A(G92gat), .B1(new_n689_), .B2(new_n595_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n588_), .A2(new_n463_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n694_), .B1(new_n691_), .B2(new_n695_), .ZN(G1337gat));
  AND2_X1   g495(.A1(new_n458_), .A2(new_n460_), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n663_), .A2(new_n289_), .A3(new_n697_), .A4(new_n616_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT108), .Z(new_n699_));
  AOI21_X1  g498(.A(new_n472_), .B1(new_n688_), .B2(new_n289_), .ZN(new_n700_));
  OR3_X1    g499(.A1(new_n699_), .A2(KEYINPUT51), .A3(new_n700_), .ZN(new_n701_));
  OAI21_X1  g500(.A(KEYINPUT51), .B1(new_n699_), .B2(new_n700_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(G1338gat));
  AOI21_X1  g502(.A(new_n459_), .B1(new_n688_), .B2(new_n653_), .ZN(new_n704_));
  OR2_X1    g503(.A1(new_n704_), .A2(KEYINPUT52), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n427_), .A2(G106gat), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(KEYINPUT109), .B1(new_n691_), .B2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT109), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n663_), .A2(new_n709_), .A3(new_n616_), .A4(new_n706_), .ZN(new_n710_));
  AOI22_X1  g509(.A1(new_n704_), .A2(KEYINPUT52), .B1(new_n708_), .B2(new_n710_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(KEYINPUT110), .B(KEYINPUT53), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n705_), .A2(new_n711_), .A3(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n705_), .B2(new_n711_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n713_), .A2(new_n714_), .ZN(G1339gat));
  NOR3_X1   g514(.A1(new_n443_), .A2(new_n441_), .A3(new_n606_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT112), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n236_), .A2(new_n240_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n204_), .B1(new_n718_), .B2(new_n237_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n236_), .A2(G229gat), .A3(G233gat), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n719_), .B1(new_n234_), .B2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n244_), .A2(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n722_), .B1(new_n559_), .B2(new_n565_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n548_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n724_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n725_));
  OAI21_X1  g524(.A(KEYINPUT12), .B1(new_n488_), .B2(new_n540_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n552_), .A2(new_n551_), .A3(new_n553_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n725_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n557_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n729_));
  OAI22_X1  g528(.A1(new_n728_), .A2(KEYINPUT55), .B1(new_n729_), .B2(new_n724_), .ZN(new_n730_));
  OAI211_X1 g529(.A(KEYINPUT55), .B(new_n549_), .C1(new_n550_), .C2(new_n554_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  OAI211_X1 g531(.A(KEYINPUT56), .B(new_n564_), .C1(new_n730_), .C2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  OAI22_X1  g533(.A1(new_n550_), .A2(new_n554_), .B1(new_n553_), .B2(new_n552_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(new_n548_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT55), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n555_), .A2(new_n737_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n736_), .A2(new_n738_), .A3(new_n731_), .ZN(new_n739_));
  AOI21_X1  g538(.A(KEYINPUT56), .B1(new_n739_), .B2(new_n564_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n723_), .B1(new_n734_), .B2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT58), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  OAI211_X1 g542(.A(KEYINPUT58), .B(new_n723_), .C1(new_n734_), .C2(new_n740_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n743_), .A2(new_n510_), .A3(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT57), .ZN(new_n746_));
  INV_X1    g545(.A(new_n505_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n567_), .A2(new_n245_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n749_), .B1(new_n734_), .B2(new_n740_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n722_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n747_), .B1(new_n750_), .B2(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n746_), .B1(new_n753_), .B2(KEYINPUT111), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n564_), .B1(new_n730_), .B2(new_n732_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT56), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n748_), .B1(new_n757_), .B2(new_n733_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n505_), .B1(new_n758_), .B2(new_n751_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT111), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n745_), .B1(new_n754_), .B2(new_n761_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n759_), .A2(new_n746_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n545_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n546_), .A2(new_n686_), .A3(new_n572_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT54), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n717_), .A2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(KEYINPUT59), .ZN(new_n769_));
  INV_X1    g568(.A(new_n763_), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n743_), .A2(new_n510_), .A3(new_n744_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT57), .B1(new_n759_), .B2(new_n760_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n753_), .A2(KEYINPUT111), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n771_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT114), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n770_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n775_), .B(new_n745_), .C1(new_n754_), .C2(new_n761_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n545_), .B1(new_n776_), .B2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n766_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(KEYINPUT113), .B(KEYINPUT59), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n780_), .A2(new_n717_), .A3(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n769_), .A2(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(G113gat), .B1(new_n783_), .B2(new_n686_), .ZN(new_n784_));
  OR2_X1    g583(.A1(new_n686_), .A2(G113gat), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n784_), .B1(new_n768_), .B2(new_n785_), .ZN(G1340gat));
  OAI21_X1  g585(.A(G120gat), .B1(new_n783_), .B2(new_n572_), .ZN(new_n787_));
  INV_X1    g586(.A(G120gat), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n788_), .B1(new_n572_), .B2(KEYINPUT60), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n789_), .B1(KEYINPUT60), .B2(new_n788_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n787_), .B1(new_n768_), .B2(new_n790_), .ZN(G1341gat));
  OAI21_X1  g590(.A(G127gat), .B1(new_n783_), .B2(new_n545_), .ZN(new_n792_));
  OR2_X1    g591(.A1(new_n545_), .A2(G127gat), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n792_), .B1(new_n768_), .B2(new_n793_), .ZN(G1342gat));
  INV_X1    g593(.A(new_n510_), .ZN(new_n795_));
  OAI21_X1  g594(.A(G134gat), .B1(new_n783_), .B2(new_n795_), .ZN(new_n796_));
  OR2_X1    g595(.A1(new_n505_), .A2(G134gat), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n796_), .B1(new_n768_), .B2(new_n797_), .ZN(G1343gat));
  INV_X1    g597(.A(new_n767_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n595_), .A2(new_n329_), .A3(new_n653_), .ZN(new_n800_));
  NOR3_X1   g599(.A1(new_n799_), .A2(new_n289_), .A3(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(new_n245_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(KEYINPUT115), .B(G141gat), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n802_), .B(new_n803_), .ZN(G1344gat));
  NAND2_X1  g603(.A1(new_n801_), .A2(new_n685_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n805_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g605(.A1(new_n801_), .A2(new_n544_), .ZN(new_n807_));
  XOR2_X1   g606(.A(KEYINPUT61), .B(G155gat), .Z(new_n808_));
  XNOR2_X1  g607(.A(new_n807_), .B(new_n808_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(KEYINPUT116), .B(KEYINPUT117), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n809_), .B(new_n811_), .ZN(G1346gat));
  INV_X1    g611(.A(new_n801_), .ZN(new_n813_));
  OR3_X1    g612(.A1(new_n813_), .A2(G162gat), .A3(new_n505_), .ZN(new_n814_));
  OAI21_X1  g613(.A(G162gat), .B1(new_n813_), .B2(new_n795_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(G1347gat));
  INV_X1    g615(.A(KEYINPUT122), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT120), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n588_), .A2(new_n441_), .A3(new_n289_), .A4(new_n427_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n819_), .A2(new_n686_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n763_), .B1(new_n762_), .B2(KEYINPUT114), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n544_), .B1(new_n821_), .B2(new_n777_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n766_), .ZN(new_n823_));
  OAI211_X1 g622(.A(KEYINPUT118), .B(new_n820_), .C1(new_n822_), .C2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(G169gat), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT118), .B1(new_n780_), .B2(new_n820_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n818_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT118), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n821_), .A2(new_n777_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n823_), .B1(new_n829_), .B2(new_n545_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n820_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n828_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n832_), .A2(KEYINPUT120), .A3(G169gat), .A4(new_n824_), .ZN(new_n833_));
  XOR2_X1   g632(.A(KEYINPUT119), .B(KEYINPUT62), .Z(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n827_), .A2(new_n833_), .A3(new_n835_), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n818_), .B(new_n834_), .C1(new_n825_), .C2(new_n826_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n830_), .A2(new_n819_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(KEYINPUT22), .B(G169gat), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n245_), .A2(new_n839_), .ZN(new_n840_));
  XOR2_X1   g639(.A(new_n840_), .B(KEYINPUT121), .Z(new_n841_));
  NAND2_X1  g640(.A1(new_n838_), .A2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n837_), .A2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n817_), .B1(new_n836_), .B2(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n827_), .A2(new_n833_), .A3(new_n835_), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n845_), .A2(KEYINPUT122), .A3(new_n837_), .A4(new_n842_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n846_), .ZN(G1348gat));
  AOI21_X1  g646(.A(G176gat), .B1(new_n838_), .B2(new_n685_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n799_), .A2(new_n819_), .ZN(new_n849_));
  INV_X1    g648(.A(G176gat), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n572_), .A2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n851_), .ZN(new_n852_));
  OR2_X1    g651(.A1(new_n852_), .A2(KEYINPUT123), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(KEYINPUT123), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n848_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT124), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n855_), .B(new_n856_), .ZN(G1349gat));
  AOI21_X1  g656(.A(G183gat), .B1(new_n849_), .B2(new_n544_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n545_), .A2(new_n333_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n858_), .B1(new_n838_), .B2(new_n859_), .ZN(G1350gat));
  NAND3_X1  g659(.A1(new_n838_), .A2(new_n253_), .A3(new_n747_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n838_), .ZN(new_n862_));
  OAI21_X1  g661(.A(G190gat), .B1(new_n862_), .B2(new_n795_), .ZN(new_n863_));
  AND2_X1   g662(.A1(new_n863_), .A2(KEYINPUT125), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n863_), .A2(KEYINPUT125), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n861_), .B1(new_n864_), .B2(new_n865_), .ZN(G1351gat));
  NOR2_X1   g665(.A1(new_n799_), .A2(new_n289_), .ZN(new_n867_));
  AND2_X1   g666(.A1(new_n588_), .A2(new_n429_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n245_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g671(.A1(new_n869_), .A2(new_n572_), .ZN(new_n873_));
  INV_X1    g672(.A(G204gat), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n873_), .B1(KEYINPUT126), .B2(new_n874_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(KEYINPUT126), .B(G204gat), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(new_n873_), .B2(new_n876_), .ZN(G1353gat));
  NOR2_X1   g676(.A1(new_n869_), .A2(new_n545_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n879_));
  AND2_X1   g678(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n878_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n881_), .B1(new_n878_), .B2(new_n879_), .ZN(G1354gat));
  XOR2_X1   g681(.A(KEYINPUT127), .B(G218gat), .Z(new_n883_));
  NOR3_X1   g682(.A1(new_n869_), .A2(new_n795_), .A3(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n870_), .A2(new_n747_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n884_), .B1(new_n885_), .B2(new_n883_), .ZN(G1355gat));
endmodule


