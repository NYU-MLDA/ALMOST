//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 0 0 1 1 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 1 0 1 1 1 0 0 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 0 1 1 0 0 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n780_, new_n781_,
    new_n782_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n804_, new_n805_, new_n806_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n934_, new_n936_, new_n937_,
    new_n939_, new_n940_, new_n941_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n960_, new_n961_, new_n962_, new_n963_, new_n965_, new_n966_,
    new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_,
    new_n975_, new_n977_, new_n978_, new_n979_, new_n981_, new_n982_;
  OR2_X1    g000(.A1(KEYINPUT78), .A2(G183gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(KEYINPUT78), .A2(G183gat), .ZN(new_n203_));
  NAND3_X1  g002(.A1(new_n202_), .A2(KEYINPUT25), .A3(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT26), .ZN(new_n205_));
  OR3_X1    g004(.A1(new_n205_), .A2(KEYINPUT79), .A3(G190gat), .ZN(new_n206_));
  INV_X1    g005(.A(G190gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT26), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT79), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT25), .ZN(new_n210_));
  AOI22_X1  g009(.A1(new_n210_), .A2(G183gat), .B1(new_n205_), .B2(G190gat), .ZN(new_n211_));
  NAND4_X1  g010(.A1(new_n204_), .A2(new_n206_), .A3(new_n209_), .A4(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT23), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT23), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n215_), .A2(G183gat), .A3(G190gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  NOR3_X1   g016(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT24), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n219_), .B1(G169gat), .B2(G176gat), .ZN(new_n220_));
  INV_X1    g019(.A(G169gat), .ZN(new_n221_));
  INV_X1    g020(.A(G176gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n218_), .B1(new_n220_), .B2(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n212_), .A2(new_n217_), .A3(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT81), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT80), .B(KEYINPUT22), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n226_), .B1(new_n227_), .B2(new_n221_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT80), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n229_), .A2(KEYINPUT22), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT22), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n231_), .A2(KEYINPUT80), .ZN(new_n232_));
  OAI211_X1 g031(.A(KEYINPUT81), .B(G169gat), .C1(new_n230_), .C2(new_n232_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n231_), .A2(G169gat), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n234_), .A2(G176gat), .ZN(new_n235_));
  AND3_X1   g034(.A1(new_n228_), .A2(new_n233_), .A3(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n214_), .A2(new_n216_), .A3(KEYINPUT82), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT82), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n213_), .A2(new_n238_), .A3(KEYINPUT23), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n202_), .A2(new_n207_), .A3(new_n203_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n237_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G169gat), .A2(G176gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n225_), .B1(new_n236_), .B2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G71gat), .B(G99gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT83), .B(G43gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n244_), .B(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G227gat), .A2(G233gat), .ZN(new_n249_));
  XOR2_X1   g048(.A(new_n249_), .B(G15gat), .Z(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT30), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n248_), .B(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT84), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G127gat), .B(G134gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G113gat), .B(G120gat), .ZN(new_n256_));
  XOR2_X1   g055(.A(new_n255_), .B(new_n256_), .Z(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT31), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n254_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n258_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n260_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n259_), .B1(new_n254_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT102), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G1gat), .B(G29gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(G85gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT0), .B(G57gat), .ZN(new_n267_));
  XOR2_X1   g066(.A(new_n266_), .B(new_n267_), .Z(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G141gat), .B(G148gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G155gat), .A2(G162gat), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n271_), .A2(KEYINPUT1), .ZN(new_n272_));
  NOR2_X1   g071(.A1(G155gat), .A2(G162gat), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n271_), .B1(new_n273_), .B2(KEYINPUT1), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT85), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n272_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT1), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n277_), .B1(G155gat), .B2(G162gat), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n278_), .A2(KEYINPUT85), .A3(new_n271_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n270_), .B1(new_n276_), .B2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n271_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n281_), .A2(new_n273_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT3), .ZN(new_n284_));
  INV_X1    g083(.A(G141gat), .ZN(new_n285_));
  INV_X1    g084(.A(G148gat), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n284_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G141gat), .A2(G148gat), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT2), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  OAI21_X1  g089(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n291_));
  AND3_X1   g090(.A1(new_n287_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(KEYINPUT86), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT86), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n295_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n283_), .B1(new_n292_), .B2(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n257_), .B1(new_n280_), .B2(new_n298_), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n294_), .A2(new_n296_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n287_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n282_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n255_), .B(new_n256_), .ZN(new_n303_));
  AND3_X1   g102(.A1(new_n278_), .A2(KEYINPUT85), .A3(new_n271_), .ZN(new_n304_));
  AOI21_X1  g103(.A(KEYINPUT85), .B1(new_n278_), .B2(new_n271_), .ZN(new_n305_));
  NOR3_X1   g104(.A1(new_n304_), .A2(new_n305_), .A3(new_n272_), .ZN(new_n306_));
  OAI211_X1 g105(.A(new_n302_), .B(new_n303_), .C1(new_n306_), .C2(new_n270_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n299_), .A2(new_n307_), .A3(KEYINPUT4), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT4), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n257_), .B(new_n309_), .C1(new_n280_), .C2(new_n298_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G225gat), .A2(G233gat), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n311_), .B(KEYINPUT93), .Z(new_n312_));
  NAND4_X1  g111(.A1(new_n308_), .A2(KEYINPUT94), .A3(new_n310_), .A4(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n299_), .A2(new_n307_), .A3(new_n311_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n310_), .A2(new_n312_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(KEYINPUT94), .B1(new_n317_), .B2(new_n308_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n269_), .B1(new_n315_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT98), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT94), .ZN(new_n321_));
  INV_X1    g120(.A(new_n308_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n321_), .B1(new_n322_), .B2(new_n316_), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n323_), .A2(new_n268_), .A3(new_n314_), .A4(new_n313_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n319_), .A2(new_n320_), .A3(new_n324_), .ZN(new_n325_));
  OAI211_X1 g124(.A(KEYINPUT98), .B(new_n269_), .C1(new_n315_), .C2(new_n318_), .ZN(new_n326_));
  AND3_X1   g125(.A1(new_n325_), .A2(KEYINPUT100), .A3(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(KEYINPUT100), .B1(new_n325_), .B2(new_n326_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT27), .ZN(new_n330_));
  XOR2_X1   g129(.A(G8gat), .B(G36gat), .Z(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT18), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G64gat), .B(G92gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G226gat), .A2(G233gat), .ZN(new_n336_));
  XOR2_X1   g135(.A(new_n336_), .B(KEYINPUT19), .Z(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT20), .ZN(new_n338_));
  OR2_X1    g137(.A1(G197gat), .A2(G204gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G197gat), .A2(G204gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT21), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT88), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n341_), .A2(KEYINPUT88), .A3(new_n342_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n339_), .A2(KEYINPUT21), .A3(new_n340_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G211gat), .B(G218gat), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n345_), .A2(new_n346_), .A3(new_n347_), .A4(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n347_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n348_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n349_), .A2(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n338_), .B1(new_n244_), .B2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n218_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n237_), .A2(new_n355_), .A3(new_n239_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT91), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n237_), .A2(KEYINPUT91), .A3(new_n355_), .A4(new_n239_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n205_), .A2(G190gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n208_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT90), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT90), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n208_), .A2(new_n361_), .A3(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT25), .B(G183gat), .ZN(new_n367_));
  AOI22_X1  g166(.A1(new_n366_), .A2(new_n367_), .B1(new_n223_), .B2(new_n220_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n360_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n347_), .A2(new_n348_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n370_), .B1(new_n344_), .B2(new_n343_), .ZN(new_n371_));
  AOI22_X1  g170(.A1(new_n371_), .A2(new_n346_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n221_), .A2(KEYINPUT22), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT92), .B1(new_n234_), .B2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n221_), .A2(KEYINPUT22), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n231_), .A2(G169gat), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT92), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n375_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(G176gat), .B1(new_n374_), .B2(new_n378_), .ZN(new_n379_));
  OR2_X1    g178(.A1(G183gat), .A2(G190gat), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n215_), .B1(G183gat), .B2(G190gat), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n213_), .A2(KEYINPUT23), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n380_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(new_n242_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n379_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n369_), .A2(new_n372_), .A3(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n228_), .A2(new_n233_), .A3(new_n235_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n388_), .A2(new_n242_), .A3(new_n241_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n389_), .A2(new_n225_), .A3(new_n349_), .A4(new_n352_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n385_), .B1(new_n360_), .B2(new_n368_), .ZN(new_n391_));
  OAI211_X1 g190(.A(KEYINPUT20), .B(new_n390_), .C1(new_n391_), .C2(new_n372_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n337_), .ZN(new_n393_));
  AOI221_X4 g192(.A(new_n335_), .B1(new_n354_), .B2(new_n387_), .C1(new_n392_), .C2(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n372_), .B1(new_n369_), .B2(new_n386_), .ZN(new_n395_));
  OAI21_X1  g194(.A(KEYINPUT20), .B1(new_n244_), .B2(new_n353_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n393_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n354_), .A2(new_n387_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n334_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n330_), .B1(new_n394_), .B2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n397_), .A2(new_n398_), .A3(new_n334_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT101), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n392_), .A2(new_n393_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT97), .B(KEYINPUT20), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n404_), .B1(new_n244_), .B2(new_n353_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n337_), .B1(new_n405_), .B2(new_n387_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n335_), .B1(new_n403_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT101), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n397_), .A2(new_n408_), .A3(new_n398_), .A4(new_n334_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n402_), .A2(KEYINPUT27), .A3(new_n407_), .A4(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G22gat), .B(G50gat), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT28), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n280_), .A2(new_n298_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT29), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n413_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  NOR4_X1   g215(.A1(new_n280_), .A2(new_n298_), .A3(KEYINPUT28), .A4(KEYINPUT29), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n412_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n414_), .A2(new_n413_), .A3(new_n415_), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n302_), .B(new_n415_), .C1(new_n306_), .C2(new_n270_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(KEYINPUT28), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n419_), .A2(new_n421_), .A3(new_n411_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n418_), .A2(new_n422_), .ZN(new_n423_));
  XOR2_X1   g222(.A(G78gat), .B(G106gat), .Z(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT29), .B1(new_n280_), .B2(new_n298_), .ZN(new_n426_));
  INV_X1    g225(.A(G233gat), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n427_), .A2(KEYINPUT87), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(KEYINPUT87), .ZN(new_n429_));
  OAI21_X1  g228(.A(G228gat), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n426_), .A2(new_n353_), .A3(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n430_), .B1(new_n426_), .B2(new_n353_), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT89), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n423_), .A2(new_n425_), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n425_), .B1(new_n423_), .B2(new_n433_), .ZN(new_n436_));
  NOR3_X1   g235(.A1(new_n431_), .A2(new_n432_), .A3(KEYINPUT89), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NOR3_X1   g237(.A1(new_n435_), .A2(new_n436_), .A3(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n423_), .A2(new_n433_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(new_n424_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n437_), .B1(new_n441_), .B2(new_n434_), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n400_), .B(new_n410_), .C1(new_n439_), .C2(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n264_), .B1(new_n329_), .B2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n325_), .A2(new_n326_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT100), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n325_), .A2(KEYINPUT100), .A3(new_n326_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n439_), .A2(new_n442_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n410_), .A2(new_n400_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n449_), .A2(new_n451_), .A3(KEYINPUT102), .A4(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n444_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n334_), .A2(KEYINPUT32), .ZN(new_n456_));
  AND3_X1   g255(.A1(new_n397_), .A2(new_n398_), .A3(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n405_), .A2(new_n387_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(new_n393_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n369_), .A2(new_n386_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(new_n353_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT20), .ZN(new_n462_));
  INV_X1    g261(.A(new_n243_), .ZN(new_n463_));
  AND2_X1   g262(.A1(new_n224_), .A2(new_n217_), .ZN(new_n464_));
  AOI22_X1  g263(.A1(new_n463_), .A2(new_n388_), .B1(new_n212_), .B2(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n462_), .B1(new_n465_), .B2(new_n372_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n461_), .A2(new_n466_), .A3(new_n337_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n456_), .B1(new_n459_), .B2(new_n467_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n457_), .A2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n469_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n394_), .A2(new_n399_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n315_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT95), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n473_), .A2(KEYINPUT33), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n472_), .A2(new_n268_), .A3(new_n323_), .A4(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n324_), .A2(new_n474_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n308_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n299_), .A2(new_n307_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT96), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(new_n312_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n479_), .A2(new_n480_), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n269_), .B(new_n478_), .C1(new_n482_), .C2(new_n483_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n471_), .A2(new_n476_), .A3(new_n477_), .A4(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n470_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(new_n450_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT99), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT99), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n486_), .A2(new_n489_), .A3(new_n450_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n263_), .B1(new_n455_), .B2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT103), .ZN(new_n493_));
  NOR3_X1   g292(.A1(new_n263_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(new_n449_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n444_), .A2(new_n454_), .A3(new_n488_), .A4(new_n490_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT103), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n496_), .A2(new_n497_), .A3(new_n263_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n493_), .A2(new_n495_), .A3(new_n498_), .ZN(new_n499_));
  XOR2_X1   g298(.A(G29gat), .B(G36gat), .Z(new_n500_));
  XOR2_X1   g299(.A(G43gat), .B(G50gat), .Z(new_n501_));
  XOR2_X1   g300(.A(new_n500_), .B(new_n501_), .Z(new_n502_));
  XOR2_X1   g301(.A(new_n502_), .B(KEYINPUT15), .Z(new_n503_));
  INV_X1    g302(.A(G1gat), .ZN(new_n504_));
  INV_X1    g303(.A(G8gat), .ZN(new_n505_));
  OAI21_X1  g304(.A(KEYINPUT14), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT74), .ZN(new_n507_));
  OR2_X1    g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(new_n507_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G15gat), .B(G22gat), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n508_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  XOR2_X1   g310(.A(G1gat), .B(G8gat), .Z(new_n512_));
  XOR2_X1   g311(.A(new_n511_), .B(new_n512_), .Z(new_n513_));
  NAND2_X1  g312(.A1(new_n503_), .A2(new_n513_), .ZN(new_n514_));
  OR2_X1    g313(.A1(new_n513_), .A2(new_n502_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G229gat), .A2(G233gat), .ZN(new_n518_));
  XOR2_X1   g317(.A(new_n518_), .B(KEYINPUT76), .Z(new_n519_));
  NAND2_X1  g318(.A1(new_n517_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT77), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n513_), .B(new_n502_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n523_), .A2(G229gat), .A3(G233gat), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n517_), .A2(KEYINPUT77), .A3(new_n519_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n522_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G113gat), .B(G141gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G169gat), .B(G197gat), .ZN(new_n528_));
  XOR2_X1   g327(.A(new_n527_), .B(new_n528_), .Z(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n526_), .A2(new_n530_), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n522_), .A2(new_n524_), .A3(new_n525_), .A4(new_n529_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G57gat), .B(G64gat), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(KEYINPUT11), .ZN(new_n535_));
  XOR2_X1   g334(.A(G71gat), .B(G78gat), .Z(new_n536_));
  NOR2_X1   g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  AND2_X1   g336(.A1(new_n535_), .A2(new_n536_), .ZN(new_n538_));
  OR2_X1    g337(.A1(new_n534_), .A2(KEYINPUT11), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n537_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G231gat), .A2(G233gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT75), .ZN(new_n543_));
  OR2_X1    g342(.A1(new_n543_), .A2(new_n513_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n513_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT17), .ZN(new_n547_));
  XOR2_X1   g346(.A(G127gat), .B(G155gat), .Z(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT16), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G183gat), .B(G211gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  OR3_X1    g350(.A1(new_n546_), .A2(new_n547_), .A3(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(KEYINPUT17), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n546_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n552_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT37), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT35), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G232gat), .A2(G233gat), .ZN(new_n559_));
  XOR2_X1   g358(.A(new_n559_), .B(KEYINPUT34), .Z(new_n560_));
  XOR2_X1   g359(.A(KEYINPUT10), .B(G99gat), .Z(new_n561_));
  INV_X1    g360(.A(G106gat), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  XOR2_X1   g362(.A(G85gat), .B(G92gat), .Z(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT9), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT9), .ZN(new_n566_));
  INV_X1    g365(.A(G85gat), .ZN(new_n567_));
  INV_X1    g366(.A(G92gat), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G99gat), .A2(G106gat), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(KEYINPUT6), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT6), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n572_), .A2(G99gat), .A3(G106gat), .ZN(new_n573_));
  AOI22_X1  g372(.A1(new_n566_), .A2(new_n569_), .B1(new_n571_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT64), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n563_), .A2(new_n565_), .A3(new_n574_), .A4(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n563_), .A2(new_n565_), .A3(new_n574_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(KEYINPUT64), .ZN(new_n578_));
  NOR2_X1   g377(.A1(G99gat), .A2(G106gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT7), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n571_), .A2(new_n573_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT8), .ZN(new_n583_));
  AND3_X1   g382(.A1(new_n582_), .A2(new_n583_), .A3(new_n564_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n583_), .B1(new_n582_), .B2(new_n564_), .ZN(new_n585_));
  OAI211_X1 g384(.A(new_n576_), .B(new_n578_), .C1(new_n584_), .C2(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n586_), .A2(new_n502_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n560_), .A2(new_n558_), .ZN(new_n588_));
  XOR2_X1   g387(.A(new_n588_), .B(KEYINPUT72), .Z(new_n589_));
  NOR2_X1   g388(.A1(new_n587_), .A2(new_n589_), .ZN(new_n590_));
  AOI211_X1 g389(.A(new_n558_), .B(new_n560_), .C1(new_n590_), .C2(KEYINPUT71), .ZN(new_n591_));
  AND3_X1   g390(.A1(new_n578_), .A2(KEYINPUT65), .A3(new_n576_), .ZN(new_n592_));
  AOI21_X1  g391(.A(KEYINPUT65), .B1(new_n578_), .B2(new_n576_), .ZN(new_n593_));
  OAI22_X1  g392(.A1(new_n592_), .A2(new_n593_), .B1(new_n585_), .B2(new_n584_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(new_n503_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(new_n590_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n591_), .B(new_n596_), .ZN(new_n597_));
  XOR2_X1   g396(.A(G190gat), .B(G218gat), .Z(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT73), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G134gat), .B(G162gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT36), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n597_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n601_), .B(KEYINPUT36), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n597_), .A2(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n557_), .B1(new_n605_), .B2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n607_), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n609_), .A2(new_n604_), .A3(KEYINPUT37), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n556_), .B1(new_n608_), .B2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT69), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT66), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n584_), .A2(new_n585_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n578_), .A2(new_n576_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT65), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n578_), .A2(KEYINPUT65), .A3(new_n576_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n614_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n540_), .A2(KEYINPUT12), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n613_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(G230gat), .A2(G233gat), .ZN(new_n622_));
  INV_X1    g421(.A(new_n620_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n594_), .A2(KEYINPUT66), .A3(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(KEYINPUT12), .B1(new_n586_), .B2(new_n540_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n586_), .A2(new_n540_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n621_), .A2(new_n622_), .A3(new_n624_), .A4(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n622_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n586_), .A2(new_n540_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n629_), .B1(new_n630_), .B2(new_n626_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(G176gat), .B(G204gat), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT68), .ZN(new_n633_));
  XOR2_X1   g432(.A(KEYINPUT67), .B(KEYINPUT5), .Z(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(G120gat), .B(G148gat), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n635_), .B(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n628_), .A2(new_n631_), .A3(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n637_), .B1(new_n628_), .B2(new_n631_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n612_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n640_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n642_), .A2(KEYINPUT69), .A3(new_n638_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT13), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n641_), .A2(new_n643_), .A3(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n644_), .B1(new_n641_), .B2(new_n643_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(KEYINPUT70), .ZN(new_n649_));
  INV_X1    g448(.A(new_n647_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(new_n645_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT70), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n611_), .B1(new_n649_), .B2(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n499_), .A2(new_n533_), .A3(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT104), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n449_), .A2(G1gat), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n656_), .A2(new_n657_), .A3(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n658_), .ZN(new_n660_));
  OAI21_X1  g459(.A(KEYINPUT104), .B1(new_n655_), .B2(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n659_), .A2(KEYINPUT38), .A3(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n498_), .A2(new_n495_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n497_), .B1(new_n496_), .B2(new_n263_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n609_), .A2(new_n604_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n533_), .ZN(new_n668_));
  NOR3_X1   g467(.A1(new_n648_), .A2(new_n668_), .A3(new_n555_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(new_n670_));
  OAI21_X1  g469(.A(G1gat), .B1(new_n670_), .B2(new_n449_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n662_), .A2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n659_), .A2(new_n661_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT38), .ZN(new_n674_));
  AOI21_X1  g473(.A(KEYINPUT105), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT105), .ZN(new_n676_));
  AOI211_X1 g475(.A(new_n676_), .B(KEYINPUT38), .C1(new_n659_), .C2(new_n661_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n672_), .B1(new_n675_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT106), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n672_), .B(KEYINPUT106), .C1(new_n675_), .C2(new_n677_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(G1324gat));
  NAND3_X1  g481(.A1(new_n656_), .A2(new_n505_), .A3(new_n452_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n667_), .A2(new_n452_), .A3(new_n669_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(KEYINPUT107), .A2(KEYINPUT39), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n505_), .B1(KEYINPUT107), .B2(KEYINPUT39), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n684_), .A2(new_n685_), .A3(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n685_), .B1(new_n684_), .B2(new_n686_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n683_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  XOR2_X1   g489(.A(new_n690_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g490(.A(G15gat), .B1(new_n670_), .B2(new_n263_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT41), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n655_), .A2(G15gat), .A3(new_n263_), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n693_), .A2(new_n694_), .ZN(G1326gat));
  OAI21_X1  g494(.A(G22gat), .B1(new_n670_), .B2(new_n450_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT42), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n450_), .A2(G22gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n697_), .B1(new_n655_), .B2(new_n698_), .ZN(G1327gat));
  NOR2_X1   g498(.A1(new_n665_), .A2(new_n668_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n666_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n701_), .A2(new_n556_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n703_), .A2(new_n648_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n700_), .A2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(G29gat), .B1(new_n706_), .B2(new_n329_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n608_), .A2(new_n610_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n708_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(KEYINPUT43), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT43), .ZN(new_n711_));
  OAI211_X1 g510(.A(new_n711_), .B(new_n708_), .C1(new_n663_), .C2(new_n664_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n651_), .A2(new_n533_), .A3(new_n555_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  AOI21_X1  g514(.A(KEYINPUT44), .B1(new_n713_), .B2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n712_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n711_), .B1(new_n499_), .B2(new_n708_), .ZN(new_n718_));
  OAI211_X1 g517(.A(KEYINPUT44), .B(new_n715_), .C1(new_n717_), .C2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(KEYINPUT108), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n714_), .B1(new_n710_), .B2(new_n712_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT108), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n721_), .A2(new_n722_), .A3(KEYINPUT44), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n716_), .B1(new_n720_), .B2(new_n723_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n329_), .A2(G29gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n707_), .B1(new_n724_), .B2(new_n725_), .ZN(G1328gat));
  INV_X1    g525(.A(KEYINPUT46), .ZN(new_n727_));
  INV_X1    g526(.A(G36gat), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n720_), .A2(new_n723_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n452_), .B1(new_n721_), .B2(KEYINPUT44), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n728_), .B1(new_n729_), .B2(new_n731_), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n700_), .A2(new_n728_), .A3(new_n452_), .A4(new_n704_), .ZN(new_n733_));
  XOR2_X1   g532(.A(KEYINPUT109), .B(KEYINPUT45), .Z(new_n734_));
  XNOR2_X1  g533(.A(new_n733_), .B(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n727_), .B1(new_n732_), .B2(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n730_), .B1(new_n720_), .B2(new_n723_), .ZN(new_n738_));
  OAI211_X1 g537(.A(KEYINPUT46), .B(new_n735_), .C1(new_n738_), .C2(new_n728_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(G1329gat));
  INV_X1    g539(.A(G43gat), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n263_), .A2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  AOI211_X1 g542(.A(new_n743_), .B(new_n716_), .C1(new_n720_), .C2(new_n723_), .ZN(new_n744_));
  AOI21_X1  g543(.A(G43gat), .B1(new_n706_), .B2(new_n262_), .ZN(new_n745_));
  OAI21_X1  g544(.A(KEYINPUT47), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n724_), .A2(new_n742_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT47), .ZN(new_n748_));
  INV_X1    g547(.A(new_n745_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n747_), .A2(new_n748_), .A3(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n746_), .A2(new_n750_), .ZN(G1330gat));
  AOI21_X1  g550(.A(G50gat), .B1(new_n706_), .B2(new_n451_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n451_), .A2(G50gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n724_), .B2(new_n753_), .ZN(G1331gat));
  INV_X1    g553(.A(new_n653_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n649_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n555_), .A2(new_n533_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n667_), .A2(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(G57gat), .B1(new_n760_), .B2(new_n449_), .ZN(new_n761_));
  OAI21_X1  g560(.A(KEYINPUT110), .B1(new_n665_), .B2(new_n533_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT110), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n499_), .A2(new_n763_), .A3(new_n668_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n762_), .A2(new_n764_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n611_), .A2(new_n651_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  OR2_X1    g566(.A1(new_n449_), .A2(G57gat), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n761_), .B1(new_n767_), .B2(new_n768_), .ZN(G1332gat));
  INV_X1    g568(.A(new_n767_), .ZN(new_n770_));
  INV_X1    g569(.A(G64gat), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n770_), .A2(new_n771_), .A3(new_n452_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n760_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n771_), .B1(new_n773_), .B2(new_n452_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT48), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n774_), .A2(new_n775_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n772_), .B1(new_n777_), .B2(new_n778_), .ZN(G1333gat));
  OAI21_X1  g578(.A(G71gat), .B1(new_n760_), .B2(new_n263_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT49), .ZN(new_n781_));
  OR2_X1    g580(.A1(new_n263_), .A2(G71gat), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n781_), .B1(new_n767_), .B2(new_n782_), .ZN(G1334gat));
  INV_X1    g582(.A(G78gat), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n770_), .A2(new_n784_), .A3(new_n451_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n784_), .B1(new_n773_), .B2(new_n451_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT50), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n786_), .A2(new_n787_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n785_), .B1(new_n789_), .B2(new_n790_), .ZN(G1335gat));
  NOR3_X1   g590(.A1(new_n651_), .A2(new_n533_), .A3(new_n556_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n713_), .A2(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n793_), .A2(G85gat), .A3(new_n329_), .ZN(new_n794_));
  NOR3_X1   g593(.A1(new_n755_), .A2(new_n756_), .A3(new_n703_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n765_), .A2(new_n329_), .A3(new_n795_), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n796_), .A2(KEYINPUT111), .A3(new_n567_), .ZN(new_n797_));
  AOI21_X1  g596(.A(KEYINPUT111), .B1(new_n796_), .B2(new_n567_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n794_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT112), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  OAI211_X1 g600(.A(KEYINPUT112), .B(new_n794_), .C1(new_n797_), .C2(new_n798_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(G1336gat));
  AND2_X1   g602(.A1(new_n765_), .A2(new_n795_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n804_), .A2(new_n568_), .A3(new_n452_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n793_), .A2(new_n452_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n805_), .B1(new_n806_), .B2(new_n568_), .ZN(G1337gat));
  NAND2_X1  g606(.A1(new_n793_), .A2(new_n262_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(G99gat), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n262_), .A2(new_n561_), .ZN(new_n810_));
  AOI22_X1  g609(.A1(new_n804_), .A2(new_n810_), .B1(KEYINPUT113), .B2(KEYINPUT51), .ZN(new_n811_));
  OR2_X1    g610(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n812_));
  AND3_X1   g611(.A1(new_n809_), .A2(new_n811_), .A3(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n812_), .B1(new_n809_), .B2(new_n811_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n813_), .A2(new_n814_), .ZN(G1338gat));
  NAND3_X1  g614(.A1(new_n804_), .A2(new_n562_), .A3(new_n451_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n713_), .A2(new_n451_), .A3(new_n792_), .ZN(new_n817_));
  XOR2_X1   g616(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n818_));
  AND3_X1   g617(.A1(new_n817_), .A2(G106gat), .A3(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n818_), .B1(new_n817_), .B2(G106gat), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n816_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(KEYINPUT53), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT53), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n816_), .B(new_n823_), .C1(new_n819_), .C2(new_n820_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n822_), .A2(new_n824_), .ZN(G1339gat));
  NAND2_X1  g624(.A1(new_n494_), .A2(new_n329_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n516_), .A2(new_n519_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n529_), .B1(new_n523_), .B2(new_n519_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n827_), .B1(KEYINPUT118), .B2(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n829_), .B1(KEYINPUT118), .B2(new_n828_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n830_), .A2(new_n532_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n831_), .A2(new_n638_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT55), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n628_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT116), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  OR2_X1    g635(.A1(new_n628_), .A2(new_n833_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n628_), .A2(KEYINPUT116), .A3(new_n833_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n621_), .A2(new_n624_), .A3(new_n627_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n629_), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n836_), .A2(new_n837_), .A3(new_n838_), .A4(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n637_), .ZN(new_n842_));
  AOI21_X1  g641(.A(KEYINPUT56), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n841_), .A2(KEYINPUT56), .A3(new_n842_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n832_), .B1(new_n843_), .B2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT58), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n832_), .B(KEYINPUT58), .C1(new_n843_), .C2(new_n845_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n848_), .A2(new_n708_), .A3(new_n849_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n668_), .A2(new_n639_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n844_), .B1(new_n843_), .B2(KEYINPUT117), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n841_), .A2(new_n842_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT56), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n853_), .A2(KEYINPUT117), .A3(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n851_), .B1(new_n852_), .B2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n641_), .A2(new_n643_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n831_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n666_), .B1(new_n856_), .B2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n850_), .B1(new_n859_), .B2(KEYINPUT57), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT57), .ZN(new_n861_));
  AOI211_X1 g660(.A(new_n861_), .B(new_n666_), .C1(new_n856_), .C2(new_n858_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n555_), .B1(new_n860_), .B2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n666_), .A2(new_n557_), .ZN(new_n864_));
  OAI21_X1  g663(.A(KEYINPUT37), .B1(new_n609_), .B2(new_n604_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n758_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT115), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n866_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(KEYINPUT115), .B1(new_n651_), .B2(new_n758_), .ZN(new_n870_));
  OAI21_X1  g669(.A(KEYINPUT54), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n867_), .A2(new_n868_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n651_), .A2(KEYINPUT115), .A3(new_n758_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n872_), .A2(new_n873_), .A3(new_n874_), .A4(new_n866_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n871_), .A2(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n826_), .B1(new_n863_), .B2(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(G113gat), .B1(new_n877_), .B2(new_n533_), .ZN(new_n878_));
  OR2_X1    g677(.A1(new_n878_), .A2(KEYINPUT119), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(KEYINPUT119), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n863_), .A2(new_n876_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n826_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(KEYINPUT59), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n826_), .A2(KEYINPUT59), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n862_), .B1(new_n860_), .B2(KEYINPUT120), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT120), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n850_), .B(new_n887_), .C1(new_n859_), .C2(KEYINPUT57), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n556_), .B1(new_n886_), .B2(new_n888_), .ZN(new_n889_));
  AND2_X1   g688(.A1(new_n871_), .A2(new_n875_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n885_), .B1(new_n889_), .B2(new_n890_), .ZN(new_n891_));
  AND2_X1   g690(.A1(new_n884_), .A2(new_n891_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(KEYINPUT121), .B(G113gat), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n533_), .A2(new_n893_), .ZN(new_n894_));
  XOR2_X1   g693(.A(new_n894_), .B(KEYINPUT122), .Z(new_n895_));
  AOI22_X1  g694(.A1(new_n879_), .A2(new_n880_), .B1(new_n892_), .B2(new_n895_), .ZN(G1340gat));
  INV_X1    g695(.A(KEYINPUT124), .ZN(new_n897_));
  INV_X1    g696(.A(new_n885_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n860_), .A2(KEYINPUT120), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n859_), .A2(KEYINPUT57), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n899_), .A2(new_n900_), .A3(new_n888_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n555_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n898_), .B1(new_n902_), .B2(new_n876_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT59), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n757_), .B1(new_n877_), .B2(new_n904_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n897_), .B1(new_n903_), .B2(new_n905_), .ZN(new_n906_));
  NAND4_X1  g705(.A1(new_n884_), .A2(new_n891_), .A3(KEYINPUT124), .A4(new_n757_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n906_), .A2(new_n907_), .A3(G120gat), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n651_), .A2(KEYINPUT60), .ZN(new_n909_));
  MUX2_X1   g708(.A(new_n909_), .B(KEYINPUT60), .S(G120gat), .Z(new_n910_));
  AND2_X1   g709(.A1(new_n877_), .A2(new_n910_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(KEYINPUT123), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n908_), .A2(new_n912_), .ZN(G1341gat));
  INV_X1    g712(.A(G127gat), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n877_), .A2(new_n914_), .A3(new_n556_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n884_), .A2(new_n891_), .A3(new_n556_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n916_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n915_), .B1(new_n917_), .B2(new_n914_), .ZN(G1342gat));
  INV_X1    g717(.A(G134gat), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n919_), .B1(new_n883_), .B2(new_n701_), .ZN(new_n920_));
  OR2_X1    g719(.A1(new_n920_), .A2(KEYINPUT125), .ZN(new_n921_));
  NAND4_X1  g720(.A1(new_n884_), .A2(new_n891_), .A3(G134gat), .A4(new_n708_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n920_), .A2(KEYINPUT125), .ZN(new_n923_));
  AND3_X1   g722(.A1(new_n921_), .A2(new_n922_), .A3(new_n923_), .ZN(G1343gat));
  AND2_X1   g723(.A1(new_n856_), .A2(new_n858_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n861_), .B1(new_n925_), .B2(new_n666_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n926_), .A2(new_n900_), .A3(new_n850_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n890_), .B1(new_n927_), .B2(new_n555_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n928_), .A2(new_n262_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n449_), .A2(new_n443_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n929_), .A2(new_n533_), .A3(new_n930_), .ZN(new_n931_));
  XOR2_X1   g730(.A(KEYINPUT126), .B(G141gat), .Z(new_n932_));
  XNOR2_X1  g731(.A(new_n931_), .B(new_n932_), .ZN(G1344gat));
  NAND3_X1  g732(.A1(new_n929_), .A2(new_n757_), .A3(new_n930_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n934_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g734(.A1(new_n929_), .A2(new_n556_), .A3(new_n930_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(KEYINPUT61), .B(G155gat), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n936_), .B(new_n937_), .ZN(G1346gat));
  INV_X1    g737(.A(G162gat), .ZN(new_n939_));
  NAND4_X1  g738(.A1(new_n929_), .A2(new_n939_), .A3(new_n666_), .A4(new_n930_), .ZN(new_n940_));
  AND3_X1   g739(.A1(new_n929_), .A2(new_n708_), .A3(new_n930_), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n940_), .B1(new_n941_), .B2(new_n939_), .ZN(G1347gat));
  NOR2_X1   g741(.A1(new_n329_), .A2(new_n453_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n943_), .A2(new_n262_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n944_), .A2(new_n451_), .ZN(new_n945_));
  OAI211_X1 g744(.A(new_n533_), .B(new_n945_), .C1(new_n889_), .C2(new_n890_), .ZN(new_n946_));
  INV_X1    g745(.A(KEYINPUT62), .ZN(new_n947_));
  AND3_X1   g746(.A1(new_n946_), .A2(new_n947_), .A3(G169gat), .ZN(new_n948_));
  AND2_X1   g747(.A1(new_n374_), .A2(new_n378_), .ZN(new_n949_));
  OR2_X1    g748(.A1(new_n946_), .A2(new_n949_), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n947_), .B1(new_n946_), .B2(G169gat), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n948_), .B1(new_n950_), .B2(new_n951_), .ZN(G1348gat));
  NAND2_X1  g751(.A1(new_n902_), .A2(new_n876_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n953_), .A2(new_n945_), .ZN(new_n954_));
  INV_X1    g753(.A(new_n954_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n955_), .A2(new_n648_), .ZN(new_n956_));
  NOR2_X1   g755(.A1(new_n928_), .A2(new_n451_), .ZN(new_n957_));
  NOR4_X1   g756(.A1(new_n755_), .A2(new_n756_), .A3(new_n222_), .A4(new_n944_), .ZN(new_n958_));
  AOI22_X1  g757(.A1(new_n956_), .A2(new_n222_), .B1(new_n957_), .B2(new_n958_), .ZN(G1349gat));
  NAND2_X1  g758(.A1(new_n202_), .A2(new_n203_), .ZN(new_n960_));
  NOR2_X1   g759(.A1(new_n944_), .A2(new_n555_), .ZN(new_n961_));
  AOI21_X1  g760(.A(new_n960_), .B1(new_n957_), .B2(new_n961_), .ZN(new_n962_));
  NOR2_X1   g761(.A1(new_n555_), .A2(new_n367_), .ZN(new_n963_));
  AOI21_X1  g762(.A(new_n962_), .B1(new_n955_), .B2(new_n963_), .ZN(G1350gat));
  OAI21_X1  g763(.A(G190gat), .B1(new_n954_), .B2(new_n866_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n666_), .A2(new_n366_), .ZN(new_n966_));
  OAI21_X1  g765(.A(new_n965_), .B1(new_n954_), .B2(new_n966_), .ZN(G1351gat));
  XNOR2_X1  g766(.A(KEYINPUT127), .B(G197gat), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n943_), .A2(new_n451_), .ZN(new_n969_));
  NOR3_X1   g768(.A1(new_n928_), .A2(new_n262_), .A3(new_n969_), .ZN(new_n970_));
  INV_X1    g769(.A(new_n970_), .ZN(new_n971_));
  OAI21_X1  g770(.A(new_n968_), .B1(new_n971_), .B2(new_n668_), .ZN(new_n972_));
  OAI211_X1 g771(.A(new_n970_), .B(new_n533_), .C1(KEYINPUT127), .C2(G197gat), .ZN(new_n973_));
  AND2_X1   g772(.A1(new_n972_), .A2(new_n973_), .ZN(G1352gat));
  NAND2_X1  g773(.A1(new_n970_), .A2(new_n757_), .ZN(new_n975_));
  XNOR2_X1  g774(.A(new_n975_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g775(.A(KEYINPUT63), .B(G211gat), .C1(new_n970_), .C2(new_n556_), .ZN(new_n977_));
  NOR2_X1   g776(.A1(new_n971_), .A2(new_n555_), .ZN(new_n978_));
  XOR2_X1   g777(.A(KEYINPUT63), .B(G211gat), .Z(new_n979_));
  AOI21_X1  g778(.A(new_n977_), .B1(new_n978_), .B2(new_n979_), .ZN(G1354gat));
  OR3_X1    g779(.A1(new_n971_), .A2(G218gat), .A3(new_n701_), .ZN(new_n981_));
  OAI21_X1  g780(.A(G218gat), .B1(new_n971_), .B2(new_n866_), .ZN(new_n982_));
  NAND2_X1  g781(.A1(new_n981_), .A2(new_n982_), .ZN(G1355gat));
endmodule


