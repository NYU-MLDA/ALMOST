//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 1 0 0 1 0 0 0 0 1 1 0 0 0 1 0 1 1 1 0 1 0 1 1 1 1 0 0 0 0 1 0 0 0 1 0 0 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n855_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n862_, new_n863_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n903_, new_n904_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n913_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_, new_n925_, new_n926_;
  NAND2_X1  g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202_));
  OAI21_X1  g001(.A(KEYINPUT84), .B1(G155gat), .B2(G162gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  NOR3_X1   g003(.A1(KEYINPUT84), .A2(G155gat), .A3(G162gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(new_n202_), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G141gat), .ZN(new_n207_));
  INV_X1    g006(.A(G148gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n207_), .A2(new_n208_), .A3(KEYINPUT3), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT3), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n210_), .B1(G141gat), .B2(G148gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G141gat), .A2(G148gat), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  AOI22_X1  g012(.A1(new_n209_), .A2(new_n211_), .B1(new_n213_), .B2(KEYINPUT2), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(KEYINPUT83), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT83), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n216_), .A2(G141gat), .A3(G148gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT2), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n215_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n206_), .B1(new_n214_), .B2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n207_), .A2(new_n208_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n215_), .A2(new_n217_), .A3(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n205_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(new_n203_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n202_), .A2(KEYINPUT1), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT1), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n226_), .A2(G155gat), .A3(G162gat), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n222_), .B1(new_n224_), .B2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT85), .B1(new_n220_), .B2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n209_), .A2(new_n211_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n213_), .A2(KEYINPUT2), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n219_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n233_), .A2(new_n224_), .A3(new_n202_), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n225_), .B(new_n227_), .C1(new_n204_), .C2(new_n205_), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n235_), .A2(new_n215_), .A3(new_n217_), .A4(new_n221_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT85), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n234_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  XOR2_X1   g037(.A(G127gat), .B(G134gat), .Z(new_n239_));
  XOR2_X1   g038(.A(G113gat), .B(G120gat), .Z(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n230_), .A2(new_n238_), .A3(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT94), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n220_), .A2(new_n229_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n244_), .B1(new_n245_), .B2(new_n241_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n243_), .A2(new_n246_), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n230_), .A2(new_n238_), .A3(new_n244_), .A4(new_n242_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n247_), .A2(KEYINPUT4), .A3(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT4), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n243_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n249_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G225gat), .A2(G233gat), .ZN(new_n253_));
  XOR2_X1   g052(.A(new_n253_), .B(KEYINPUT95), .Z(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G1gat), .B(G29gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(G85gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT0), .B(G57gat), .ZN(new_n258_));
  XOR2_X1   g057(.A(new_n257_), .B(new_n258_), .Z(new_n259_));
  AOI21_X1  g058(.A(new_n254_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n255_), .A2(new_n259_), .A3(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT99), .ZN(new_n263_));
  INV_X1    g062(.A(new_n259_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n254_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n265_), .B1(new_n249_), .B2(new_n251_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n264_), .B1(new_n266_), .B2(new_n260_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n262_), .A2(new_n263_), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(G197gat), .ZN(new_n269_));
  INV_X1    g068(.A(G204gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G197gat), .A2(G204gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT21), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT88), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n273_), .A2(KEYINPUT88), .A3(new_n274_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n271_), .A2(KEYINPUT21), .A3(new_n272_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G211gat), .B(G218gat), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n277_), .A2(new_n278_), .A3(new_n279_), .A4(new_n280_), .ZN(new_n281_));
  OR2_X1    g080(.A1(new_n279_), .A2(new_n280_), .ZN(new_n282_));
  AND2_X1   g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT25), .B(G183gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(KEYINPUT26), .B(G190gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT78), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(G169gat), .A2(G176gat), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  OR2_X1    g089(.A1(new_n290_), .A2(KEYINPUT24), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G183gat), .A2(G190gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT23), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G169gat), .A2(G176gat), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n290_), .A2(KEYINPUT24), .A3(new_n294_), .ZN(new_n295_));
  AND3_X1   g094(.A1(new_n291_), .A2(new_n293_), .A3(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n288_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT80), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT22), .B(G169gat), .ZN(new_n299_));
  INV_X1    g098(.A(G176gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT79), .ZN(new_n302_));
  AOI22_X1  g101(.A1(new_n301_), .A2(new_n302_), .B1(G169gat), .B2(G176gat), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n299_), .A2(KEYINPUT79), .A3(new_n300_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n298_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n301_), .A2(new_n302_), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n306_), .A2(new_n298_), .A3(new_n294_), .A4(new_n304_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT23), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n292_), .A2(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n310_));
  OAI211_X1 g109(.A(new_n309_), .B(new_n310_), .C1(G183gat), .C2(G190gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n307_), .A2(new_n311_), .ZN(new_n312_));
  OAI211_X1 g111(.A(new_n283_), .B(new_n297_), .C1(new_n305_), .C2(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n301_), .A2(new_n311_), .A3(new_n294_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  OR2_X1    g114(.A1(KEYINPUT92), .A2(KEYINPUT24), .ZN(new_n316_));
  NAND2_X1  g115(.A1(KEYINPUT92), .A2(KEYINPUT24), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n318_), .A2(new_n290_), .A3(new_n294_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n316_), .A2(new_n289_), .A3(new_n317_), .ZN(new_n320_));
  AND3_X1   g119(.A1(new_n319_), .A2(new_n293_), .A3(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(G190gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(KEYINPUT26), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT26), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(G190gat), .ZN(new_n325_));
  AND3_X1   g124(.A1(new_n323_), .A2(new_n325_), .A3(KEYINPUT91), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(KEYINPUT91), .B1(new_n323_), .B2(new_n325_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n327_), .A2(new_n284_), .A3(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT93), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n321_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n332_));
  XOR2_X1   g131(.A(KEYINPUT25), .B(G183gat), .Z(new_n333_));
  NOR3_X1   g132(.A1(new_n326_), .A2(new_n328_), .A3(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n319_), .A2(new_n293_), .A3(new_n320_), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT93), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n315_), .B1(new_n332_), .B2(new_n336_), .ZN(new_n337_));
  OAI211_X1 g136(.A(new_n313_), .B(KEYINPUT20), .C1(new_n283_), .C2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G226gat), .A2(G233gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n338_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n341_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(KEYINPUT20), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n344_), .B1(new_n337_), .B2(new_n283_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n297_), .B1(new_n312_), .B2(new_n305_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n281_), .A2(new_n282_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n345_), .A2(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G8gat), .B(G36gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT18), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G64gat), .B(G92gat), .ZN(new_n352_));
  XOR2_X1   g151(.A(new_n351_), .B(new_n352_), .Z(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT32), .ZN(new_n354_));
  AND3_X1   g153(.A1(new_n342_), .A2(new_n349_), .A3(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n314_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n356_));
  OAI21_X1  g155(.A(KEYINPUT20), .B1(new_n347_), .B2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT98), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  OAI211_X1 g158(.A(KEYINPUT98), .B(KEYINPUT20), .C1(new_n347_), .C2(new_n356_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n359_), .A2(new_n348_), .A3(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(new_n341_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT20), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n331_), .B1(new_n321_), .B2(new_n330_), .ZN(new_n364_));
  NOR3_X1   g163(.A1(new_n334_), .A2(new_n335_), .A3(KEYINPUT93), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n314_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n363_), .B1(new_n366_), .B2(new_n347_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n367_), .A2(new_n343_), .A3(new_n313_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n354_), .B1(new_n362_), .B2(new_n368_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n355_), .A2(new_n369_), .ZN(new_n370_));
  OAI211_X1 g169(.A(KEYINPUT99), .B(new_n264_), .C1(new_n266_), .C2(new_n260_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n268_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT100), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n353_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n343_), .B1(new_n367_), .B2(new_n313_), .ZN(new_n376_));
  AND2_X1   g175(.A1(new_n345_), .A2(new_n348_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n375_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n342_), .A2(new_n349_), .A3(new_n353_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n254_), .B1(new_n249_), .B2(new_n251_), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n247_), .A2(new_n248_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n264_), .B1(new_n381_), .B2(new_n265_), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n378_), .B(new_n379_), .C1(new_n380_), .C2(new_n382_), .ZN(new_n383_));
  XOR2_X1   g182(.A(KEYINPUT97), .B(KEYINPUT33), .Z(new_n384_));
  NOR2_X1   g183(.A1(new_n266_), .A2(new_n260_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n384_), .B1(new_n385_), .B2(new_n259_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n383_), .A2(new_n386_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n255_), .A2(KEYINPUT33), .A3(new_n259_), .A4(new_n261_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT96), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n385_), .A2(KEYINPUT96), .A3(KEYINPUT33), .A4(new_n259_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n387_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT29), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n347_), .B1(new_n245_), .B2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G228gat), .A2(G233gat), .ZN(new_n396_));
  XOR2_X1   g195(.A(new_n396_), .B(KEYINPUT87), .Z(new_n397_));
  NAND2_X1  g196(.A1(new_n395_), .A2(new_n397_), .ZN(new_n398_));
  OR2_X1    g197(.A1(new_n283_), .A2(new_n397_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n230_), .A2(new_n238_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n400_), .A2(new_n394_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n398_), .B1(new_n399_), .B2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G78gat), .B(G106gat), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n402_), .B(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT89), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n406_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n400_), .A2(new_n394_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  XOR2_X1   g210(.A(G22gat), .B(G50gat), .Z(new_n412_));
  INV_X1    g211(.A(new_n410_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n400_), .A2(new_n394_), .A3(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n411_), .A2(new_n412_), .A3(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n411_), .A2(new_n414_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n412_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n405_), .A2(new_n408_), .A3(new_n415_), .A4(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n402_), .B(new_n403_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n418_), .A2(new_n415_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n420_), .B1(new_n421_), .B2(new_n407_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n419_), .A2(new_n422_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n268_), .A2(new_n370_), .A3(KEYINPUT100), .A4(new_n371_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n374_), .A2(new_n393_), .A3(new_n423_), .A4(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT30), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n346_), .A2(new_n426_), .ZN(new_n427_));
  XOR2_X1   g226(.A(G15gat), .B(G43gat), .Z(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n297_), .B(KEYINPUT30), .C1(new_n312_), .C2(new_n305_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n427_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n429_), .B1(new_n427_), .B2(new_n430_), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT31), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n427_), .A2(new_n430_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n428_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT31), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n436_), .A2(new_n437_), .A3(new_n431_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G227gat), .A2(G233gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(G71gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(G99gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(KEYINPUT81), .B(KEYINPUT82), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n441_), .B(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(new_n242_), .ZN(new_n444_));
  AND3_X1   g243(.A1(new_n434_), .A2(new_n438_), .A3(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n444_), .B1(new_n434_), .B2(new_n438_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n378_), .A2(new_n379_), .ZN(new_n448_));
  XOR2_X1   g247(.A(KEYINPUT101), .B(KEYINPUT27), .Z(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT27), .ZN(new_n451_));
  AOI22_X1  g250(.A1(new_n338_), .A2(new_n341_), .B1(new_n348_), .B2(new_n345_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n451_), .B1(new_n452_), .B2(new_n353_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n362_), .A2(new_n368_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(new_n375_), .ZN(new_n455_));
  AOI22_X1  g254(.A1(new_n448_), .A2(new_n450_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n268_), .A2(new_n371_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n423_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n447_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n456_), .A2(new_n447_), .A3(new_n423_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  AOI22_X1  g261(.A1(new_n425_), .A2(new_n460_), .B1(new_n457_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G229gat), .A2(G233gat), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G29gat), .B(G36gat), .ZN(new_n466_));
  AND2_X1   g265(.A1(new_n466_), .A2(KEYINPUT72), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n466_), .A2(KEYINPUT72), .ZN(new_n468_));
  XOR2_X1   g267(.A(G43gat), .B(G50gat), .Z(new_n469_));
  OR3_X1    g268(.A1(new_n467_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n469_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G15gat), .B(G22gat), .ZN(new_n473_));
  INV_X1    g272(.A(G1gat), .ZN(new_n474_));
  INV_X1    g273(.A(G8gat), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT14), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n473_), .A2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G1gat), .B(G8gat), .ZN(new_n478_));
  XOR2_X1   g277(.A(new_n477_), .B(new_n478_), .Z(new_n479_));
  AOI21_X1  g278(.A(new_n465_), .B1(new_n472_), .B2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n472_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT15), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT15), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n472_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n479_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n482_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n480_), .A2(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(KEYINPUT77), .B1(new_n472_), .B2(new_n479_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n488_), .B1(new_n472_), .B2(new_n479_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n481_), .A2(KEYINPUT77), .A3(new_n485_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n489_), .A2(new_n465_), .A3(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n487_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G113gat), .B(G141gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G169gat), .B(G197gat), .ZN(new_n494_));
  XOR2_X1   g293(.A(new_n493_), .B(new_n494_), .Z(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n492_), .A2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n487_), .A2(new_n491_), .A3(new_n495_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n463_), .A2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G57gat), .B(G64gat), .ZN(new_n502_));
  OR2_X1    g301(.A1(new_n502_), .A2(KEYINPUT11), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(KEYINPUT11), .ZN(new_n504_));
  XOR2_X1   g303(.A(G71gat), .B(G78gat), .Z(new_n505_));
  NAND3_X1  g304(.A1(new_n503_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  OR2_X1    g305(.A1(new_n504_), .A2(new_n505_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  AND2_X1   g307(.A1(G231gat), .A2(G233gat), .ZN(new_n509_));
  XOR2_X1   g308(.A(new_n508_), .B(new_n509_), .Z(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(KEYINPUT76), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(new_n485_), .ZN(new_n512_));
  XOR2_X1   g311(.A(G127gat), .B(G155gat), .Z(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT16), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G183gat), .B(G211gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT17), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n512_), .A2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n511_), .B(new_n479_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n516_), .B(KEYINPUT17), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n519_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(G85gat), .ZN(new_n525_));
  INV_X1    g324(.A(G92gat), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G85gat), .A2(G92gat), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n527_), .A2(KEYINPUT9), .A3(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G99gat), .A2(G106gat), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(KEYINPUT6), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT6), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n532_), .A2(G99gat), .A3(G106gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n531_), .A2(new_n533_), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n528_), .A2(KEYINPUT9), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n529_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(KEYINPUT10), .B(G99gat), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT65), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n537_), .B1(new_n540_), .B2(G106gat), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT8), .ZN(new_n542_));
  OAI21_X1  g341(.A(KEYINPUT66), .B1(G99gat), .B2(G106gat), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT67), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT7), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT67), .ZN(new_n547_));
  OAI21_X1  g346(.A(KEYINPUT66), .B1(new_n547_), .B2(new_n545_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(G99gat), .A2(G106gat), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n546_), .A2(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n532_), .B1(G99gat), .B2(G106gat), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n530_), .A2(KEYINPUT6), .ZN(new_n553_));
  OAI21_X1  g352(.A(KEYINPUT69), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT69), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n531_), .A2(new_n533_), .A3(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n551_), .A2(new_n554_), .A3(new_n556_), .ZN(new_n557_));
  AND2_X1   g356(.A1(G85gat), .A2(G92gat), .ZN(new_n558_));
  NOR2_X1   g357(.A1(G85gat), .A2(G92gat), .ZN(new_n559_));
  OAI21_X1  g358(.A(KEYINPUT68), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT68), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n527_), .A2(new_n561_), .A3(new_n528_), .ZN(new_n562_));
  AND2_X1   g361(.A1(new_n560_), .A2(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n542_), .B1(new_n557_), .B2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n560_), .A2(new_n562_), .A3(new_n542_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n565_), .B1(new_n551_), .B2(new_n534_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n541_), .B1(new_n564_), .B2(new_n566_), .ZN(new_n567_));
  OR2_X1    g366(.A1(new_n567_), .A2(new_n481_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n482_), .A2(new_n567_), .A3(new_n484_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT73), .ZN(new_n570_));
  XNOR2_X1  g369(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G232gat), .A2(G233gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT35), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n568_), .A2(new_n569_), .A3(new_n570_), .A4(new_n576_), .ZN(new_n577_));
  AOI211_X1 g376(.A(new_n575_), .B(new_n574_), .C1(new_n569_), .C2(KEYINPUT73), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n574_), .A2(new_n575_), .ZN(new_n579_));
  AND3_X1   g378(.A1(new_n568_), .A2(new_n569_), .A3(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n577_), .B1(new_n578_), .B2(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G190gat), .B(G218gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT74), .ZN(new_n583_));
  XOR2_X1   g382(.A(G134gat), .B(G162gat), .Z(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT36), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n581_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n585_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n589_), .A2(KEYINPUT36), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n581_), .A2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n588_), .A2(KEYINPUT37), .A3(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n591_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT75), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n581_), .A2(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n587_), .B1(new_n581_), .B2(new_n594_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n593_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n524_), .B(new_n592_), .C1(new_n597_), .C2(KEYINPUT37), .ZN(new_n598_));
  NAND2_X1  g397(.A1(G230gat), .A2(G233gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT64), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n508_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n554_), .A2(new_n556_), .ZN(new_n603_));
  AOI22_X1  g402(.A1(new_n545_), .A2(new_n544_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n563_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n566_), .B1(new_n605_), .B2(KEYINPUT8), .ZN(new_n606_));
  INV_X1    g405(.A(new_n541_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n602_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  OAI211_X1 g407(.A(new_n508_), .B(new_n541_), .C1(new_n564_), .C2(new_n566_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n608_), .A2(KEYINPUT12), .A3(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT12), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n567_), .A2(new_n611_), .A3(new_n602_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n601_), .B1(new_n610_), .B2(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n600_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n614_));
  OR2_X1    g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G120gat), .B(G148gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT5), .ZN(new_n617_));
  XOR2_X1   g416(.A(G176gat), .B(G204gat), .Z(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n615_), .A2(new_n619_), .ZN(new_n620_));
  OR3_X1    g419(.A1(new_n613_), .A2(new_n614_), .A3(new_n619_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n620_), .A2(new_n621_), .A3(KEYINPUT70), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT70), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n615_), .A2(new_n623_), .A3(new_n619_), .ZN(new_n624_));
  AND3_X1   g423(.A1(new_n622_), .A2(KEYINPUT13), .A3(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(KEYINPUT13), .B1(new_n622_), .B2(new_n624_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n598_), .A2(new_n627_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n501_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n457_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n629_), .A2(new_n474_), .A3(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT38), .ZN(new_n632_));
  OAI211_X1 g431(.A(new_n524_), .B(new_n499_), .C1(new_n625_), .C2(new_n626_), .ZN(new_n633_));
  NOR3_X1   g432(.A1(new_n463_), .A2(new_n633_), .A3(new_n597_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n474_), .B1(new_n634_), .B2(new_n630_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT102), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n632_), .A2(new_n636_), .ZN(G1324gat));
  NAND2_X1  g436(.A1(new_n425_), .A2(new_n460_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n462_), .A2(new_n457_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n456_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n597_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n633_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n640_), .A2(new_n641_), .A3(new_n642_), .A4(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(G8gat), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(KEYINPUT39), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT39), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n644_), .A2(new_n647_), .A3(G8gat), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n629_), .A2(new_n475_), .A3(new_n641_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(KEYINPUT103), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT103), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n649_), .A2(new_n653_), .A3(new_n650_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n652_), .A2(new_n654_), .A3(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n655_), .B1(new_n652_), .B2(new_n654_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n656_), .A2(new_n657_), .ZN(G1325gat));
  INV_X1    g457(.A(G15gat), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n659_), .B1(new_n634_), .B2(new_n447_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT41), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n629_), .A2(new_n659_), .A3(new_n447_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1326gat));
  INV_X1    g462(.A(G22gat), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n423_), .B(KEYINPUT105), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n664_), .B1(new_n634_), .B2(new_n665_), .ZN(new_n666_));
  XOR2_X1   g465(.A(new_n666_), .B(KEYINPUT42), .Z(new_n667_));
  INV_X1    g466(.A(new_n629_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n665_), .A2(new_n664_), .ZN(new_n669_));
  XOR2_X1   g468(.A(new_n669_), .B(KEYINPUT106), .Z(new_n670_));
  OAI21_X1  g469(.A(new_n667_), .B1(new_n668_), .B2(new_n670_), .ZN(G1327gat));
  NOR2_X1   g470(.A1(new_n627_), .A2(new_n500_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(new_n523_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT43), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n592_), .B1(new_n597_), .B2(KEYINPUT37), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n640_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n676_), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n463_), .A2(KEYINPUT43), .A3(new_n678_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n674_), .B1(new_n677_), .B2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT44), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  OAI211_X1 g481(.A(new_n674_), .B(KEYINPUT44), .C1(new_n677_), .C2(new_n679_), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n682_), .A2(G29gat), .A3(new_n630_), .A4(new_n683_), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n627_), .A2(new_n642_), .A3(new_n524_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n501_), .A2(new_n685_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n686_), .A2(new_n457_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n684_), .B1(G29gat), .B2(new_n687_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT107), .ZN(G1328gat));
  NOR2_X1   g488(.A1(new_n456_), .A2(G36gat), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n501_), .A2(new_n685_), .A3(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT45), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n691_), .B(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n682_), .A2(new_n641_), .A3(new_n683_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n694_), .B2(G36gat), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT108), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT46), .ZN(new_n697_));
  AND3_X1   g496(.A1(new_n695_), .A2(new_n696_), .A3(new_n697_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n696_), .A2(new_n697_), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n695_), .A2(new_n699_), .A3(new_n700_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n698_), .A2(new_n701_), .ZN(G1329gat));
  INV_X1    g501(.A(G43gat), .ZN(new_n703_));
  INV_X1    g502(.A(new_n447_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n703_), .B1(new_n686_), .B2(new_n704_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT109), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n682_), .A2(G43gat), .A3(new_n447_), .A4(new_n683_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g508(.A(new_n686_), .ZN(new_n710_));
  AOI21_X1  g509(.A(G50gat), .B1(new_n710_), .B2(new_n665_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n682_), .A2(new_n683_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n459_), .A2(G50gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n711_), .B1(new_n712_), .B2(new_n713_), .ZN(G1331gat));
  NOR2_X1   g513(.A1(new_n463_), .A2(new_n597_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n627_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n716_), .A2(new_n499_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n715_), .A2(new_n524_), .A3(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(G57gat), .B1(new_n718_), .B2(new_n457_), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n463_), .A2(new_n716_), .A3(new_n499_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n720_), .A2(new_n524_), .A3(new_n678_), .ZN(new_n721_));
  OR2_X1    g520(.A1(new_n457_), .A2(G57gat), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n719_), .B1(new_n721_), .B2(new_n722_), .ZN(G1332gat));
  OAI21_X1  g522(.A(G64gat), .B1(new_n718_), .B2(new_n456_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT48), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n456_), .A2(G64gat), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n725_), .B1(new_n721_), .B2(new_n726_), .ZN(G1333gat));
  OAI21_X1  g526(.A(G71gat), .B1(new_n718_), .B2(new_n704_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT49), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n704_), .A2(G71gat), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n729_), .B1(new_n721_), .B2(new_n730_), .ZN(G1334gat));
  NAND4_X1  g530(.A1(new_n715_), .A2(new_n524_), .A3(new_n717_), .A4(new_n665_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(G78gat), .ZN(new_n733_));
  XNOR2_X1  g532(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n733_), .B(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(G78gat), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n665_), .A2(new_n736_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n735_), .B1(new_n721_), .B2(new_n737_), .ZN(G1335gat));
  AND3_X1   g537(.A1(new_n720_), .A2(new_n597_), .A3(new_n523_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n739_), .A2(new_n525_), .A3(new_n630_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n677_), .A2(new_n679_), .ZN(new_n741_));
  NOR4_X1   g540(.A1(new_n741_), .A2(new_n524_), .A3(new_n499_), .A4(new_n716_), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n742_), .A2(new_n630_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n740_), .B1(new_n743_), .B2(new_n525_), .ZN(G1336gat));
  NAND3_X1  g543(.A1(new_n739_), .A2(new_n526_), .A3(new_n641_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n742_), .A2(new_n641_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n745_), .B1(new_n746_), .B2(new_n526_), .ZN(G1337gat));
  NOR2_X1   g546(.A1(new_n704_), .A2(new_n540_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n739_), .A2(new_n748_), .ZN(new_n749_));
  NOR3_X1   g548(.A1(new_n716_), .A2(new_n524_), .A3(new_n499_), .ZN(new_n750_));
  OAI211_X1 g549(.A(new_n750_), .B(new_n447_), .C1(new_n677_), .C2(new_n679_), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n751_), .A2(KEYINPUT111), .A3(G99gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(KEYINPUT111), .B1(new_n751_), .B2(G99gat), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n749_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g554(.A(G106gat), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n739_), .A2(new_n756_), .A3(new_n459_), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n750_), .B(new_n459_), .C1(new_n677_), .C2(new_n679_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT52), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n758_), .A2(new_n759_), .A3(G106gat), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n758_), .B2(G106gat), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n757_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g562(.A(KEYINPUT112), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n764_), .B1(new_n499_), .B2(new_n621_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n499_), .A2(new_n764_), .A3(new_n621_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT113), .ZN(new_n769_));
  OAI21_X1  g568(.A(KEYINPUT115), .B1(new_n613_), .B2(new_n769_), .ZN(new_n770_));
  OAI21_X1  g569(.A(KEYINPUT55), .B1(new_n613_), .B2(KEYINPUT115), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n610_), .A2(new_n612_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT114), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT114), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n610_), .A2(new_n775_), .A3(new_n612_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n774_), .A2(new_n601_), .A3(new_n776_), .ZN(new_n777_));
  OAI211_X1 g576(.A(KEYINPUT115), .B(KEYINPUT55), .C1(new_n613_), .C2(new_n769_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n619_), .B1(new_n772_), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT56), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  OAI211_X1 g581(.A(KEYINPUT56), .B(new_n619_), .C1(new_n772_), .C2(new_n779_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n768_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n498_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n489_), .A2(new_n464_), .A3(new_n490_), .ZN(new_n786_));
  AOI21_X1  g585(.A(KEYINPUT116), .B1(new_n786_), .B2(new_n496_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n464_), .B1(new_n472_), .B2(new_n479_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n787_), .B1(new_n486_), .B2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n786_), .A2(KEYINPUT116), .A3(new_n496_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n785_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n791_), .A2(new_n622_), .A3(new_n624_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n642_), .B1(new_n784_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT57), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n767_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n797_), .A2(new_n765_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n783_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n770_), .A2(new_n771_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n800_), .A2(new_n778_), .A3(new_n777_), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT56), .B1(new_n801_), .B2(new_n619_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n798_), .B1(new_n799_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n792_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n804_), .A2(KEYINPUT57), .A3(new_n642_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n791_), .A2(new_n621_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n806_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n807_));
  OAI211_X1 g606(.A(KEYINPUT117), .B(new_n676_), .C1(new_n807_), .C2(KEYINPUT58), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(KEYINPUT58), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n806_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n811_), .B1(new_n799_), .B2(new_n802_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT58), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(KEYINPUT117), .B1(new_n814_), .B2(new_n676_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n796_), .B(new_n805_), .C1(new_n810_), .C2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n523_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n818_), .B1(new_n628_), .B2(new_n500_), .ZN(new_n819_));
  NOR4_X1   g618(.A1(new_n598_), .A2(new_n627_), .A3(KEYINPUT54), .A4(new_n499_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n457_), .B1(new_n817_), .B2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n823_), .A2(KEYINPUT59), .A3(new_n462_), .ZN(new_n824_));
  AOI21_X1  g623(.A(KEYINPUT57), .B1(new_n804_), .B2(new_n642_), .ZN(new_n825_));
  AOI211_X1 g624(.A(new_n795_), .B(new_n597_), .C1(new_n803_), .C2(new_n792_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n676_), .B1(new_n807_), .B2(KEYINPUT58), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT117), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n830_), .A2(new_n809_), .A3(new_n808_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n524_), .B1(new_n827_), .B2(new_n831_), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n630_), .B(new_n462_), .C1(new_n832_), .C2(new_n821_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT59), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n824_), .A2(new_n835_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n500_), .A2(KEYINPUT118), .ZN(new_n837_));
  MUX2_X1   g636(.A(KEYINPUT118), .B(new_n837_), .S(G113gat), .Z(new_n838_));
  INV_X1    g637(.A(G113gat), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n823_), .A2(new_n462_), .A3(new_n499_), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n836_), .A2(new_n838_), .B1(new_n839_), .B2(new_n840_), .ZN(G1340gat));
  AOI21_X1  g640(.A(new_n716_), .B1(new_n824_), .B2(new_n835_), .ZN(new_n842_));
  INV_X1    g641(.A(G120gat), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n843_), .B1(new_n716_), .B2(KEYINPUT60), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n843_), .A2(KEYINPUT60), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n844_), .B1(KEYINPUT119), .B2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n846_), .B1(KEYINPUT119), .B2(new_n844_), .ZN(new_n847_));
  OAI22_X1  g646(.A1(new_n842_), .A2(new_n843_), .B1(new_n833_), .B2(new_n847_), .ZN(G1341gat));
  AOI21_X1  g647(.A(new_n523_), .B1(new_n824_), .B2(new_n835_), .ZN(new_n849_));
  INV_X1    g648(.A(G127gat), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n524_), .A2(new_n850_), .ZN(new_n851_));
  OAI22_X1  g650(.A1(new_n849_), .A2(new_n850_), .B1(new_n833_), .B2(new_n851_), .ZN(G1342gat));
  AOI21_X1  g651(.A(new_n678_), .B1(new_n824_), .B2(new_n835_), .ZN(new_n853_));
  INV_X1    g652(.A(G134gat), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n597_), .A2(new_n854_), .ZN(new_n855_));
  OAI22_X1  g654(.A1(new_n853_), .A2(new_n854_), .B1(new_n833_), .B2(new_n855_), .ZN(G1343gat));
  NAND2_X1  g655(.A1(new_n704_), .A2(new_n459_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n857_), .A2(new_n641_), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n630_), .B(new_n858_), .C1(new_n832_), .C2(new_n821_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n859_), .A2(new_n500_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(new_n207_), .ZN(G1344gat));
  NOR2_X1   g660(.A1(new_n859_), .A2(new_n716_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(KEYINPUT120), .B(G148gat), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n862_), .B(new_n863_), .ZN(G1345gat));
  OAI21_X1  g663(.A(KEYINPUT121), .B1(new_n859_), .B2(new_n523_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT121), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n823_), .A2(new_n866_), .A3(new_n524_), .A4(new_n858_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(KEYINPUT61), .B(G155gat), .ZN(new_n868_));
  AND3_X1   g667(.A1(new_n865_), .A2(new_n867_), .A3(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n868_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1346gat));
  INV_X1    g670(.A(G162gat), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n859_), .A2(new_n872_), .A3(new_n678_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n859_), .B2(new_n642_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT122), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  OAI211_X1 g675(.A(KEYINPUT122), .B(new_n872_), .C1(new_n859_), .C2(new_n642_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n873_), .B1(new_n876_), .B2(new_n877_), .ZN(G1347gat));
  AOI21_X1  g677(.A(new_n821_), .B1(new_n816_), .B2(new_n523_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n641_), .A2(new_n457_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n881_), .A2(new_n704_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n883_), .A2(new_n665_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n880_), .A2(new_n499_), .A3(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT62), .ZN(new_n886_));
  AND3_X1   g685(.A1(new_n885_), .A2(new_n886_), .A3(G169gat), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n886_), .B1(new_n885_), .B2(G169gat), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n880_), .A2(new_n884_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n499_), .A2(new_n299_), .ZN(new_n890_));
  XOR2_X1   g689(.A(new_n890_), .B(KEYINPUT123), .Z(new_n891_));
  OAI22_X1  g690(.A1(new_n887_), .A2(new_n888_), .B1(new_n889_), .B2(new_n891_), .ZN(G1348gat));
  NAND3_X1  g691(.A1(new_n880_), .A2(new_n627_), .A3(new_n884_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n879_), .A2(new_n459_), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n883_), .A2(new_n716_), .A3(new_n300_), .ZN(new_n895_));
  AOI22_X1  g694(.A1(new_n893_), .A2(new_n300_), .B1(new_n894_), .B2(new_n895_), .ZN(G1349gat));
  NOR3_X1   g695(.A1(new_n889_), .A2(new_n284_), .A3(new_n523_), .ZN(new_n897_));
  NOR4_X1   g696(.A1(new_n879_), .A2(new_n459_), .A3(new_n523_), .A4(new_n883_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT124), .ZN(new_n899_));
  OR2_X1    g698(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  AOI21_X1  g699(.A(G183gat), .B1(new_n898_), .B2(new_n899_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n897_), .B1(new_n900_), .B2(new_n901_), .ZN(G1350gat));
  OAI21_X1  g701(.A(G190gat), .B1(new_n889_), .B2(new_n678_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n597_), .A2(new_n329_), .A3(new_n327_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n903_), .B1(new_n889_), .B2(new_n904_), .ZN(G1351gat));
  NOR2_X1   g704(.A1(new_n857_), .A2(new_n881_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n906_), .ZN(new_n907_));
  OAI21_X1  g706(.A(KEYINPUT125), .B1(new_n879_), .B2(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT125), .ZN(new_n909_));
  OAI211_X1 g708(.A(new_n909_), .B(new_n906_), .C1(new_n832_), .C2(new_n821_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n500_), .B1(new_n908_), .B2(new_n910_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(new_n269_), .ZN(G1352gat));
  AOI21_X1  g711(.A(new_n716_), .B1(new_n908_), .B2(new_n910_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n913_), .B(new_n914_), .ZN(G1353gat));
  AOI21_X1  g714(.A(new_n523_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n916_));
  INV_X1    g715(.A(new_n916_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n917_), .B1(new_n908_), .B2(new_n910_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(KEYINPUT127), .ZN(new_n920_));
  INV_X1    g719(.A(new_n920_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n918_), .B(new_n921_), .ZN(G1354gat));
  NAND2_X1  g721(.A1(new_n908_), .A2(new_n910_), .ZN(new_n923_));
  INV_X1    g722(.A(G218gat), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n923_), .A2(new_n924_), .A3(new_n597_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n678_), .B1(new_n908_), .B2(new_n910_), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n925_), .B1(new_n924_), .B2(new_n926_), .ZN(G1355gat));
endmodule


