//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 0 1 1 1 0 0 1 0 1 0 0 0 0 0 0 1 0 0 1 0 0 0 0 1 1 0 0 1 0 1 0 0 1 0 1 0 0 1 0 1 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n804_, new_n805_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n873_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n951_, new_n952_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n959_, new_n961_,
    new_n962_, new_n963_, new_n965_, new_n966_, new_n967_, new_n968_,
    new_n969_, new_n970_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n982_,
    new_n983_, new_n985_, new_n986_, new_n987_, new_n989_, new_n990_,
    new_n991_, new_n992_, new_n993_, new_n994_, new_n995_, new_n996_,
    new_n998_, new_n999_, new_n1000_, new_n1002_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1009_, new_n1010_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(new_n202_), .B(KEYINPUT64), .Z(new_n203_));
  XOR2_X1   g002(.A(G71gat), .B(G78gat), .Z(new_n204_));
  XNOR2_X1  g003(.A(G57gat), .B(G64gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(new_n204_), .B1(KEYINPUT11), .B2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(KEYINPUT11), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  XOR2_X1   g008(.A(G85gat), .B(G92gat), .Z(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT68), .ZN(new_n213_));
  AOI21_X1  g012(.A(KEYINPUT67), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT7), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n212_), .A2(KEYINPUT67), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT7), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n216_), .B1(new_n214_), .B2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G99gat), .A2(G106gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(KEYINPUT6), .ZN(new_n221_));
  AOI211_X1 g020(.A(KEYINPUT8), .B(new_n211_), .C1(new_n219_), .C2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  XOR2_X1   g022(.A(KEYINPUT69), .B(KEYINPUT6), .Z(new_n224_));
  INV_X1    g023(.A(new_n220_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT69), .B(KEYINPUT6), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(new_n220_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n226_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT70), .ZN(new_n230_));
  OR2_X1    g029(.A1(new_n218_), .A2(new_n214_), .ZN(new_n231_));
  AOI22_X1  g030(.A1(new_n229_), .A2(new_n230_), .B1(new_n231_), .B2(new_n216_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n226_), .A2(KEYINPUT70), .A3(new_n228_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n211_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT8), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n223_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  XOR2_X1   g035(.A(KEYINPUT10), .B(G99gat), .Z(new_n237_));
  INV_X1    g036(.A(G106gat), .ZN(new_n238_));
  INV_X1    g037(.A(G85gat), .ZN(new_n239_));
  INV_X1    g038(.A(G92gat), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT65), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n242_), .A2(KEYINPUT9), .ZN(new_n243_));
  AOI22_X1  g042(.A1(new_n237_), .A2(new_n238_), .B1(new_n241_), .B2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n243_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n242_), .A2(KEYINPUT9), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n210_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n244_), .A2(new_n221_), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT66), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n209_), .B1(new_n236_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n228_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n227_), .A2(new_n220_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n230_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n254_), .A2(new_n233_), .A3(new_n219_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n235_), .B1(new_n255_), .B2(new_n210_), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n250_), .B(new_n209_), .C1(new_n256_), .C2(new_n222_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT12), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n251_), .A2(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n250_), .B1(new_n256_), .B2(new_n222_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT12), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n260_), .A2(new_n261_), .A3(new_n208_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n203_), .B1(new_n259_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT71), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n260_), .A2(new_n208_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n203_), .B1(new_n266_), .B2(new_n257_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n264_), .A2(new_n265_), .A3(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n203_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n266_), .A2(KEYINPUT12), .A3(new_n257_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n270_), .B1(new_n271_), .B2(new_n262_), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT71), .B1(new_n272_), .B2(new_n267_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G120gat), .B(G148gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(G204gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT5), .B(G176gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  XOR2_X1   g076(.A(new_n277_), .B(KEYINPUT72), .Z(new_n278_));
  NAND3_X1  g077(.A1(new_n269_), .A2(new_n273_), .A3(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n264_), .A2(new_n268_), .A3(new_n277_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT13), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n279_), .A2(KEYINPUT13), .A3(new_n280_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(KEYINPUT73), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G169gat), .A2(G176gat), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT86), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(G183gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(KEYINPUT83), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT83), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(G183gat), .ZN(new_n293_));
  INV_X1    g092(.A(G190gat), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n291_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G183gat), .A2(G190gat), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT23), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n289_), .B1(new_n295_), .B2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(G169gat), .ZN(new_n302_));
  AOI21_X1  g101(.A(G176gat), .B1(new_n302_), .B2(KEYINPUT22), .ZN(new_n303_));
  OR2_X1    g102(.A1(KEYINPUT87), .A2(KEYINPUT22), .ZN(new_n304_));
  NAND2_X1  g103(.A1(KEYINPUT87), .A2(KEYINPUT22), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n302_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT88), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n303_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n304_), .A2(new_n305_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n309_), .A2(new_n307_), .A3(G169gat), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n301_), .B1(new_n308_), .B2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n294_), .A2(KEYINPUT26), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT84), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n294_), .A2(KEYINPUT84), .A3(KEYINPUT26), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT26), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(G190gat), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT85), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n318_), .A2(KEYINPUT85), .A3(G190gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT25), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n324_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n326_));
  OAI211_X1 g125(.A(new_n317_), .B(new_n323_), .C1(new_n325_), .C2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n287_), .B(KEYINPUT86), .ZN(new_n328_));
  INV_X1    g127(.A(G176gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n302_), .A2(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n328_), .A2(KEYINPUT24), .A3(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n298_), .A2(new_n299_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT24), .ZN(new_n333_));
  INV_X1    g132(.A(new_n330_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n332_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n327_), .A2(new_n331_), .A3(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n312_), .A2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT30), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT89), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT31), .ZN(new_n340_));
  OR2_X1    g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n339_), .A2(new_n340_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  XOR2_X1   g142(.A(G71gat), .B(G99gat), .Z(new_n344_));
  NAND2_X1  g143(.A1(G227gat), .A2(G233gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  XOR2_X1   g145(.A(G15gat), .B(G43gat), .Z(new_n347_));
  XOR2_X1   g146(.A(new_n346_), .B(new_n347_), .Z(new_n348_));
  XOR2_X1   g147(.A(G127gat), .B(G134gat), .Z(new_n349_));
  XOR2_X1   g148(.A(G113gat), .B(G120gat), .Z(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n348_), .B(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n343_), .A2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n341_), .A2(new_n342_), .A3(new_n353_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT101), .B(KEYINPUT0), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G1gat), .B(G29gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G57gat), .B(G85gat), .ZN(new_n361_));
  XOR2_X1   g160(.A(new_n360_), .B(new_n361_), .Z(new_n362_));
  NAND2_X1  g161(.A1(G155gat), .A2(G162gat), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT90), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT1), .ZN(new_n366_));
  NAND3_X1  g165(.A1(KEYINPUT90), .A2(G155gat), .A3(G162gat), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n365_), .A2(new_n366_), .A3(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT91), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT91), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n365_), .A2(new_n370_), .A3(new_n366_), .A4(new_n367_), .ZN(new_n371_));
  OR2_X1    g170(.A1(G155gat), .A2(G162gat), .ZN(new_n372_));
  INV_X1    g171(.A(new_n367_), .ZN(new_n373_));
  AOI21_X1  g172(.A(KEYINPUT90), .B1(G155gat), .B2(G162gat), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT1), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n369_), .A2(new_n371_), .A3(new_n372_), .A4(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G141gat), .A2(G148gat), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(G141gat), .A2(G148gat), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n376_), .A2(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n372_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n379_), .B(KEYINPUT3), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n377_), .B(KEYINPUT2), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n382_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n381_), .A2(new_n386_), .ZN(new_n387_));
  XOR2_X1   g186(.A(KEYINPUT100), .B(KEYINPUT4), .Z(new_n388_));
  NAND3_X1  g187(.A1(new_n387_), .A2(new_n352_), .A3(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G225gat), .A2(G233gat), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n387_), .A2(new_n352_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n385_), .B1(new_n376_), .B2(new_n380_), .ZN(new_n394_));
  AOI21_X1  g193(.A(KEYINPUT99), .B1(new_n394_), .B2(new_n351_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n387_), .A2(KEYINPUT99), .A3(new_n352_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n392_), .B1(new_n398_), .B2(KEYINPUT4), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n391_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n362_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n398_), .A2(new_n390_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n362_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT4), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n404_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n405_));
  OAI211_X1 g204(.A(new_n402_), .B(new_n403_), .C1(new_n405_), .C2(new_n392_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n401_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT29), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n394_), .A2(new_n408_), .ZN(new_n409_));
  XOR2_X1   g208(.A(G211gat), .B(G218gat), .Z(new_n410_));
  INV_X1    g209(.A(G204gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(G197gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT92), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT92), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n414_), .A2(new_n411_), .A3(G197gat), .ZN(new_n415_));
  INV_X1    g214(.A(G197gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(G204gat), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n413_), .A2(new_n415_), .A3(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n410_), .B1(new_n418_), .B2(KEYINPUT21), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT93), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n412_), .A2(new_n417_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n420_), .B1(new_n421_), .B2(KEYINPUT21), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT21), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n412_), .A2(new_n417_), .A3(KEYINPUT93), .A4(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n419_), .A2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n410_), .A2(KEYINPUT21), .A3(new_n421_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n428_), .B1(new_n394_), .B2(new_n408_), .ZN(new_n429_));
  INV_X1    g228(.A(G228gat), .ZN(new_n430_));
  INV_X1    g229(.A(G233gat), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n429_), .A2(new_n432_), .ZN(new_n433_));
  OAI221_X1 g232(.A(new_n428_), .B1(new_n430_), .B2(new_n431_), .C1(new_n394_), .C2(new_n408_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n409_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n433_), .A2(new_n434_), .A3(new_n409_), .ZN(new_n437_));
  XOR2_X1   g236(.A(G22gat), .B(G50gat), .Z(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(KEYINPUT28), .ZN(new_n439_));
  XOR2_X1   g238(.A(G78gat), .B(G106gat), .Z(new_n440_));
  XOR2_X1   g239(.A(new_n439_), .B(new_n440_), .Z(new_n441_));
  NAND3_X1  g240(.A1(new_n436_), .A2(new_n437_), .A3(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n441_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n437_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n443_), .B1(new_n444_), .B2(new_n435_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n442_), .A2(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G8gat), .B(G36gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n447_), .B(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G64gat), .B(G92gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n449_), .B(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G226gat), .A2(G233gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(KEYINPUT19), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT20), .ZN(new_n456_));
  AND2_X1   g255(.A1(KEYINPUT94), .A2(KEYINPUT24), .ZN(new_n457_));
  NOR2_X1   g256(.A1(KEYINPUT94), .A2(KEYINPUT24), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n332_), .B1(new_n334_), .B2(new_n459_), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n330_), .B(new_n287_), .C1(new_n457_), .C2(new_n458_), .ZN(new_n461_));
  AND2_X1   g260(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n313_), .B(new_n319_), .C1(new_n462_), .C2(new_n326_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n461_), .A2(new_n463_), .A3(KEYINPUT95), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(KEYINPUT95), .B1(new_n461_), .B2(new_n463_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n460_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(KEYINPUT22), .B(G169gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(new_n329_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(G183gat), .A2(G190gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n296_), .A2(KEYINPUT23), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n297_), .A2(G183gat), .A3(G190gat), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n470_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n473_), .A2(KEYINPUT96), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT96), .ZN(new_n475_));
  AOI211_X1 g274(.A(new_n475_), .B(new_n470_), .C1(new_n471_), .C2(new_n472_), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n328_), .B(new_n469_), .C1(new_n474_), .C2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n467_), .A2(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n456_), .B1(new_n478_), .B2(new_n428_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n427_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n480_), .B1(new_n419_), .B2(new_n425_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n481_), .A2(new_n312_), .A3(new_n336_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n455_), .B1(new_n479_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n337_), .A2(new_n428_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n467_), .A2(new_n481_), .A3(new_n477_), .ZN(new_n485_));
  AND4_X1   g284(.A1(KEYINPUT20), .A2(new_n484_), .A3(new_n455_), .A4(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n452_), .B1(new_n483_), .B2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n460_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n466_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n488_), .B1(new_n489_), .B2(new_n464_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n469_), .A2(new_n328_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n474_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n476_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n491_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n428_), .B1(new_n490_), .B2(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n495_), .A2(KEYINPUT20), .A3(new_n482_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(new_n454_), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n484_), .A2(new_n485_), .A3(KEYINPUT20), .A4(new_n455_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n497_), .A2(new_n451_), .A3(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n487_), .A2(KEYINPUT98), .A3(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT27), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT98), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n497_), .A2(new_n502_), .A3(new_n451_), .A4(new_n498_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n500_), .A2(new_n501_), .A3(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n484_), .A2(KEYINPUT20), .A3(new_n485_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(new_n454_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n479_), .A2(new_n455_), .A3(new_n482_), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  OAI211_X1 g307(.A(KEYINPUT27), .B(new_n499_), .C1(new_n508_), .C2(new_n451_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n504_), .A2(new_n509_), .ZN(new_n510_));
  NOR4_X1   g309(.A1(new_n357_), .A2(new_n407_), .A3(new_n446_), .A4(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n446_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n451_), .A2(KEYINPUT32), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n513_), .B1(new_n483_), .B2(new_n486_), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n506_), .A2(new_n507_), .A3(KEYINPUT32), .A4(new_n451_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n407_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(KEYINPUT104), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT104), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n407_), .A2(new_n519_), .A3(new_n516_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n403_), .B1(new_n398_), .B2(new_n391_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n398_), .A2(KEYINPUT4), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n389_), .A2(new_n390_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(KEYINPUT102), .B1(new_n523_), .B2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT102), .ZN(new_n527_));
  NOR3_X1   g326(.A1(new_n405_), .A2(new_n527_), .A3(new_n524_), .ZN(new_n528_));
  OAI211_X1 g327(.A(KEYINPUT103), .B(new_n522_), .C1(new_n526_), .C2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT33), .ZN(new_n530_));
  INV_X1    g329(.A(new_n392_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n400_), .B1(new_n523_), .B2(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n530_), .B1(new_n532_), .B2(new_n403_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n406_), .A2(KEYINPUT33), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n529_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n500_), .A2(new_n503_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n398_), .A2(new_n391_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(new_n362_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n523_), .A2(KEYINPUT102), .A3(new_n525_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n527_), .B1(new_n405_), .B2(new_n524_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n538_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n536_), .B1(new_n541_), .B2(KEYINPUT103), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n535_), .A2(new_n542_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n512_), .B1(new_n521_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT105), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n446_), .A2(new_n401_), .A3(new_n406_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n545_), .B1(new_n510_), .B2(new_n546_), .ZN(new_n547_));
  AND3_X1   g346(.A1(new_n446_), .A2(new_n401_), .A3(new_n406_), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n548_), .A2(KEYINPUT105), .A3(new_n504_), .A4(new_n509_), .ZN(new_n549_));
  AND2_X1   g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n544_), .A2(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n511_), .B1(new_n551_), .B2(new_n357_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT37), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT74), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G232gat), .A2(G233gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT34), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT35), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G29gat), .B(G50gat), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  XOR2_X1   g360(.A(G36gat), .B(G43gat), .Z(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G36gat), .B(G43gat), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n560_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT15), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n260_), .A2(new_n567_), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n250_), .B(new_n566_), .C1(new_n256_), .C2(new_n222_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n557_), .A2(new_n558_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n559_), .B1(new_n568_), .B2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n260_), .A2(new_n567_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n559_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n573_), .A2(new_n574_), .A3(new_n570_), .A4(new_n569_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n554_), .B1(new_n572_), .B2(new_n575_), .ZN(new_n576_));
  XOR2_X1   g375(.A(G190gat), .B(G218gat), .Z(new_n577_));
  XNOR2_X1  g376(.A(G134gat), .B(G162gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(KEYINPUT36), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n581_), .B1(new_n572_), .B2(new_n575_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n580_), .A2(KEYINPUT36), .ZN(new_n583_));
  NOR3_X1   g382(.A1(new_n576_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n583_), .ZN(new_n585_));
  AOI221_X4 g384(.A(new_n554_), .B1(new_n585_), .B2(new_n581_), .C1(new_n572_), .C2(new_n575_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n553_), .B1(new_n584_), .B2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n576_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n572_), .A2(new_n575_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n581_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n588_), .A2(new_n591_), .A3(new_n585_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n586_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n592_), .A2(new_n593_), .A3(KEYINPUT37), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n587_), .A2(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G113gat), .B(G141gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(G169gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(new_n416_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(G229gat), .A2(G233gat), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(G8gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(KEYINPUT75), .B(G1gat), .ZN(new_n602_));
  OAI21_X1  g401(.A(KEYINPUT14), .B1(new_n602_), .B2(new_n601_), .ZN(new_n603_));
  INV_X1    g402(.A(G1gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G15gat), .B(G22gat), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n603_), .A2(new_n604_), .A3(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n604_), .B1(new_n603_), .B2(new_n605_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n601_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n603_), .A2(new_n605_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(G1gat), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n611_), .A2(G8gat), .A3(new_n606_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n609_), .A2(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n600_), .B1(new_n613_), .B2(new_n567_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT78), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT77), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n566_), .A2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n563_), .A2(KEYINPUT77), .A3(new_n565_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  AOI211_X1 g418(.A(new_n615_), .B(new_n619_), .C1(new_n609_), .C2(new_n612_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n609_), .A2(new_n612_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n619_), .ZN(new_n622_));
  AOI21_X1  g421(.A(KEYINPUT78), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n614_), .B1(new_n620_), .B2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT79), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n613_), .A2(new_n619_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n627_), .B1(new_n620_), .B2(new_n623_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(new_n600_), .ZN(new_n629_));
  OAI211_X1 g428(.A(new_n614_), .B(KEYINPUT79), .C1(new_n623_), .C2(new_n620_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n626_), .A2(new_n629_), .A3(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n598_), .B1(new_n631_), .B2(KEYINPUT80), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT80), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n626_), .A2(new_n629_), .A3(new_n633_), .A4(new_n630_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(KEYINPUT81), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT81), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n632_), .A2(new_n637_), .A3(new_n634_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n626_), .A2(new_n629_), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n639_), .A2(KEYINPUT82), .A3(new_n630_), .A4(new_n598_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT82), .ZN(new_n641_));
  INV_X1    g440(.A(new_n598_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n641_), .B1(new_n631_), .B2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n640_), .A2(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n636_), .A2(new_n638_), .A3(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(G231gat), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n613_), .B1(new_n646_), .B2(new_n431_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n621_), .A2(G231gat), .A3(G233gat), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(new_n209_), .ZN(new_n650_));
  XOR2_X1   g449(.A(KEYINPUT76), .B(KEYINPUT16), .Z(new_n651_));
  XNOR2_X1  g450(.A(G127gat), .B(G155gat), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n651_), .B(new_n652_), .ZN(new_n653_));
  XOR2_X1   g452(.A(G183gat), .B(G211gat), .Z(new_n654_));
  XNOR2_X1  g453(.A(new_n653_), .B(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT17), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n650_), .A2(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n655_), .B(KEYINPUT17), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n659_), .B1(new_n650_), .B2(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n595_), .A2(new_n645_), .A3(new_n661_), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n286_), .A2(new_n552_), .A3(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n407_), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n664_), .A2(KEYINPUT106), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(KEYINPUT106), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n663_), .A2(new_n602_), .A3(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT38), .ZN(new_n669_));
  AOI221_X4 g468(.A(KEYINPUT104), .B1(new_n514_), .B2(new_n515_), .C1(new_n401_), .C2(new_n406_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n519_), .B1(new_n407_), .B2(new_n516_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n522_), .B1(new_n526_), .B2(new_n528_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT103), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n532_), .A2(new_n530_), .A3(new_n403_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n406_), .A2(KEYINPUT33), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n675_), .A2(new_n678_), .A3(new_n536_), .A4(new_n529_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n446_), .B1(new_n672_), .B2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n547_), .A2(new_n549_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n357_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n511_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n584_), .A2(new_n586_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT107), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n645_), .A2(new_n661_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n687_), .B1(new_n688_), .B2(new_n285_), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n279_), .A2(KEYINPUT13), .A3(new_n280_), .ZN(new_n690_));
  AOI21_X1  g489(.A(KEYINPUT13), .B1(new_n279_), .B2(new_n280_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n692_), .A2(KEYINPUT107), .A3(new_n645_), .A4(new_n661_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n689_), .A2(new_n693_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n686_), .A2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  OAI21_X1  g495(.A(G1gat), .B1(new_n696_), .B2(new_n664_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n669_), .A2(new_n697_), .ZN(G1324gat));
  INV_X1    g497(.A(KEYINPUT40), .ZN(new_n699_));
  INV_X1    g498(.A(new_n510_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n700_), .A2(G8gat), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n663_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n686_), .A2(new_n694_), .A3(new_n700_), .ZN(new_n704_));
  OAI21_X1  g503(.A(KEYINPUT39), .B1(new_n704_), .B2(new_n601_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n686_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n694_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n706_), .A2(new_n707_), .A3(new_n510_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT39), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n708_), .A2(new_n709_), .A3(G8gat), .ZN(new_n710_));
  AOI211_X1 g509(.A(KEYINPUT108), .B(new_n703_), .C1(new_n705_), .C2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n705_), .A2(new_n710_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n713_), .B2(new_n702_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n699_), .B1(new_n711_), .B2(new_n714_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n704_), .A2(KEYINPUT39), .A3(new_n601_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n709_), .B1(new_n708_), .B2(G8gat), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n702_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(KEYINPUT108), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n713_), .A2(new_n712_), .A3(new_n702_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n719_), .A2(KEYINPUT40), .A3(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n715_), .A2(new_n721_), .ZN(G1325gat));
  INV_X1    g521(.A(KEYINPUT109), .ZN(new_n723_));
  INV_X1    g522(.A(new_n357_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n695_), .A2(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n723_), .B1(new_n725_), .B2(G15gat), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n686_), .A2(new_n694_), .A3(new_n357_), .ZN(new_n727_));
  INV_X1    g526(.A(G15gat), .ZN(new_n728_));
  NOR3_X1   g527(.A1(new_n727_), .A2(KEYINPUT109), .A3(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(KEYINPUT110), .B1(new_n726_), .B2(new_n729_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n725_), .A2(new_n723_), .A3(G15gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(KEYINPUT109), .B1(new_n727_), .B2(new_n728_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT110), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n731_), .A2(new_n732_), .A3(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n730_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT41), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n663_), .A2(new_n728_), .A3(new_n724_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n730_), .A2(KEYINPUT41), .A3(new_n734_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n737_), .A2(new_n738_), .A3(new_n739_), .ZN(G1326gat));
  INV_X1    g539(.A(G22gat), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n663_), .A2(new_n741_), .A3(new_n446_), .ZN(new_n742_));
  OAI21_X1  g541(.A(G22gat), .B1(new_n696_), .B2(new_n512_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(KEYINPUT111), .B(KEYINPUT42), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n743_), .A2(new_n744_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n742_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT112), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  OAI211_X1 g548(.A(KEYINPUT112), .B(new_n742_), .C1(new_n745_), .C2(new_n746_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1327gat));
  INV_X1    g550(.A(new_n661_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n692_), .A2(new_n645_), .A3(new_n752_), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n552_), .A2(new_n685_), .A3(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(G29gat), .B1(new_n754_), .B2(new_n407_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(KEYINPUT113), .B(KEYINPUT43), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT114), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n595_), .A2(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(KEYINPUT114), .B1(new_n587_), .B2(new_n594_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n756_), .B1(new_n552_), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT115), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT43), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n587_), .A2(new_n763_), .A3(new_n594_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n762_), .B1(new_n684_), .B2(new_n765_), .ZN(new_n766_));
  AOI211_X1 g565(.A(KEYINPUT115), .B(new_n764_), .C1(new_n682_), .C2(new_n683_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n761_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n753_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n768_), .A2(KEYINPUT44), .A3(new_n769_), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n770_), .A2(G29gat), .A3(new_n667_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n768_), .A2(new_n769_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT44), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n755_), .B1(new_n771_), .B2(new_n774_), .ZN(G1328gat));
  INV_X1    g574(.A(KEYINPUT46), .ZN(new_n776_));
  INV_X1    g575(.A(G36gat), .ZN(new_n777_));
  OAI21_X1  g576(.A(KEYINPUT115), .B1(new_n552_), .B2(new_n764_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n684_), .A2(new_n762_), .A3(new_n765_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n753_), .B1(new_n780_), .B2(new_n761_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n700_), .B1(new_n781_), .B2(KEYINPUT44), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n777_), .B1(new_n782_), .B2(new_n774_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n754_), .A2(new_n777_), .A3(new_n510_), .ZN(new_n784_));
  OR2_X1    g583(.A1(new_n784_), .A2(KEYINPUT45), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(KEYINPUT45), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n776_), .B1(new_n783_), .B2(new_n788_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n781_), .A2(KEYINPUT44), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n770_), .A2(new_n510_), .ZN(new_n791_));
  OAI21_X1  g590(.A(G36gat), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n792_), .A2(new_n787_), .A3(KEYINPUT46), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n789_), .A2(new_n793_), .ZN(G1329gat));
  NAND2_X1  g593(.A1(new_n754_), .A2(new_n724_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(KEYINPUT116), .B(G43gat), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n770_), .A2(G43gat), .A3(new_n724_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n797_), .B1(new_n798_), .B2(new_n790_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT47), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT47), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n801_), .B(new_n797_), .C1(new_n798_), .C2(new_n790_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n802_), .ZN(G1330gat));
  AOI21_X1  g602(.A(G50gat), .B1(new_n754_), .B2(new_n446_), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n770_), .A2(G50gat), .A3(new_n446_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n804_), .B1(new_n805_), .B2(new_n774_), .ZN(G1331gat));
  NOR3_X1   g605(.A1(new_n584_), .A2(new_n553_), .A3(new_n586_), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT37), .B1(new_n592_), .B2(new_n593_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n636_), .A2(new_n638_), .A3(new_n644_), .A4(new_n661_), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n692_), .A2(new_n809_), .A3(new_n810_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n684_), .A2(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(G57gat), .B1(new_n812_), .B2(new_n667_), .ZN(new_n813_));
  XOR2_X1   g612(.A(new_n813_), .B(KEYINPUT117), .Z(new_n814_));
  XNOR2_X1  g613(.A(new_n692_), .B(KEYINPUT73), .ZN(new_n815_));
  NOR4_X1   g614(.A1(new_n686_), .A2(new_n815_), .A3(new_n645_), .A4(new_n752_), .ZN(new_n816_));
  XOR2_X1   g615(.A(KEYINPUT118), .B(G57gat), .Z(new_n817_));
  NOR2_X1   g616(.A1(new_n664_), .A2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n814_), .B1(new_n816_), .B2(new_n818_), .ZN(G1332gat));
  INV_X1    g618(.A(new_n812_), .ZN(new_n820_));
  OR3_X1    g619(.A1(new_n820_), .A2(G64gat), .A3(new_n700_), .ZN(new_n821_));
  INV_X1    g620(.A(G64gat), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n822_), .B1(new_n816_), .B2(new_n510_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(KEYINPUT119), .B(KEYINPUT48), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  AND2_X1   g624(.A1(new_n823_), .A2(new_n825_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n823_), .A2(new_n825_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n821_), .B1(new_n826_), .B2(new_n827_), .ZN(G1333gat));
  NAND2_X1  g627(.A1(new_n816_), .A2(new_n724_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(G71gat), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n830_), .A2(KEYINPUT49), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n830_), .A2(KEYINPUT49), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n357_), .A2(G71gat), .ZN(new_n833_));
  XOR2_X1   g632(.A(new_n833_), .B(KEYINPUT120), .Z(new_n834_));
  OAI22_X1  g633(.A1(new_n831_), .A2(new_n832_), .B1(new_n820_), .B2(new_n834_), .ZN(G1334gat));
  OR3_X1    g634(.A1(new_n820_), .A2(G78gat), .A3(new_n512_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n816_), .A2(new_n446_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(G78gat), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n838_), .A2(KEYINPUT50), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n838_), .A2(KEYINPUT50), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n836_), .B1(new_n839_), .B2(new_n840_), .ZN(G1335gat));
  NOR3_X1   g640(.A1(new_n815_), .A2(new_n645_), .A3(new_n661_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n552_), .A2(new_n685_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n845_), .A2(new_n239_), .A3(new_n667_), .ZN(new_n846_));
  NOR3_X1   g645(.A1(new_n692_), .A2(new_n645_), .A3(new_n661_), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n768_), .A2(new_n847_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n848_), .A2(new_n407_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n846_), .B1(new_n849_), .B2(new_n239_), .ZN(G1336gat));
  NAND3_X1  g649(.A1(new_n845_), .A2(new_n240_), .A3(new_n510_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n848_), .A2(new_n510_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n851_), .B1(new_n852_), .B2(new_n240_), .ZN(G1337gat));
  NAND4_X1  g652(.A1(new_n842_), .A2(new_n724_), .A3(new_n237_), .A4(new_n843_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(KEYINPUT121), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT51), .ZN(new_n856_));
  AND2_X1   g655(.A1(new_n848_), .A2(new_n724_), .ZN(new_n857_));
  INV_X1    g656(.A(G99gat), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n855_), .B(new_n856_), .C1(new_n857_), .C2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT121), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n854_), .B(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n858_), .B1(new_n848_), .B2(new_n724_), .ZN(new_n862_));
  OAI21_X1  g661(.A(KEYINPUT51), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n859_), .A2(new_n863_), .ZN(G1338gat));
  NAND3_X1  g663(.A1(new_n845_), .A2(new_n238_), .A3(new_n446_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n768_), .A2(new_n446_), .A3(new_n847_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT52), .ZN(new_n867_));
  AND3_X1   g666(.A1(new_n866_), .A2(new_n867_), .A3(G106gat), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n867_), .B1(new_n866_), .B2(G106gat), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n865_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(KEYINPUT53), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n872_), .B(new_n865_), .C1(new_n868_), .C2(new_n869_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n871_), .A2(new_n873_), .ZN(G1339gat));
  INV_X1    g673(.A(KEYINPUT57), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n599_), .B1(new_n613_), .B2(new_n567_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n876_), .B1(new_n620_), .B2(new_n623_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(new_n642_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n878_), .B1(new_n599_), .B2(new_n628_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n879_), .B1(new_n640_), .B2(new_n643_), .ZN(new_n880_));
  AND2_X1   g679(.A1(new_n281_), .A2(new_n880_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n271_), .A2(new_n270_), .A3(new_n262_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n882_), .B1(new_n272_), .B2(KEYINPUT55), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT55), .ZN(new_n884_));
  AOI211_X1 g683(.A(new_n884_), .B(new_n270_), .C1(new_n271_), .C2(new_n262_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n278_), .B1(new_n883_), .B2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(KEYINPUT56), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT56), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n888_), .B(new_n278_), .C1(new_n883_), .C2(new_n885_), .ZN(new_n889_));
  AND3_X1   g688(.A1(new_n887_), .A2(new_n280_), .A3(new_n889_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n881_), .B1(new_n890_), .B2(new_n645_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n685_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n875_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n281_), .A2(new_n880_), .ZN(new_n894_));
  AND3_X1   g693(.A1(new_n636_), .A2(new_n638_), .A3(new_n644_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n887_), .A2(new_n280_), .A3(new_n889_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n894_), .B1(new_n895_), .B2(new_n896_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n897_), .A2(KEYINPUT57), .A3(new_n685_), .ZN(new_n898_));
  NAND4_X1  g697(.A1(new_n887_), .A2(new_n880_), .A3(new_n280_), .A4(new_n889_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT58), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n595_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n901_), .B1(new_n900_), .B2(new_n899_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n893_), .A2(new_n898_), .A3(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n752_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n810_), .A2(KEYINPUT122), .ZN(new_n905_));
  AOI22_X1  g704(.A1(new_n635_), .A2(KEYINPUT81), .B1(new_n643_), .B2(new_n640_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT122), .ZN(new_n907_));
  NAND4_X1  g706(.A1(new_n906_), .A2(new_n907_), .A3(new_n638_), .A4(new_n661_), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n905_), .A2(new_n692_), .A3(new_n595_), .A4(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(KEYINPUT123), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n285_), .A2(new_n809_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT123), .ZN(new_n912_));
  NAND4_X1  g711(.A1(new_n911_), .A2(new_n912_), .A3(new_n908_), .A4(new_n905_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n910_), .A2(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT54), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n910_), .A2(new_n913_), .A3(KEYINPUT54), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n904_), .A2(new_n916_), .A3(new_n917_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n357_), .A2(new_n446_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n919_), .A2(new_n700_), .A3(new_n667_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n920_), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT124), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(KEYINPUT59), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n918_), .A2(new_n921_), .A3(new_n923_), .ZN(new_n924_));
  AND3_X1   g723(.A1(new_n910_), .A2(new_n913_), .A3(KEYINPUT54), .ZN(new_n925_));
  AOI21_X1  g724(.A(KEYINPUT54), .B1(new_n910_), .B2(new_n913_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n925_), .A2(new_n926_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n920_), .B1(new_n927_), .B2(new_n904_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(KEYINPUT124), .B(KEYINPUT59), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n924_), .B1(new_n928_), .B2(new_n929_), .ZN(new_n930_));
  OAI21_X1  g729(.A(G113gat), .B1(new_n930_), .B2(new_n895_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n918_), .A2(new_n921_), .ZN(new_n932_));
  OR3_X1    g731(.A1(new_n932_), .A2(G113gat), .A3(new_n895_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n931_), .A2(new_n933_), .ZN(G1340gat));
  INV_X1    g733(.A(KEYINPUT60), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n935_), .B1(new_n692_), .B2(G120gat), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n918_), .A2(new_n921_), .A3(new_n936_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n937_), .A2(new_n286_), .ZN(new_n938_));
  OAI21_X1  g737(.A(G120gat), .B1(new_n930_), .B2(new_n938_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n928_), .A2(new_n935_), .A3(new_n936_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n939_), .A2(new_n940_), .ZN(G1341gat));
  NAND3_X1  g740(.A1(new_n918_), .A2(new_n661_), .A3(new_n921_), .ZN(new_n942_));
  INV_X1    g741(.A(G127gat), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n942_), .A2(new_n943_), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT125), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n944_), .A2(new_n945_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n752_), .A2(new_n943_), .ZN(new_n947_));
  OAI211_X1 g746(.A(new_n924_), .B(new_n947_), .C1(new_n928_), .C2(new_n929_), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n942_), .A2(KEYINPUT125), .A3(new_n943_), .ZN(new_n949_));
  AND3_X1   g748(.A1(new_n946_), .A2(new_n948_), .A3(new_n949_), .ZN(G1342gat));
  OAI21_X1  g749(.A(G134gat), .B1(new_n930_), .B2(new_n595_), .ZN(new_n951_));
  OR3_X1    g750(.A1(new_n932_), .A2(G134gat), .A3(new_n685_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n951_), .A2(new_n952_), .ZN(G1343gat));
  INV_X1    g752(.A(new_n667_), .ZN(new_n954_));
  NOR4_X1   g753(.A1(new_n954_), .A2(new_n724_), .A3(new_n512_), .A4(new_n510_), .ZN(new_n955_));
  AND2_X1   g754(.A1(new_n918_), .A2(new_n955_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n956_), .A2(new_n645_), .ZN(new_n957_));
  XNOR2_X1  g756(.A(new_n957_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g757(.A1(new_n956_), .A2(new_n286_), .ZN(new_n959_));
  XNOR2_X1  g758(.A(new_n959_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g759(.A1(new_n918_), .A2(new_n955_), .ZN(new_n961_));
  NOR2_X1   g760(.A1(new_n961_), .A2(new_n752_), .ZN(new_n962_));
  XOR2_X1   g761(.A(KEYINPUT61), .B(G155gat), .Z(new_n963_));
  XNOR2_X1  g762(.A(new_n962_), .B(new_n963_), .ZN(G1346gat));
  INV_X1    g763(.A(G162gat), .ZN(new_n965_));
  NOR3_X1   g764(.A1(new_n961_), .A2(new_n965_), .A3(new_n760_), .ZN(new_n966_));
  OAI21_X1  g765(.A(new_n965_), .B1(new_n961_), .B2(new_n685_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n967_), .A2(KEYINPUT126), .ZN(new_n968_));
  INV_X1    g767(.A(KEYINPUT126), .ZN(new_n969_));
  OAI211_X1 g768(.A(new_n969_), .B(new_n965_), .C1(new_n961_), .C2(new_n685_), .ZN(new_n970_));
  AOI21_X1  g769(.A(new_n966_), .B1(new_n968_), .B2(new_n970_), .ZN(G1347gat));
  NAND3_X1  g770(.A1(new_n954_), .A2(new_n919_), .A3(new_n510_), .ZN(new_n972_));
  INV_X1    g771(.A(new_n972_), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n918_), .A2(new_n973_), .ZN(new_n974_));
  OAI21_X1  g773(.A(G169gat), .B1(new_n974_), .B2(new_n895_), .ZN(new_n975_));
  INV_X1    g774(.A(KEYINPUT62), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n975_), .A2(new_n976_), .ZN(new_n977_));
  OAI211_X1 g776(.A(KEYINPUT62), .B(G169gat), .C1(new_n974_), .C2(new_n895_), .ZN(new_n978_));
  AOI21_X1  g777(.A(new_n972_), .B1(new_n927_), .B2(new_n904_), .ZN(new_n979_));
  NAND3_X1  g778(.A1(new_n979_), .A2(new_n468_), .A3(new_n645_), .ZN(new_n980_));
  NAND3_X1  g779(.A1(new_n977_), .A2(new_n978_), .A3(new_n980_), .ZN(G1348gat));
  NOR3_X1   g780(.A1(new_n974_), .A2(new_n329_), .A3(new_n815_), .ZN(new_n982_));
  AOI21_X1  g781(.A(G176gat), .B1(new_n979_), .B2(new_n285_), .ZN(new_n983_));
  NOR2_X1   g782(.A1(new_n982_), .A2(new_n983_), .ZN(G1349gat));
  OAI211_X1 g783(.A(new_n291_), .B(new_n293_), .C1(new_n974_), .C2(new_n752_), .ZN(new_n985_));
  NOR2_X1   g784(.A1(new_n462_), .A2(new_n326_), .ZN(new_n986_));
  NAND3_X1  g785(.A1(new_n979_), .A2(new_n986_), .A3(new_n661_), .ZN(new_n987_));
  AND2_X1   g786(.A1(new_n985_), .A2(new_n987_), .ZN(G1350gat));
  AOI21_X1  g787(.A(new_n294_), .B1(new_n979_), .B2(new_n809_), .ZN(new_n989_));
  AND3_X1   g788(.A1(new_n892_), .A2(new_n313_), .A3(new_n319_), .ZN(new_n990_));
  AND3_X1   g789(.A1(new_n918_), .A2(new_n973_), .A3(new_n990_), .ZN(new_n991_));
  OAI21_X1  g790(.A(KEYINPUT127), .B1(new_n989_), .B2(new_n991_), .ZN(new_n992_));
  OAI21_X1  g791(.A(G190gat), .B1(new_n974_), .B2(new_n595_), .ZN(new_n993_));
  INV_X1    g792(.A(KEYINPUT127), .ZN(new_n994_));
  NAND2_X1  g793(.A1(new_n979_), .A2(new_n990_), .ZN(new_n995_));
  NAND3_X1  g794(.A1(new_n993_), .A2(new_n994_), .A3(new_n995_), .ZN(new_n996_));
  NAND2_X1  g795(.A1(new_n992_), .A2(new_n996_), .ZN(G1351gat));
  NOR3_X1   g796(.A1(new_n724_), .A2(new_n700_), .A3(new_n546_), .ZN(new_n998_));
  NAND2_X1  g797(.A1(new_n918_), .A2(new_n998_), .ZN(new_n999_));
  NOR2_X1   g798(.A1(new_n999_), .A2(new_n895_), .ZN(new_n1000_));
  XNOR2_X1  g799(.A(new_n1000_), .B(new_n416_), .ZN(G1352gat));
  NOR2_X1   g800(.A1(new_n999_), .A2(new_n815_), .ZN(new_n1002_));
  XNOR2_X1  g801(.A(new_n1002_), .B(new_n411_), .ZN(G1353gat));
  NOR2_X1   g802(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1004_));
  OAI21_X1  g803(.A(new_n1004_), .B1(new_n999_), .B2(new_n752_), .ZN(new_n1005_));
  XOR2_X1   g804(.A(KEYINPUT63), .B(G211gat), .Z(new_n1006_));
  NAND4_X1  g805(.A1(new_n918_), .A2(new_n661_), .A3(new_n998_), .A4(new_n1006_), .ZN(new_n1007_));
  AND2_X1   g806(.A1(new_n1005_), .A2(new_n1007_), .ZN(G1354gat));
  OAI21_X1  g807(.A(G218gat), .B1(new_n999_), .B2(new_n595_), .ZN(new_n1009_));
  OR2_X1    g808(.A1(new_n685_), .A2(G218gat), .ZN(new_n1010_));
  OAI21_X1  g809(.A(new_n1009_), .B1(new_n999_), .B2(new_n1010_), .ZN(G1355gat));
endmodule


