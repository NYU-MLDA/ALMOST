//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 1 1 1 0 1 0 1 1 0 0 0 0 0 1 0 0 1 0 1 0 1 1 1 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 0 0 0 0 1 1 1 1 0 0 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n659_, new_n660_, new_n661_, new_n663_, new_n664_,
    new_n665_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n707_, new_n708_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n807_,
    new_n808_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n841_, new_n842_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n871_, new_n872_, new_n873_, new_n874_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n894_;
  INV_X1    g000(.A(G155gat), .ZN(new_n202_));
  INV_X1    g001(.A(G162gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n202_), .A2(new_n203_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT1), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n204_), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT88), .ZN(new_n208_));
  INV_X1    g007(.A(new_n205_), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n208_), .B1(KEYINPUT1), .B2(new_n209_), .ZN(new_n210_));
  OR2_X1    g009(.A1(G141gat), .A2(G148gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G141gat), .A2(G148gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(KEYINPUT89), .ZN(new_n214_));
  AOI22_X1  g013(.A1(KEYINPUT2), .A2(new_n214_), .B1(new_n211_), .B2(KEYINPUT3), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n214_), .A2(KEYINPUT2), .ZN(new_n216_));
  OAI211_X1 g015(.A(new_n215_), .B(new_n216_), .C1(KEYINPUT3), .C2(new_n211_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(new_n209_), .A3(new_n204_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n213_), .A2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(G127gat), .B(G134gat), .ZN(new_n220_));
  INV_X1    g019(.A(G113gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n220_), .B(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n222_), .B(G120gat), .ZN(new_n223_));
  OR3_X1    g022(.A1(new_n219_), .A2(KEYINPUT96), .A3(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n223_), .B1(new_n219_), .B2(KEYINPUT96), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(KEYINPUT4), .A3(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT4), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n219_), .A2(new_n227_), .A3(new_n223_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT99), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G225gat), .A2(G233gat), .ZN(new_n231_));
  XOR2_X1   g030(.A(new_n231_), .B(KEYINPUT97), .Z(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT98), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n228_), .A2(new_n229_), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n226_), .A2(new_n230_), .A3(new_n233_), .A4(new_n234_), .ZN(new_n235_));
  AND2_X1   g034(.A1(new_n224_), .A2(new_n225_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n232_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n235_), .A2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G1gat), .B(G29gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(G85gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT0), .ZN(new_n242_));
  INV_X1    g041(.A(G57gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n239_), .A2(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n235_), .A2(new_n238_), .A3(new_n244_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT27), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G169gat), .A2(G176gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT24), .ZN(new_n252_));
  NOR2_X1   g051(.A1(G169gat), .A2(G176gat), .ZN(new_n253_));
  MUX2_X1   g052(.A(new_n252_), .B(KEYINPUT24), .S(new_n253_), .Z(new_n254_));
  INV_X1    g053(.A(G190gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT26), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT26), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(G190gat), .ZN(new_n258_));
  AND2_X1   g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT25), .B(G183gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(G183gat), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT23), .B1(new_n262_), .B2(new_n255_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT23), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n264_), .A2(G183gat), .A3(G190gat), .ZN(new_n265_));
  AOI21_X1  g064(.A(KEYINPUT86), .B1(new_n263_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT86), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G183gat), .A2(G190gat), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n267_), .B1(new_n268_), .B2(KEYINPUT23), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n254_), .B(new_n261_), .C1(new_n266_), .C2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT94), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n263_), .A2(new_n265_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n272_), .B1(G183gat), .B2(G190gat), .ZN(new_n273_));
  XOR2_X1   g072(.A(KEYINPUT22), .B(G169gat), .Z(new_n274_));
  OAI211_X1 g073(.A(new_n273_), .B(new_n251_), .C1(G176gat), .C2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n271_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT21), .ZN(new_n277_));
  INV_X1    g076(.A(G204gat), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n278_), .A2(G197gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT90), .B(G204gat), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n279_), .B1(new_n280_), .B2(G197gat), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n277_), .B1(new_n281_), .B2(KEYINPUT91), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G211gat), .B(G218gat), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  OAI211_X1 g083(.A(new_n282_), .B(new_n284_), .C1(KEYINPUT91), .C2(new_n281_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n284_), .B1(new_n281_), .B2(new_n277_), .ZN(new_n286_));
  INV_X1    g085(.A(G197gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n280_), .A2(new_n287_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n288_), .B1(new_n287_), .B2(new_n278_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n286_), .B1(new_n277_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n285_), .A2(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT20), .B1(new_n276_), .B2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G226gat), .A2(G233gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT19), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  XOR2_X1   g094(.A(KEYINPUT81), .B(G183gat), .Z(new_n296_));
  INV_X1    g095(.A(KEYINPUT25), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT82), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT82), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n297_), .A2(new_n262_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT81), .B(G183gat), .ZN(new_n301_));
  OAI211_X1 g100(.A(new_n299_), .B(new_n300_), .C1(new_n301_), .C2(new_n297_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT83), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n258_), .B(new_n303_), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n298_), .A2(new_n302_), .A3(new_n256_), .A4(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n305_), .A2(new_n272_), .A3(new_n254_), .ZN(new_n306_));
  INV_X1    g105(.A(G169gat), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n307_), .A2(KEYINPUT85), .ZN(new_n308_));
  NAND2_X1  g107(.A1(KEYINPUT84), .A2(KEYINPUT22), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(G176gat), .ZN(new_n311_));
  OAI21_X1  g110(.A(KEYINPUT22), .B1(KEYINPUT84), .B2(G169gat), .ZN(new_n312_));
  OAI211_X1 g111(.A(new_n310_), .B(new_n311_), .C1(new_n308_), .C2(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n266_), .A2(new_n269_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n296_), .A2(G190gat), .ZN(new_n315_));
  OAI211_X1 g114(.A(new_n251_), .B(new_n313_), .C1(new_n314_), .C2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n306_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(new_n291_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT95), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n295_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n276_), .A2(new_n291_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(KEYINPUT20), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n317_), .A2(new_n291_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n294_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  AND2_X1   g124(.A1(new_n321_), .A2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G8gat), .B(G36gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT18), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(G64gat), .ZN(new_n329_));
  INV_X1    g128(.A(G92gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  AND2_X1   g130(.A1(new_n326_), .A2(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n326_), .A2(new_n331_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n250_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n326_), .A2(new_n331_), .ZN(new_n335_));
  NOR3_X1   g134(.A1(new_n323_), .A2(new_n294_), .A3(new_n324_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n275_), .A2(new_n270_), .ZN(new_n337_));
  OAI211_X1 g136(.A(new_n320_), .B(KEYINPUT20), .C1(new_n291_), .C2(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n336_), .B1(new_n338_), .B2(new_n294_), .ZN(new_n339_));
  OAI211_X1 g138(.A(new_n335_), .B(KEYINPUT27), .C1(new_n331_), .C2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n334_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  AND2_X1   g141(.A1(new_n213_), .A2(new_n218_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT29), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n291_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G228gat), .A2(G233gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(G50gat), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT28), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n343_), .A2(new_n349_), .A3(new_n344_), .ZN(new_n350_));
  INV_X1    g149(.A(G22gat), .ZN(new_n351_));
  OAI21_X1  g150(.A(KEYINPUT28), .B1(new_n219_), .B2(KEYINPUT29), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n350_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n351_), .B1(new_n350_), .B2(new_n352_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n348_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n350_), .A2(new_n352_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(G22gat), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n358_), .A2(G50gat), .A3(new_n353_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G78gat), .B(G106gat), .ZN(new_n360_));
  XOR2_X1   g159(.A(new_n360_), .B(KEYINPUT92), .Z(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT93), .ZN(new_n363_));
  AND3_X1   g162(.A1(new_n356_), .A2(new_n359_), .A3(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n361_), .B1(new_n356_), .B2(new_n359_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n347_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n356_), .A2(new_n359_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(new_n362_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n347_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n356_), .A2(new_n359_), .A3(new_n363_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n368_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n317_), .B(KEYINPUT30), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(new_n223_), .ZN(new_n373_));
  XOR2_X1   g172(.A(G71gat), .B(G99gat), .Z(new_n374_));
  NAND2_X1  g173(.A1(G227gat), .A2(G233gat), .ZN(new_n375_));
  XOR2_X1   g174(.A(new_n374_), .B(new_n375_), .Z(new_n376_));
  XNOR2_X1  g175(.A(new_n373_), .B(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(KEYINPUT87), .B(G15gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(KEYINPUT31), .B(G43gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n377_), .A2(new_n381_), .ZN(new_n382_));
  OR2_X1    g181(.A1(new_n373_), .A2(new_n376_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n373_), .A2(new_n376_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n383_), .A2(new_n380_), .A3(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n382_), .A2(new_n385_), .ZN(new_n386_));
  AND3_X1   g185(.A1(new_n366_), .A2(new_n371_), .A3(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n386_), .B1(new_n366_), .B2(new_n371_), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n249_), .B(new_n342_), .C1(new_n387_), .C2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n247_), .A2(KEYINPUT100), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(KEYINPUT33), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n332_), .A2(new_n333_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n236_), .A2(new_n233_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n226_), .A2(new_n234_), .A3(new_n230_), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n245_), .B(new_n393_), .C1(new_n394_), .C2(new_n232_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT33), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n247_), .A2(KEYINPUT100), .A3(new_n396_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n391_), .A2(new_n392_), .A3(new_n395_), .A4(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n331_), .A2(KEYINPUT32), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n326_), .A2(new_n399_), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n248_), .B(new_n400_), .C1(new_n339_), .C2(new_n399_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n398_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n366_), .A2(new_n371_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n402_), .A2(new_n386_), .A3(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n389_), .A2(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT69), .B(KEYINPUT12), .ZN(new_n406_));
  NOR2_X1   g205(.A1(G99gat), .A2(G106gat), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT7), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT67), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n408_), .A2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(KEYINPUT67), .B(KEYINPUT7), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n411_), .B1(new_n412_), .B2(new_n408_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G99gat), .A2(G106gat), .ZN(new_n414_));
  AND2_X1   g213(.A1(KEYINPUT68), .A2(KEYINPUT6), .ZN(new_n415_));
  NOR2_X1   g214(.A1(KEYINPUT68), .A2(KEYINPUT6), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n414_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT68), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT6), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  AND2_X1   g219(.A1(G99gat), .A2(G106gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(KEYINPUT68), .A2(KEYINPUT6), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n420_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n417_), .A2(new_n423_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n413_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(G85gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(new_n330_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G85gat), .A2(G92gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT8), .B1(new_n425_), .B2(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n429_), .A2(KEYINPUT8), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n419_), .A2(KEYINPUT65), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT65), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT6), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n432_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n421_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n432_), .A2(new_n434_), .A3(new_n414_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n431_), .B1(new_n438_), .B2(new_n413_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n428_), .A2(KEYINPUT9), .ZN(new_n440_));
  INV_X1    g239(.A(G99gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT10), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT10), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(G99gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(G106gat), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n440_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n427_), .A2(KEYINPUT9), .A3(new_n428_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n447_), .A2(new_n436_), .A3(new_n437_), .A4(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT66), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n437_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n414_), .B1(new_n432_), .B2(new_n434_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n454_), .A2(KEYINPUT66), .A3(new_n448_), .A4(new_n447_), .ZN(new_n455_));
  AOI22_X1  g254(.A1(new_n430_), .A2(new_n439_), .B1(new_n451_), .B2(new_n455_), .ZN(new_n456_));
  XOR2_X1   g255(.A(G71gat), .B(G78gat), .Z(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G57gat), .B(G64gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT11), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n458_), .A2(new_n460_), .ZN(new_n461_));
  OR2_X1    g260(.A1(new_n459_), .A2(KEYINPUT11), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n457_), .A2(KEYINPUT11), .A3(new_n459_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n461_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n406_), .B1(new_n456_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n451_), .A2(new_n455_), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n417_), .A2(new_n423_), .ZN(new_n468_));
  AOI22_X1  g267(.A1(new_n441_), .A2(new_n446_), .B1(new_n409_), .B2(KEYINPUT67), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT67), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT7), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n410_), .A2(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n469_), .B1(new_n407_), .B2(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n429_), .B1(new_n468_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT8), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n439_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n467_), .A2(new_n476_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(KEYINPUT69), .A2(KEYINPUT12), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n477_), .A2(new_n464_), .A3(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G230gat), .A2(G233gat), .ZN(new_n481_));
  XOR2_X1   g280(.A(new_n481_), .B(KEYINPUT64), .Z(new_n482_));
  NAND2_X1  g281(.A1(new_n456_), .A2(new_n465_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n466_), .A2(new_n480_), .A3(new_n482_), .A4(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n482_), .ZN(new_n485_));
  AND3_X1   g284(.A1(new_n467_), .A2(new_n476_), .A3(new_n465_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n465_), .B1(new_n467_), .B2(new_n476_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n485_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G120gat), .B(G148gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G176gat), .B(G204gat), .ZN(new_n492_));
  XOR2_X1   g291(.A(new_n491_), .B(new_n492_), .Z(new_n493_));
  NAND3_X1  g292(.A1(new_n484_), .A2(new_n488_), .A3(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n493_), .B1(new_n484_), .B2(new_n488_), .ZN(new_n496_));
  AND2_X1   g295(.A1(KEYINPUT71), .A2(KEYINPUT13), .ZN(new_n497_));
  OR3_X1    g296(.A1(new_n495_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(KEYINPUT71), .A2(KEYINPUT13), .ZN(new_n499_));
  OAI22_X1  g298(.A1(new_n495_), .A2(new_n496_), .B1(new_n497_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n498_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT77), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G29gat), .B(G36gat), .ZN(new_n504_));
  INV_X1    g303(.A(G43gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(G50gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n504_), .B(G43gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(new_n348_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G15gat), .B(G22gat), .ZN(new_n510_));
  INV_X1    g309(.A(G1gat), .ZN(new_n511_));
  INV_X1    g310(.A(G8gat), .ZN(new_n512_));
  OAI21_X1  g311(.A(KEYINPUT14), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n510_), .A2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G1gat), .B(G8gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  OR2_X1    g315(.A1(new_n514_), .A2(new_n515_), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n507_), .A2(new_n509_), .A3(new_n516_), .A4(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  AOI22_X1  g318(.A1(new_n507_), .A2(new_n509_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n503_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n520_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n522_), .A2(KEYINPUT77), .A3(new_n518_), .ZN(new_n523_));
  AND2_X1   g322(.A1(G229gat), .A2(G233gat), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n521_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n517_), .A2(new_n516_), .ZN(new_n526_));
  AND3_X1   g325(.A1(new_n507_), .A2(new_n509_), .A3(KEYINPUT15), .ZN(new_n527_));
  AOI21_X1  g326(.A(KEYINPUT15), .B1(new_n507_), .B2(new_n509_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n526_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n524_), .B(KEYINPUT78), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n529_), .A2(new_n518_), .A3(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n525_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G169gat), .B(G197gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G113gat), .B(G141gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(KEYINPUT79), .B(KEYINPUT80), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n533_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n538_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n525_), .A2(new_n532_), .A3(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n502_), .A2(new_n543_), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n405_), .A2(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n477_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n456_), .A2(new_n507_), .A3(new_n509_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G232gat), .A2(G233gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT34), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n549_), .A2(KEYINPUT35), .ZN(new_n550_));
  XOR2_X1   g349(.A(new_n550_), .B(KEYINPUT73), .Z(new_n551_));
  NAND3_X1  g350(.A1(new_n546_), .A2(new_n547_), .A3(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n549_), .A2(KEYINPUT35), .ZN(new_n553_));
  XOR2_X1   g352(.A(new_n553_), .B(KEYINPUT72), .Z(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  OR2_X1    g354(.A1(new_n552_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n552_), .A2(new_n555_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G190gat), .B(G218gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(G134gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(new_n203_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n556_), .A2(KEYINPUT36), .A3(new_n557_), .A4(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n556_), .A2(new_n557_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT74), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n561_), .A2(KEYINPUT36), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n563_), .A2(new_n564_), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n565_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n562_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT37), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  OAI211_X1 g370(.A(KEYINPUT37), .B(new_n562_), .C1(new_n567_), .C2(new_n568_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n526_), .B(new_n464_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G231gat), .A2(G233gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT75), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G127gat), .B(G155gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT16), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(G183gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(G211gat), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(KEYINPUT17), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT76), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n578_), .A2(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n577_), .B1(KEYINPUT17), .B2(new_n582_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n586_), .B1(KEYINPUT17), .B2(new_n582_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n574_), .A2(new_n589_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n545_), .A2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n591_), .A2(new_n511_), .A3(new_n248_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n592_), .A2(KEYINPUT38), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n592_), .A2(KEYINPUT38), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT101), .ZN(new_n595_));
  INV_X1    g394(.A(new_n569_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(new_n588_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n545_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(new_n248_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n595_), .B1(new_n601_), .B2(G1gat), .ZN(new_n602_));
  AOI211_X1 g401(.A(KEYINPUT101), .B(new_n511_), .C1(new_n600_), .C2(new_n248_), .ZN(new_n603_));
  OAI22_X1  g402(.A1(new_n593_), .A2(new_n594_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(KEYINPUT102), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT102), .ZN(new_n606_));
  OAI221_X1 g405(.A(new_n606_), .B1(new_n602_), .B2(new_n603_), .C1(new_n593_), .C2(new_n594_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n607_), .ZN(G1324gat));
  NAND3_X1  g407(.A1(new_n591_), .A2(new_n512_), .A3(new_n341_), .ZN(new_n609_));
  OAI21_X1  g408(.A(G8gat), .B1(new_n599_), .B2(new_n342_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n610_), .A2(KEYINPUT39), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n610_), .A2(KEYINPUT39), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n609_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT40), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(G1325gat));
  OAI21_X1  g414(.A(G15gat), .B1(new_n599_), .B2(new_n386_), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n616_), .B(KEYINPUT41), .Z(new_n617_));
  INV_X1    g416(.A(G15gat), .ZN(new_n618_));
  INV_X1    g417(.A(new_n386_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n591_), .A2(new_n618_), .A3(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n617_), .A2(new_n620_), .ZN(G1326gat));
  INV_X1    g420(.A(KEYINPUT103), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n403_), .B(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  OAI21_X1  g423(.A(G22gat), .B1(new_n599_), .B2(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(KEYINPUT104), .B(KEYINPUT42), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n591_), .A2(new_n351_), .A3(new_n623_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(G1327gat));
  NOR2_X1   g428(.A1(new_n596_), .A2(new_n588_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n545_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(G29gat), .B1(new_n632_), .B2(new_n248_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n544_), .A2(new_n589_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT43), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n636_), .B1(new_n405_), .B2(new_n574_), .ZN(new_n637_));
  AOI211_X1 g436(.A(KEYINPUT43), .B(new_n573_), .C1(new_n389_), .C2(new_n404_), .ZN(new_n638_));
  OAI211_X1 g437(.A(KEYINPUT44), .B(new_n635_), .C1(new_n637_), .C2(new_n638_), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n639_), .A2(G29gat), .A3(new_n248_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n635_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT44), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n633_), .B1(new_n640_), .B2(new_n643_), .ZN(G1328gat));
  INV_X1    g443(.A(G36gat), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n545_), .A2(new_n645_), .A3(new_n341_), .A4(new_n630_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n646_), .A2(KEYINPUT45), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n646_), .A2(KEYINPUT45), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT105), .ZN(new_n649_));
  OAI22_X1  g448(.A1(new_n647_), .A2(new_n648_), .B1(new_n649_), .B2(KEYINPUT46), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n342_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n645_), .B1(new_n651_), .B2(new_n639_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n649_), .A2(KEYINPUT46), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT106), .Z(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  OR3_X1    g454(.A1(new_n650_), .A2(new_n652_), .A3(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n655_), .B1(new_n650_), .B2(new_n652_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(G1329gat));
  OAI21_X1  g457(.A(new_n505_), .B1(new_n631_), .B2(new_n386_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n643_), .A2(G43gat), .A3(new_n639_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n659_), .B1(new_n660_), .B2(new_n386_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g461(.A(new_n403_), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n643_), .A2(G50gat), .A3(new_n663_), .A4(new_n639_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n348_), .B1(new_n631_), .B2(new_n624_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1331gat));
  NOR2_X1   g465(.A1(new_n501_), .A2(new_n542_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n405_), .A2(new_n667_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n668_), .A2(new_n597_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n243_), .B1(new_n669_), .B2(new_n248_), .ZN(new_n670_));
  NOR3_X1   g469(.A1(new_n668_), .A2(new_n589_), .A3(new_n574_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n249_), .A2(G57gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n670_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT107), .ZN(G1332gat));
  INV_X1    g473(.A(G64gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n675_), .B1(new_n669_), .B2(new_n341_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT48), .Z(new_n677_));
  NAND3_X1  g476(.A1(new_n671_), .A2(new_n675_), .A3(new_n341_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1333gat));
  NAND2_X1  g478(.A1(new_n669_), .A2(new_n619_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(G71gat), .ZN(new_n681_));
  XNOR2_X1  g480(.A(KEYINPUT108), .B(KEYINPUT49), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n681_), .B(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n671_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n386_), .A2(G71gat), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT109), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n683_), .B1(new_n684_), .B2(new_n686_), .ZN(G1334gat));
  INV_X1    g486(.A(G78gat), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n671_), .A2(new_n688_), .A3(new_n623_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n669_), .B2(new_n623_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT50), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n690_), .A2(new_n691_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n689_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT110), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n694_), .B(new_n695_), .ZN(G1335gat));
  NOR3_X1   g495(.A1(new_n668_), .A2(new_n596_), .A3(new_n588_), .ZN(new_n697_));
  AOI21_X1  g496(.A(G85gat), .B1(new_n697_), .B2(new_n248_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n637_), .A2(new_n638_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT111), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n501_), .A2(new_n588_), .A3(new_n542_), .ZN(new_n702_));
  OAI21_X1  g501(.A(KEYINPUT111), .B1(new_n637_), .B2(new_n638_), .ZN(new_n703_));
  AND3_X1   g502(.A1(new_n701_), .A2(new_n702_), .A3(new_n703_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n249_), .A2(new_n426_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n698_), .B1(new_n704_), .B2(new_n705_), .ZN(G1336gat));
  AOI21_X1  g505(.A(G92gat), .B1(new_n697_), .B2(new_n341_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n342_), .A2(new_n330_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n707_), .B1(new_n704_), .B2(new_n708_), .ZN(G1337gat));
  NAND4_X1  g508(.A1(new_n701_), .A2(new_n619_), .A3(new_n702_), .A4(new_n703_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(G99gat), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n697_), .A2(new_n445_), .A3(new_n619_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT51), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n714_), .A2(KEYINPUT112), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n713_), .B(new_n715_), .ZN(G1338gat));
  OAI211_X1 g515(.A(new_n663_), .B(new_n702_), .C1(new_n637_), .C2(new_n638_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(G106gat), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT113), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n717_), .A2(KEYINPUT113), .A3(G106gat), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n720_), .A2(KEYINPUT52), .A3(new_n721_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n697_), .A2(new_n446_), .A3(new_n663_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT52), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n718_), .A2(new_n719_), .A3(new_n724_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n722_), .A2(new_n723_), .A3(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT53), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT53), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n722_), .A2(new_n728_), .A3(new_n723_), .A4(new_n725_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(G1339gat));
  NOR2_X1   g529(.A1(new_n341_), .A2(new_n249_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(new_n388_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT55), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n466_), .A2(new_n483_), .A3(new_n480_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n734_), .B2(new_n485_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n484_), .A2(KEYINPUT114), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n484_), .A2(KEYINPUT114), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n735_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n493_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n484_), .A2(KEYINPUT114), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n486_), .B1(new_n487_), .B2(new_n479_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT114), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n741_), .A2(new_n742_), .A3(new_n482_), .A4(new_n466_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n482_), .B1(new_n741_), .B2(new_n466_), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n740_), .B(new_n743_), .C1(new_n744_), .C2(new_n733_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n738_), .A2(new_n739_), .A3(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT56), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n738_), .A2(new_n745_), .A3(KEYINPUT56), .A4(new_n739_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n495_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n521_), .A2(new_n523_), .A3(new_n531_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n529_), .A2(new_n518_), .A3(new_n530_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n751_), .A2(new_n752_), .A3(new_n538_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n541_), .A2(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(KEYINPUT58), .B1(new_n750_), .B2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n750_), .A2(KEYINPUT58), .A3(new_n754_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n756_), .A2(new_n574_), .A3(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n542_), .A2(new_n494_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n759_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n754_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT115), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n754_), .B(KEYINPUT115), .C1(new_n495_), .C2(new_n496_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n596_), .B1(new_n760_), .B2(new_n765_), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n766_), .A2(KEYINPUT116), .A3(KEYINPUT57), .ZN(new_n767_));
  AOI21_X1  g566(.A(KEYINPUT57), .B1(new_n766_), .B2(KEYINPUT116), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n758_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT117), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n758_), .B(KEYINPUT117), .C1(new_n767_), .C2(new_n768_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n771_), .A2(new_n589_), .A3(new_n772_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n573_), .A2(new_n543_), .A3(new_n501_), .A4(new_n588_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT54), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n732_), .B1(new_n773_), .B2(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(G113gat), .B1(new_n776_), .B2(new_n542_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n773_), .A2(new_n775_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n732_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT59), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n766_), .A2(KEYINPUT116), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT57), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n766_), .A2(KEYINPUT116), .A3(KEYINPUT57), .ZN(new_n785_));
  AND3_X1   g584(.A1(new_n750_), .A2(KEYINPUT58), .A3(new_n754_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n786_), .A2(new_n755_), .ZN(new_n787_));
  AOI22_X1  g586(.A1(new_n784_), .A2(new_n785_), .B1(new_n787_), .B2(new_n574_), .ZN(new_n788_));
  OAI21_X1  g587(.A(KEYINPUT118), .B1(new_n788_), .B2(new_n588_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT118), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n769_), .A2(new_n790_), .A3(new_n589_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n789_), .A2(new_n775_), .A3(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT59), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n792_), .A2(new_n793_), .A3(new_n779_), .ZN(new_n794_));
  AND2_X1   g593(.A1(new_n781_), .A2(new_n794_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n543_), .A2(new_n221_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n777_), .B1(new_n795_), .B2(new_n796_), .ZN(G1340gat));
  OAI211_X1 g596(.A(new_n794_), .B(new_n502_), .C1(new_n793_), .C2(new_n776_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT119), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT119), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n781_), .A2(new_n800_), .A3(new_n502_), .A4(new_n794_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n799_), .A2(new_n801_), .A3(G120gat), .ZN(new_n802_));
  INV_X1    g601(.A(G120gat), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n803_), .B1(new_n501_), .B2(KEYINPUT60), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n776_), .B(new_n804_), .C1(KEYINPUT60), .C2(new_n803_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n802_), .A2(new_n805_), .ZN(G1341gat));
  AOI21_X1  g605(.A(G127gat), .B1(new_n776_), .B2(new_n588_), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n588_), .A2(G127gat), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n807_), .B1(new_n795_), .B2(new_n808_), .ZN(G1342gat));
  INV_X1    g608(.A(G134gat), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n573_), .A2(new_n810_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n794_), .B(new_n811_), .C1(new_n793_), .C2(new_n776_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n810_), .B1(new_n780_), .B2(new_n596_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n814_), .B(KEYINPUT120), .ZN(G1343gat));
  INV_X1    g614(.A(new_n387_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n816_), .B1(new_n773_), .B2(new_n775_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT121), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n817_), .A2(new_n818_), .A3(new_n731_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n818_), .B1(new_n817_), .B2(new_n731_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n542_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(KEYINPUT122), .B(G141gat), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n817_), .A2(new_n731_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT121), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n819_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n823_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n827_), .A2(new_n542_), .A3(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n824_), .A2(new_n829_), .ZN(G1344gat));
  OAI21_X1  g629(.A(new_n502_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(G148gat), .ZN(new_n832_));
  INV_X1    g631(.A(G148gat), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n827_), .A2(new_n833_), .A3(new_n502_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n832_), .A2(new_n834_), .ZN(G1345gat));
  XNOR2_X1  g634(.A(KEYINPUT61), .B(G155gat), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n836_), .B1(new_n827_), .B2(new_n588_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n836_), .ZN(new_n838_));
  AOI211_X1 g637(.A(new_n589_), .B(new_n838_), .C1(new_n826_), .C2(new_n819_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n837_), .A2(new_n839_), .ZN(G1346gat));
  AOI21_X1  g639(.A(G162gat), .B1(new_n827_), .B2(new_n569_), .ZN(new_n841_));
  AOI211_X1 g640(.A(new_n203_), .B(new_n573_), .C1(new_n826_), .C2(new_n819_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n841_), .A2(new_n842_), .ZN(G1347gat));
  NOR2_X1   g642(.A1(new_n342_), .A2(new_n248_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n619_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n845_), .A2(new_n623_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n792_), .A2(new_n542_), .A3(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(G169gat), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT62), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  OR2_X1    g649(.A1(new_n847_), .A2(new_n274_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n847_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n850_), .A2(new_n851_), .A3(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT123), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n850_), .A2(new_n851_), .A3(KEYINPUT123), .A4(new_n852_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(G1348gat));
  INV_X1    g656(.A(new_n792_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n846_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(G176gat), .B1(new_n860_), .B2(new_n502_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n663_), .B1(new_n773_), .B2(new_n775_), .ZN(new_n862_));
  NOR3_X1   g661(.A1(new_n845_), .A2(new_n311_), .A3(new_n501_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n861_), .B1(new_n862_), .B2(new_n863_), .ZN(G1349gat));
  INV_X1    g663(.A(new_n845_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n862_), .A2(new_n588_), .A3(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT124), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n866_), .B(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n589_), .A2(new_n260_), .ZN(new_n869_));
  AOI22_X1  g668(.A1(new_n868_), .A2(new_n301_), .B1(new_n860_), .B2(new_n869_), .ZN(G1350gat));
  NAND2_X1  g669(.A1(new_n569_), .A2(new_n259_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(KEYINPUT125), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n860_), .A2(new_n872_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n858_), .A2(new_n573_), .A3(new_n859_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n873_), .B1(new_n255_), .B2(new_n874_), .ZN(G1351gat));
  NAND2_X1  g674(.A1(new_n817_), .A2(new_n844_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT126), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n817_), .A2(KEYINPUT126), .A3(new_n844_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(G197gat), .B1(new_n880_), .B2(new_n542_), .ZN(new_n881_));
  AOI211_X1 g680(.A(new_n287_), .B(new_n543_), .C1(new_n878_), .C2(new_n879_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n881_), .A2(new_n882_), .ZN(G1352gat));
  NAND3_X1  g682(.A1(new_n880_), .A2(new_n502_), .A3(new_n280_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n501_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n278_), .B2(new_n885_), .ZN(G1353gat));
  OR2_X1    g685(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n887_), .B1(new_n880_), .B2(new_n588_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(KEYINPUT63), .B(G211gat), .ZN(new_n889_));
  AOI211_X1 g688(.A(new_n589_), .B(new_n889_), .C1(new_n878_), .C2(new_n879_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n888_), .A2(new_n890_), .ZN(G1354gat));
  AOI21_X1  g690(.A(G218gat), .B1(new_n880_), .B2(new_n569_), .ZN(new_n892_));
  INV_X1    g691(.A(G218gat), .ZN(new_n893_));
  AOI211_X1 g692(.A(new_n893_), .B(new_n573_), .C1(new_n878_), .C2(new_n879_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n892_), .A2(new_n894_), .ZN(G1355gat));
endmodule


