//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 1 1 0 1 0 1 0 0 1 1 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 0 0 0 1 0 1 1 0 0 0 0 1 1 1 0 0 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n645_, new_n646_, new_n647_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n753_, new_n754_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n848_, new_n849_, new_n850_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n859_, new_n860_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n894_,
    new_n895_, new_n897_, new_n898_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_;
  XOR2_X1   g000(.A(G71gat), .B(G78gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G57gat), .B(G64gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(new_n202_), .B1(KEYINPUT11), .B2(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT69), .ZN(new_n205_));
  AND2_X1   g004(.A1(new_n203_), .A2(KEYINPUT11), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  XOR2_X1   g006(.A(KEYINPUT10), .B(G99gat), .Z(new_n208_));
  INV_X1    g007(.A(G106gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  OR2_X1    g009(.A1(new_n210_), .A2(KEYINPUT65), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G85gat), .A2(G92gat), .ZN(new_n212_));
  AND2_X1   g011(.A1(G85gat), .A2(G92gat), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n212_), .B1(new_n213_), .B2(KEYINPUT9), .ZN(new_n214_));
  XOR2_X1   g013(.A(KEYINPUT66), .B(G85gat), .Z(new_n215_));
  INV_X1    g014(.A(G92gat), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n214_), .B1(new_n217_), .B2(KEYINPUT9), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n210_), .A2(KEYINPUT65), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G99gat), .A2(G106gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(KEYINPUT6), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n211_), .A2(new_n218_), .A3(new_n219_), .A4(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT67), .ZN(new_n223_));
  OR4_X1    g022(.A1(new_n223_), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n224_));
  OAI22_X1  g023(.A1(new_n223_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n221_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n213_), .A2(new_n212_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n228_), .B1(KEYINPUT68), .B2(KEYINPUT8), .ZN(new_n229_));
  NAND2_X1  g028(.A1(KEYINPUT68), .A2(KEYINPUT8), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n230_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n222_), .B1(new_n229_), .B2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n207_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT70), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT12), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n233_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  OR2_X1    g035(.A1(new_n207_), .A2(new_n232_), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n233_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n239_), .B1(KEYINPUT70), .B2(KEYINPUT12), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G230gat), .A2(G233gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT64), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n238_), .A2(new_n240_), .A3(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT71), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n237_), .A2(new_n233_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n242_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n238_), .A2(new_n240_), .A3(KEYINPUT71), .A4(new_n242_), .ZN(new_n249_));
  AND3_X1   g048(.A1(new_n245_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G120gat), .B(G148gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT5), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G176gat), .B(G204gat), .ZN(new_n253_));
  XOR2_X1   g052(.A(new_n252_), .B(new_n253_), .Z(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT72), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n250_), .A2(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n245_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n257_), .A2(KEYINPUT72), .A3(new_n254_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  OR2_X1    g058(.A1(KEYINPUT73), .A2(KEYINPUT13), .ZN(new_n260_));
  NAND2_X1  g059(.A1(KEYINPUT73), .A2(KEYINPUT13), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n259_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n256_), .A2(KEYINPUT73), .A3(new_n258_), .A4(KEYINPUT13), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT79), .B(G15gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(G22gat), .ZN(new_n266_));
  XOR2_X1   g065(.A(KEYINPUT80), .B(G8gat), .Z(new_n267_));
  INV_X1    g066(.A(G1gat), .ZN(new_n268_));
  OAI21_X1  g067(.A(KEYINPUT14), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n266_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G1gat), .B(G8gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  XOR2_X1   g071(.A(G29gat), .B(G36gat), .Z(new_n273_));
  XNOR2_X1  g072(.A(G43gat), .B(G50gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n272_), .B(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G229gat), .A2(G233gat), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n272_), .A2(new_n275_), .ZN(new_n281_));
  XOR2_X1   g080(.A(new_n275_), .B(KEYINPUT15), .Z(new_n282_));
  AOI21_X1  g081(.A(new_n281_), .B1(new_n272_), .B2(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n280_), .B1(new_n279_), .B2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G113gat), .B(G141gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G169gat), .B(G197gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n284_), .B(new_n287_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n264_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(G228gat), .ZN(new_n290_));
  INV_X1    g089(.A(G233gat), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  OR2_X1    g092(.A1(G197gat), .A2(G204gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G197gat), .A2(G204gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(KEYINPUT90), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT90), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n294_), .A2(new_n298_), .A3(new_n295_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(G211gat), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n301_), .A2(G218gat), .ZN(new_n302_));
  INV_X1    g101(.A(G218gat), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n303_), .A2(G211gat), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n300_), .A2(KEYINPUT21), .A3(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n305_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT89), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT21), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n308_), .B1(new_n296_), .B2(new_n309_), .ZN(new_n310_));
  AND2_X1   g109(.A1(G197gat), .A2(G204gat), .ZN(new_n311_));
  NOR2_X1   g110(.A1(G197gat), .A2(G204gat), .ZN(new_n312_));
  OAI211_X1 g111(.A(new_n308_), .B(new_n309_), .C1(new_n311_), .C2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n307_), .B1(new_n310_), .B2(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n294_), .A2(KEYINPUT21), .A3(new_n295_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT88), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT88), .ZN(new_n318_));
  NAND4_X1  g117(.A1(new_n294_), .A2(new_n318_), .A3(KEYINPUT21), .A4(new_n295_), .ZN(new_n319_));
  AND2_X1   g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n306_), .B1(new_n315_), .B2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G155gat), .A2(G162gat), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(G155gat), .A2(G162gat), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  OR2_X1    g125(.A1(G141gat), .A2(G148gat), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT85), .B1(new_n327_), .B2(KEYINPUT3), .ZN(new_n328_));
  NOR2_X1   g127(.A1(G141gat), .A2(G148gat), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT85), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT3), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n329_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G141gat), .A2(G148gat), .ZN(new_n333_));
  OR2_X1    g132(.A1(new_n333_), .A2(KEYINPUT2), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(KEYINPUT2), .ZN(new_n335_));
  AOI22_X1  g134(.A1(new_n328_), .A2(new_n332_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n337_));
  XOR2_X1   g136(.A(new_n337_), .B(KEYINPUT86), .Z(new_n338_));
  AOI21_X1  g137(.A(new_n326_), .B1(new_n336_), .B2(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n324_), .B1(KEYINPUT1), .B2(new_n322_), .ZN(new_n340_));
  OR2_X1    g139(.A1(new_n322_), .A2(KEYINPUT1), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n342_), .A2(new_n327_), .A3(new_n333_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(KEYINPUT87), .B1(new_n339_), .B2(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n333_), .B(KEYINPUT2), .ZN(new_n346_));
  INV_X1    g145(.A(new_n332_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n330_), .B1(new_n329_), .B2(new_n331_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n346_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n337_), .B(KEYINPUT86), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n325_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT87), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n351_), .A2(new_n352_), .A3(new_n343_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n345_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT29), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n293_), .B(new_n321_), .C1(new_n354_), .C2(new_n355_), .ZN(new_n356_));
  XOR2_X1   g155(.A(KEYINPUT91), .B(KEYINPUT29), .Z(new_n357_));
  OAI21_X1  g156(.A(new_n357_), .B1(new_n339_), .B2(new_n344_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n293_), .B1(new_n358_), .B2(new_n321_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G78gat), .B(G106gat), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  AND3_X1   g161(.A1(new_n356_), .A2(new_n360_), .A3(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n362_), .B1(new_n356_), .B2(new_n360_), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT92), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n321_), .A2(new_n293_), .ZN(new_n366_));
  AND2_X1   g165(.A1(new_n345_), .A2(new_n353_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n366_), .B1(new_n367_), .B2(KEYINPUT29), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n361_), .B1(new_n368_), .B2(new_n359_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT92), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n356_), .A2(new_n360_), .A3(new_n362_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n369_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  XOR2_X1   g171(.A(G22gat), .B(G50gat), .Z(new_n373_));
  INV_X1    g172(.A(KEYINPUT28), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n354_), .A2(new_n374_), .A3(new_n355_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n374_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n373_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n377_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n373_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n379_), .A2(new_n375_), .A3(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n378_), .A2(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n365_), .A2(new_n372_), .A3(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n369_), .A2(new_n371_), .ZN(new_n384_));
  NAND4_X1  g183(.A1(new_n384_), .A2(KEYINPUT92), .A3(new_n381_), .A4(new_n378_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n383_), .A2(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(G169gat), .A2(G176gat), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT24), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G183gat), .A2(G190gat), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT23), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n389_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G169gat), .A2(G176gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(KEYINPUT24), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n396_), .A2(new_n387_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n394_), .A2(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT25), .B(G183gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT26), .B(G190gat), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT83), .ZN(new_n401_));
  AND3_X1   g200(.A1(new_n399_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n401_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n398_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(KEYINPUT22), .B(G169gat), .ZN(new_n405_));
  INV_X1    g204(.A(G176gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  OAI211_X1 g206(.A(new_n392_), .B(new_n393_), .C1(G183gat), .C2(G190gat), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n407_), .A2(new_n408_), .A3(new_n395_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n404_), .A2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(KEYINPUT30), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G71gat), .B(G99gat), .ZN(new_n412_));
  INV_X1    g211(.A(G43gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n412_), .B(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G227gat), .A2(G233gat), .ZN(new_n415_));
  XOR2_X1   g214(.A(new_n415_), .B(G15gat), .Z(new_n416_));
  XNOR2_X1  g215(.A(new_n414_), .B(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n411_), .B(new_n417_), .ZN(new_n418_));
  XOR2_X1   g217(.A(new_n418_), .B(KEYINPUT31), .Z(new_n419_));
  XNOR2_X1  g218(.A(G127gat), .B(G134gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G113gat), .B(G120gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(KEYINPUT84), .ZN(new_n423_));
  OR2_X1    g222(.A1(new_n419_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n419_), .A2(new_n423_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n423_), .A2(new_n345_), .A3(new_n353_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n351_), .A2(new_n422_), .A3(new_n343_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G225gat), .A2(G233gat), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT98), .B1(new_n429_), .B2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT98), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n427_), .A2(new_n433_), .A3(new_n428_), .A4(new_n430_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n432_), .A2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G1gat), .B(G29gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(KEYINPUT0), .ZN(new_n437_));
  INV_X1    g236(.A(G57gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(G85gat), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT4), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n427_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n441_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n431_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  AND3_X1   g244(.A1(new_n435_), .A2(new_n440_), .A3(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n440_), .B1(new_n435_), .B2(new_n445_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n426_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT27), .ZN(new_n451_));
  XOR2_X1   g250(.A(G8gat), .B(G36gat), .Z(new_n452_));
  XNOR2_X1  g251(.A(G64gat), .B(G92gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT96), .ZN(new_n458_));
  OAI21_X1  g257(.A(KEYINPUT20), .B1(new_n321_), .B2(new_n410_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT95), .ZN(new_n460_));
  AND3_X1   g259(.A1(new_n407_), .A2(new_n408_), .A3(new_n395_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n388_), .B1(G169gat), .B2(G176gat), .ZN(new_n462_));
  INV_X1    g261(.A(G169gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n406_), .ZN(new_n464_));
  AOI22_X1  g263(.A1(new_n399_), .A2(new_n400_), .B1(new_n462_), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT94), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n394_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(G183gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(KEYINPUT25), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT25), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(G183gat), .ZN(new_n471_));
  INV_X1    g270(.A(G190gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT26), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT26), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(G190gat), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n469_), .A2(new_n471_), .A3(new_n473_), .A4(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n464_), .A2(KEYINPUT24), .A3(new_n395_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n466_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n461_), .B1(new_n467_), .B2(new_n479_), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT21), .B1(new_n302_), .B2(new_n304_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n481_), .B1(new_n297_), .B2(new_n299_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n309_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(KEYINPUT89), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n305_), .B1(new_n484_), .B2(new_n313_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n317_), .A2(new_n319_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n482_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n460_), .B1(new_n480_), .B2(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n476_), .A2(new_n466_), .A3(new_n477_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n394_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n409_), .B1(new_n491_), .B2(new_n478_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n321_), .A2(new_n492_), .A3(KEYINPUT95), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n459_), .B1(new_n488_), .B2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G226gat), .A2(G233gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n458_), .B1(new_n494_), .B2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT20), .ZN(new_n499_));
  AND2_X1   g298(.A1(new_n404_), .A2(new_n409_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n499_), .B1(new_n500_), .B2(new_n487_), .ZN(new_n501_));
  NOR3_X1   g300(.A1(new_n480_), .A2(new_n487_), .A3(new_n460_), .ZN(new_n502_));
  AOI21_X1  g301(.A(KEYINPUT95), .B1(new_n321_), .B2(new_n492_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n501_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n497_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n504_), .A2(KEYINPUT96), .A3(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n498_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n480_), .A2(new_n487_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n321_), .A2(new_n410_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n508_), .A2(new_n509_), .A3(KEYINPUT20), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n510_), .A2(new_n505_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n457_), .B1(new_n507_), .B2(new_n512_), .ZN(new_n513_));
  AOI211_X1 g312(.A(new_n511_), .B(new_n456_), .C1(new_n498_), .C2(new_n506_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n451_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT102), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  OAI211_X1 g316(.A(KEYINPUT102), .B(new_n451_), .C1(new_n513_), .C2(new_n514_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n507_), .A2(new_n512_), .A3(new_n457_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n508_), .A2(new_n509_), .A3(KEYINPUT20), .A4(new_n505_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n522_), .B1(new_n497_), .B2(new_n504_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n451_), .B1(new_n523_), .B2(new_n456_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n520_), .A2(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(KEYINPUT103), .B1(new_n519_), .B2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT103), .ZN(new_n527_));
  INV_X1    g326(.A(new_n525_), .ZN(new_n528_));
  AOI211_X1 g327(.A(new_n527_), .B(new_n528_), .C1(new_n517_), .C2(new_n518_), .ZN(new_n529_));
  OAI211_X1 g328(.A(new_n386_), .B(new_n450_), .C1(new_n526_), .C2(new_n529_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n513_), .A2(new_n514_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n444_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n532_), .A2(new_n430_), .A3(new_n442_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT33), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n534_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n440_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(KEYINPUT33), .B1(new_n435_), .B2(new_n445_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n446_), .A2(KEYINPUT33), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n531_), .A2(new_n538_), .A3(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT99), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n531_), .A2(new_n538_), .A3(new_n539_), .A4(KEYINPUT99), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n457_), .A2(KEYINPUT32), .ZN(new_n544_));
  OAI211_X1 g343(.A(new_n521_), .B(new_n544_), .C1(new_n494_), .C2(new_n505_), .ZN(new_n545_));
  OR2_X1    g344(.A1(new_n545_), .A2(KEYINPUT101), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(KEYINPUT101), .ZN(new_n547_));
  NOR3_X1   g346(.A1(new_n494_), .A2(new_n458_), .A3(new_n497_), .ZN(new_n548_));
  AOI21_X1  g347(.A(KEYINPUT96), .B1(new_n504_), .B2(new_n505_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n512_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  XOR2_X1   g349(.A(new_n544_), .B(KEYINPUT100), .Z(new_n551_));
  OAI211_X1 g350(.A(new_n546_), .B(new_n547_), .C1(new_n550_), .C2(new_n551_), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n448_), .A2(new_n552_), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n542_), .A2(new_n543_), .A3(new_n386_), .A4(new_n553_), .ZN(new_n554_));
  AOI211_X1 g353(.A(new_n528_), .B(new_n449_), .C1(new_n517_), .C2(new_n518_), .ZN(new_n555_));
  OAI211_X1 g354(.A(new_n554_), .B(new_n426_), .C1(new_n555_), .C2(new_n386_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n530_), .A2(new_n556_), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n289_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G231gat), .A2(G233gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n207_), .B(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(new_n272_), .ZN(new_n561_));
  XOR2_X1   g360(.A(G127gat), .B(G155gat), .Z(new_n562_));
  XNOR2_X1  g361(.A(G183gat), .B(G211gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(KEYINPUT81), .B(KEYINPUT16), .Z(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n561_), .A2(KEYINPUT17), .A3(new_n566_), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n567_), .B(KEYINPUT82), .Z(new_n568_));
  XNOR2_X1  g367(.A(new_n566_), .B(KEYINPUT17), .ZN(new_n569_));
  OR2_X1    g368(.A1(new_n561_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G190gat), .B(G218gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT75), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G134gat), .B(G162gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n576_), .A2(KEYINPUT36), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G232gat), .A2(G233gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT34), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(KEYINPUT35), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n580_), .A2(KEYINPUT35), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n582_), .B1(new_n232_), .B2(new_n282_), .ZN(new_n583_));
  OAI211_X1 g382(.A(new_n222_), .B(new_n276_), .C1(new_n229_), .C2(new_n231_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n581_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n583_), .A2(new_n581_), .A3(new_n584_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(KEYINPUT76), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT76), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n583_), .A2(new_n588_), .A3(new_n584_), .A4(new_n581_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n585_), .B1(new_n587_), .B2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n576_), .A2(KEYINPUT36), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n578_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n590_), .A2(KEYINPUT77), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n587_), .A2(new_n589_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n585_), .ZN(new_n596_));
  AOI221_X4 g395(.A(KEYINPUT77), .B1(new_n578_), .B2(new_n591_), .C1(new_n595_), .C2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n594_), .A2(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n571_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n558_), .A2(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(G1gat), .B1(new_n601_), .B2(new_n448_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n264_), .B(KEYINPUT74), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT78), .ZN(new_n604_));
  AOI21_X1  g403(.A(KEYINPUT37), .B1(new_n599_), .B2(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n592_), .A2(new_n593_), .ZN(new_n606_));
  OAI211_X1 g405(.A(new_n604_), .B(KEYINPUT37), .C1(new_n606_), .C2(new_n597_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n605_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n571_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n611_), .A2(new_n288_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n603_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT104), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n613_), .A2(new_n614_), .A3(new_n557_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n614_), .B1(new_n613_), .B2(new_n557_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n448_), .A2(G1gat), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT105), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT38), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n617_), .A2(KEYINPUT105), .A3(new_n618_), .ZN(new_n623_));
  AND3_X1   g422(.A1(new_n621_), .A2(new_n622_), .A3(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n622_), .B1(new_n621_), .B2(new_n623_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n602_), .B1(new_n624_), .B2(new_n625_), .ZN(G1324gat));
  NOR2_X1   g425(.A1(new_n526_), .A2(new_n529_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(new_n267_), .ZN(new_n628_));
  NOR3_X1   g427(.A1(new_n615_), .A2(new_n616_), .A3(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n627_), .ZN(new_n630_));
  OR3_X1    g429(.A1(new_n601_), .A2(KEYINPUT106), .A3(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(KEYINPUT106), .B1(new_n601_), .B2(new_n630_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n631_), .A2(G8gat), .A3(new_n632_), .ZN(new_n633_));
  OR2_X1    g432(.A1(new_n633_), .A2(KEYINPUT39), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(KEYINPUT39), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n629_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  XOR2_X1   g435(.A(KEYINPUT107), .B(KEYINPUT40), .Z(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(G1325gat));
  OAI21_X1  g437(.A(G15gat), .B1(new_n601_), .B2(new_n426_), .ZN(new_n639_));
  XOR2_X1   g438(.A(KEYINPUT108), .B(KEYINPUT41), .Z(new_n640_));
  XNOR2_X1  g439(.A(new_n639_), .B(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n613_), .A2(new_n557_), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n426_), .A2(G15gat), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n641_), .B1(new_n642_), .B2(new_n643_), .ZN(G1326gat));
  OAI21_X1  g443(.A(G22gat), .B1(new_n601_), .B2(new_n386_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT42), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n386_), .A2(G22gat), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n646_), .B1(new_n642_), .B2(new_n647_), .ZN(G1327gat));
  INV_X1    g447(.A(new_n599_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n610_), .A2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n558_), .A2(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT111), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(G29gat), .B1(new_n653_), .B2(new_n449_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n289_), .A2(new_n571_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n609_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n557_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT109), .ZN(new_n659_));
  AOI21_X1  g458(.A(KEYINPUT43), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n609_), .B1(new_n530_), .B2(new_n556_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT43), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n661_), .A2(KEYINPUT109), .A3(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n656_), .B1(new_n660_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT110), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT44), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n664_), .A2(new_n665_), .A3(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n386_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n550_), .A2(new_n456_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(new_n520_), .ZN(new_n670_));
  AOI21_X1  g469(.A(KEYINPUT102), .B1(new_n670_), .B2(new_n451_), .ZN(new_n671_));
  AOI211_X1 g470(.A(new_n516_), .B(KEYINPUT27), .C1(new_n669_), .C2(new_n520_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n525_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(new_n527_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n519_), .A2(KEYINPUT103), .A3(new_n525_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n668_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n668_), .B1(new_n673_), .B2(new_n449_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n426_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n386_), .B1(new_n448_), .B2(new_n552_), .ZN(new_n679_));
  AND3_X1   g478(.A1(new_n531_), .A2(new_n538_), .A3(new_n539_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n679_), .B1(new_n680_), .B2(KEYINPUT99), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n678_), .B1(new_n681_), .B2(new_n542_), .ZN(new_n682_));
  AOI22_X1  g481(.A1(new_n676_), .A2(new_n450_), .B1(new_n677_), .B2(new_n682_), .ZN(new_n683_));
  OAI211_X1 g482(.A(new_n659_), .B(KEYINPUT43), .C1(new_n683_), .C2(new_n609_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n662_), .B1(new_n661_), .B2(KEYINPUT109), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n655_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(KEYINPUT110), .B1(new_n686_), .B2(KEYINPUT44), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n667_), .A2(new_n687_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n664_), .A2(new_n666_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  AND3_X1   g489(.A1(new_n690_), .A2(G29gat), .A3(new_n449_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n654_), .B1(new_n688_), .B2(new_n691_), .ZN(G1328gat));
  INV_X1    g491(.A(G36gat), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n627_), .A2(new_n693_), .ZN(new_n694_));
  XOR2_X1   g493(.A(KEYINPUT113), .B(KEYINPUT45), .Z(new_n695_));
  OR3_X1    g494(.A1(new_n652_), .A2(new_n694_), .A3(new_n695_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n695_), .B1(new_n652_), .B2(new_n694_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT112), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n630_), .B1(new_n686_), .B2(KEYINPUT44), .ZN(new_n700_));
  AOI211_X1 g499(.A(new_n699_), .B(new_n693_), .C1(new_n688_), .C2(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n665_), .B1(new_n664_), .B2(new_n666_), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n686_), .A2(KEYINPUT110), .A3(KEYINPUT44), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n700_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(KEYINPUT112), .B1(new_n704_), .B2(G36gat), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n698_), .B1(new_n701_), .B2(new_n705_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(KEYINPUT114), .A2(KEYINPUT46), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  OAI221_X1 g507(.A(new_n698_), .B1(KEYINPUT114), .B2(KEYINPUT46), .C1(new_n701_), .C2(new_n705_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1329gat));
  AOI21_X1  g509(.A(G43gat), .B1(new_n653_), .B2(new_n678_), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n689_), .A2(new_n413_), .A3(new_n426_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n711_), .B1(new_n688_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT47), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n713_), .B(new_n714_), .ZN(G1330gat));
  AOI21_X1  g514(.A(G50gat), .B1(new_n653_), .B2(new_n668_), .ZN(new_n716_));
  AND3_X1   g515(.A1(new_n690_), .A2(G50gat), .A3(new_n668_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n716_), .B1(new_n688_), .B2(new_n717_), .ZN(G1331gat));
  INV_X1    g517(.A(new_n288_), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n603_), .A2(new_n683_), .A3(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(new_n600_), .ZN(new_n721_));
  OAI21_X1  g520(.A(G57gat), .B1(new_n721_), .B2(new_n448_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n264_), .A2(new_n288_), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n683_), .A2(new_n723_), .A3(new_n611_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n724_), .A2(new_n438_), .A3(new_n449_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n722_), .A2(new_n725_), .ZN(G1332gat));
  INV_X1    g525(.A(G64gat), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n724_), .A2(new_n727_), .A3(new_n627_), .ZN(new_n728_));
  OAI21_X1  g527(.A(G64gat), .B1(new_n721_), .B2(new_n630_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n729_), .A2(KEYINPUT48), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n729_), .A2(KEYINPUT48), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n728_), .B1(new_n730_), .B2(new_n731_), .ZN(G1333gat));
  INV_X1    g531(.A(G71gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n724_), .A2(new_n733_), .A3(new_n678_), .ZN(new_n734_));
  OAI21_X1  g533(.A(G71gat), .B1(new_n721_), .B2(new_n426_), .ZN(new_n735_));
  OR2_X1    g534(.A1(new_n735_), .A2(KEYINPUT116), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(KEYINPUT116), .ZN(new_n737_));
  XNOR2_X1  g536(.A(KEYINPUT115), .B(KEYINPUT49), .ZN(new_n738_));
  AND3_X1   g537(.A1(new_n736_), .A2(new_n737_), .A3(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n734_), .B1(new_n739_), .B2(new_n740_), .ZN(G1334gat));
  INV_X1    g540(.A(G78gat), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n724_), .A2(new_n742_), .A3(new_n668_), .ZN(new_n743_));
  OAI21_X1  g542(.A(G78gat), .B1(new_n721_), .B2(new_n386_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n744_), .A2(KEYINPUT50), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n744_), .A2(KEYINPUT50), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n743_), .B1(new_n745_), .B2(new_n746_), .ZN(G1335gat));
  AND2_X1   g546(.A1(new_n720_), .A2(new_n650_), .ZN(new_n748_));
  AOI21_X1  g547(.A(G85gat), .B1(new_n748_), .B2(new_n449_), .ZN(new_n749_));
  AOI211_X1 g548(.A(new_n610_), .B(new_n723_), .C1(new_n684_), .C2(new_n685_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n448_), .A2(new_n215_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n749_), .B1(new_n750_), .B2(new_n751_), .ZN(G1336gat));
  NAND3_X1  g551(.A1(new_n748_), .A2(new_n216_), .A3(new_n627_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n750_), .A2(new_n627_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n753_), .B1(new_n754_), .B2(new_n216_), .ZN(G1337gat));
  NAND3_X1  g554(.A1(new_n748_), .A2(new_n208_), .A3(new_n678_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT117), .ZN(new_n757_));
  INV_X1    g556(.A(G99gat), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n750_), .A2(new_n678_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n757_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT51), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT51), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n757_), .B(new_n762_), .C1(new_n758_), .C2(new_n759_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(G1338gat));
  NAND3_X1  g563(.A1(new_n748_), .A2(new_n209_), .A3(new_n668_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n750_), .A2(new_n668_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(G106gat), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n767_), .A2(KEYINPUT52), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n767_), .A2(KEYINPUT52), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n765_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g570(.A(KEYINPUT57), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT121), .ZN(new_n773_));
  INV_X1    g572(.A(new_n254_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n250_), .A2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n719_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n238_), .A2(new_n240_), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT119), .B1(new_n777_), .B2(new_n247_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT119), .ZN(new_n779_));
  AOI211_X1 g578(.A(new_n779_), .B(new_n242_), .C1(new_n238_), .C2(new_n240_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781_));
  OAI22_X1  g580(.A1(new_n778_), .A2(new_n780_), .B1(new_n781_), .B2(new_n243_), .ZN(new_n782_));
  XOR2_X1   g581(.A(KEYINPUT118), .B(KEYINPUT55), .Z(new_n783_));
  AND3_X1   g582(.A1(new_n245_), .A2(new_n249_), .A3(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT120), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n782_), .A2(new_n784_), .A3(new_n785_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n243_), .A2(new_n781_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n777_), .A2(new_n247_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n779_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n777_), .A2(KEYINPUT119), .A3(new_n247_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n787_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n245_), .A2(new_n249_), .A3(new_n783_), .ZN(new_n792_));
  AOI21_X1  g591(.A(KEYINPUT120), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n254_), .B1(new_n786_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT56), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n785_), .B1(new_n782_), .B2(new_n784_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n791_), .A2(KEYINPUT120), .A3(new_n792_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n799_), .A2(KEYINPUT56), .A3(new_n254_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n776_), .B1(new_n796_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n287_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n802_), .B1(new_n283_), .B2(new_n279_), .ZN(new_n803_));
  OR2_X1    g602(.A1(new_n277_), .A2(new_n279_), .ZN(new_n804_));
  AOI22_X1  g603(.A1(new_n284_), .A2(new_n802_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n259_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n649_), .B(new_n773_), .C1(new_n801_), .C2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n796_), .A2(new_n800_), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n775_), .A2(new_n805_), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT58), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT56), .B1(new_n799_), .B2(new_n254_), .ZN(new_n812_));
  AOI211_X1 g611(.A(new_n795_), .B(new_n774_), .C1(new_n797_), .C2(new_n798_), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n810_), .B(KEYINPUT58), .C1(new_n812_), .C2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n657_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n808_), .B1(new_n811_), .B2(new_n815_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n812_), .A2(new_n813_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n806_), .B1(new_n817_), .B2(new_n776_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n773_), .B1(new_n818_), .B2(new_n649_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n571_), .B1(new_n816_), .B2(new_n819_), .ZN(new_n820_));
  NOR3_X1   g619(.A1(new_n611_), .A2(new_n264_), .A3(new_n719_), .ZN(new_n821_));
  XOR2_X1   g620(.A(new_n821_), .B(KEYINPUT54), .Z(new_n822_));
  NAND2_X1  g621(.A1(new_n820_), .A2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n676_), .A2(new_n449_), .A3(new_n678_), .ZN(new_n824_));
  XOR2_X1   g623(.A(new_n824_), .B(KEYINPUT122), .Z(new_n825_));
  AND2_X1   g624(.A1(new_n823_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(G113gat), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(new_n827_), .A3(new_n719_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(KEYINPUT59), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n823_), .A2(new_n825_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT59), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n288_), .B1(new_n829_), .B2(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n828_), .B1(new_n833_), .B2(new_n827_), .ZN(G1340gat));
  INV_X1    g633(.A(KEYINPUT60), .ZN(new_n835_));
  INV_X1    g634(.A(G120gat), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n264_), .A2(new_n835_), .A3(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n837_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n826_), .A2(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n603_), .B1(new_n829_), .B2(new_n832_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n839_), .B1(new_n840_), .B2(new_n836_), .ZN(G1341gat));
  AOI21_X1  g640(.A(G127gat), .B1(new_n826_), .B2(new_n610_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n829_), .A2(new_n832_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT123), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n610_), .A2(new_n844_), .A3(G127gat), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n845_), .B1(new_n844_), .B2(G127gat), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n842_), .B1(new_n843_), .B2(new_n846_), .ZN(G1342gat));
  INV_X1    g646(.A(G134gat), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n826_), .A2(new_n848_), .A3(new_n599_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n609_), .B1(new_n829_), .B2(new_n832_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n849_), .B1(new_n850_), .B2(new_n848_), .ZN(G1343gat));
  NOR2_X1   g650(.A1(new_n678_), .A2(new_n386_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n853_), .B1(new_n820_), .B2(new_n822_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n627_), .A2(new_n448_), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n719_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g657(.A(new_n603_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n856_), .A2(new_n859_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(G148gat), .ZN(G1345gat));
  NAND4_X1  g660(.A1(new_n823_), .A2(new_n610_), .A3(new_n852_), .A4(new_n855_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT124), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT124), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n854_), .A2(new_n864_), .A3(new_n610_), .A4(new_n855_), .ZN(new_n865_));
  XOR2_X1   g664(.A(KEYINPUT61), .B(G155gat), .Z(new_n866_));
  AND3_X1   g665(.A1(new_n863_), .A2(new_n865_), .A3(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n866_), .B1(new_n863_), .B2(new_n865_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n867_), .A2(new_n868_), .ZN(G1346gat));
  INV_X1    g668(.A(G162gat), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n856_), .A2(new_n870_), .A3(new_n599_), .ZN(new_n871_));
  AND2_X1   g670(.A1(new_n856_), .A2(new_n657_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n871_), .B1(new_n872_), .B2(new_n870_), .ZN(G1347gat));
  INV_X1    g672(.A(KEYINPUT62), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n627_), .A2(new_n386_), .A3(new_n450_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n875_), .B1(new_n820_), .B2(new_n822_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n719_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n874_), .B1(new_n877_), .B2(G169gat), .ZN(new_n878_));
  AOI211_X1 g677(.A(KEYINPUT62), .B(new_n463_), .C1(new_n876_), .C2(new_n719_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n875_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n823_), .A2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n719_), .A2(new_n405_), .ZN(new_n882_));
  XOR2_X1   g681(.A(new_n882_), .B(KEYINPUT125), .Z(new_n883_));
  OAI22_X1  g682(.A1(new_n878_), .A2(new_n879_), .B1(new_n881_), .B2(new_n883_), .ZN(G1348gat));
  OAI21_X1  g683(.A(G176gat), .B1(new_n881_), .B2(new_n603_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n876_), .A2(new_n406_), .A3(new_n264_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(G1349gat));
  OAI21_X1  g686(.A(G183gat), .B1(new_n881_), .B2(new_n571_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT126), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n876_), .A2(new_n610_), .A3(new_n399_), .ZN(new_n890_));
  AND3_X1   g689(.A1(new_n888_), .A2(new_n889_), .A3(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n889_), .B1(new_n888_), .B2(new_n890_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n891_), .A2(new_n892_), .ZN(G1350gat));
  OAI21_X1  g692(.A(G190gat), .B1(new_n881_), .B2(new_n609_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n876_), .A2(new_n599_), .A3(new_n400_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1351gat));
  NOR2_X1   g695(.A1(new_n630_), .A2(new_n449_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n854_), .A2(new_n719_), .A3(new_n897_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g698(.A1(new_n854_), .A2(new_n859_), .A3(new_n897_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(G204gat), .ZN(G1353gat));
  NAND3_X1  g700(.A1(new_n854_), .A2(new_n610_), .A3(new_n897_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT63), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n301_), .ZN(new_n905_));
  OAI21_X1  g704(.A(KEYINPUT127), .B1(new_n903_), .B2(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT127), .ZN(new_n907_));
  NAND4_X1  g706(.A1(new_n902_), .A2(new_n907_), .A3(new_n904_), .A4(new_n301_), .ZN(new_n908_));
  XOR2_X1   g707(.A(KEYINPUT63), .B(G211gat), .Z(new_n909_));
  AOI22_X1  g708(.A1(new_n906_), .A2(new_n908_), .B1(new_n903_), .B2(new_n909_), .ZN(G1354gat));
  NAND4_X1  g709(.A1(new_n854_), .A2(new_n303_), .A3(new_n599_), .A4(new_n897_), .ZN(new_n911_));
  AND3_X1   g710(.A1(new_n854_), .A2(new_n657_), .A3(new_n897_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n911_), .B1(new_n912_), .B2(new_n303_), .ZN(G1355gat));
endmodule


