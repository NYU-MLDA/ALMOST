//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 0 1 1 0 0 1 1 1 0 0 1 0 1 1 1 0 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 0 1 0 1 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n710_, new_n711_, new_n712_, new_n713_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n826_, new_n827_, new_n828_, new_n830_, new_n831_,
    new_n832_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n850_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n927_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(G183gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT25), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT25), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G183gat), .ZN(new_n206_));
  INV_X1    g005(.A(G190gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT26), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT26), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G190gat), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n204_), .A2(new_n206_), .A3(new_n208_), .A4(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT24), .ZN(new_n212_));
  INV_X1    g011(.A(G169gat), .ZN(new_n213_));
  INV_X1    g012(.A(G176gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n212_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n214_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n216_), .A2(KEYINPUT24), .A3(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT23), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(G183gat), .A3(G190gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n211_), .A2(new_n215_), .A3(new_n218_), .A4(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n219_), .A2(new_n221_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n203_), .A2(new_n207_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  OR3_X1    g027(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n229_));
  OAI21_X1  g028(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n228_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n224_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT79), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT79), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n224_), .A2(new_n234_), .A3(new_n231_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G71gat), .B(G99gat), .ZN(new_n237_));
  INV_X1    g036(.A(G43gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n236_), .B(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G227gat), .A2(G233gat), .ZN(new_n243_));
  INV_X1    g042(.A(G15gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT30), .ZN(new_n246_));
  XOR2_X1   g045(.A(G127gat), .B(G134gat), .Z(new_n247_));
  INV_X1    g046(.A(G120gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(G113gat), .ZN(new_n249_));
  INV_X1    g048(.A(G113gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(G120gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n249_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n247_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G127gat), .B(G134gat), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n254_), .A2(new_n249_), .A3(new_n251_), .ZN(new_n255_));
  AND2_X1   g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n246_), .B(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n242_), .B(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G1gat), .B(G29gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(G85gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT0), .B(G57gat), .ZN(new_n262_));
  XOR2_X1   g061(.A(new_n261_), .B(new_n262_), .Z(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G155gat), .A2(G162gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(KEYINPUT1), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(KEYINPUT81), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT81), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n265_), .A2(new_n268_), .A3(KEYINPUT1), .ZN(new_n269_));
  INV_X1    g068(.A(G155gat), .ZN(new_n270_));
  INV_X1    g069(.A(G162gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT1), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n273_), .A2(G155gat), .A3(G162gat), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n267_), .A2(new_n269_), .A3(new_n272_), .A4(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G141gat), .A2(G148gat), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(G141gat), .A2(G148gat), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n275_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT3), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n278_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT2), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n276_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n285_));
  OAI21_X1  g084(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n282_), .A2(new_n284_), .A3(new_n285_), .A4(new_n286_), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n272_), .A2(new_n265_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n280_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT4), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n290_), .A2(new_n291_), .A3(new_n256_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G225gat), .A2(G233gat), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n279_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n274_), .A2(new_n272_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n268_), .B1(new_n265_), .B2(KEYINPUT1), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n296_), .B1(new_n299_), .B2(new_n269_), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n287_), .A2(new_n288_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n256_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT91), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n253_), .A2(new_n255_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n280_), .A2(new_n304_), .A3(new_n289_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n302_), .A2(new_n303_), .A3(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n290_), .A2(KEYINPUT91), .A3(new_n256_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n295_), .B1(new_n308_), .B2(KEYINPUT4), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n294_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n264_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n308_), .A2(new_n293_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n291_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n312_), .B(new_n263_), .C1(new_n313_), .C2(new_n295_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n311_), .A2(KEYINPUT95), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT95), .ZN(new_n316_));
  OAI211_X1 g115(.A(new_n316_), .B(new_n264_), .C1(new_n309_), .C2(new_n310_), .ZN(new_n317_));
  INV_X1    g116(.A(G218gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(G211gat), .ZN(new_n319_));
  INV_X1    g118(.A(G211gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(G218gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(G197gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(G204gat), .ZN(new_n324_));
  INV_X1    g123(.A(G204gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(G197gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n324_), .A2(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n322_), .B1(KEYINPUT21), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT84), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n329_), .B1(new_n325_), .B2(G197gat), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n323_), .A2(KEYINPUT84), .A3(G204gat), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT21), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n330_), .A2(new_n331_), .A3(new_n332_), .A4(new_n326_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n328_), .A2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n330_), .A2(new_n331_), .A3(new_n326_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n332_), .B1(new_n319_), .B2(new_n321_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT85), .ZN(new_n337_));
  AND3_X1   g136(.A1(new_n335_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n337_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n334_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  AND3_X1   g139(.A1(new_n224_), .A2(new_n234_), .A3(new_n231_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n234_), .B1(new_n224_), .B2(new_n231_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n340_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n335_), .A2(new_n336_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT85), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n335_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n346_));
  AOI22_X1  g145(.A1(new_n345_), .A2(new_n346_), .B1(new_n333_), .B2(new_n328_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT22), .B(G169gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(new_n214_), .ZN(new_n349_));
  AND2_X1   g148(.A1(new_n217_), .A2(KEYINPUT90), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n217_), .A2(KEYINPUT90), .ZN(new_n351_));
  OAI211_X1 g150(.A(new_n349_), .B(new_n228_), .C1(new_n350_), .C2(new_n351_), .ZN(new_n352_));
  AND2_X1   g151(.A1(new_n352_), .A2(new_n224_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n347_), .A2(new_n353_), .ZN(new_n354_));
  XOR2_X1   g153(.A(KEYINPUT94), .B(KEYINPUT20), .Z(new_n355_));
  NAND3_X1  g154(.A1(new_n343_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G226gat), .A2(G233gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT88), .ZN(new_n358_));
  XOR2_X1   g157(.A(KEYINPUT87), .B(KEYINPUT19), .Z(new_n359_));
  OR2_X1    g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n359_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n356_), .A2(new_n362_), .ZN(new_n363_));
  XOR2_X1   g162(.A(G8gat), .B(G36gat), .Z(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT18), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G64gat), .B(G92gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n367_), .A2(KEYINPUT32), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n347_), .A2(new_n233_), .A3(new_n235_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT89), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n362_), .A2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n360_), .A2(KEYINPUT89), .A3(new_n361_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n352_), .A2(new_n224_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n340_), .A2(new_n374_), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n369_), .A2(new_n373_), .A3(KEYINPUT20), .A4(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n363_), .A2(new_n368_), .A3(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT93), .ZN(new_n378_));
  INV_X1    g177(.A(new_n373_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n369_), .A2(KEYINPUT20), .A3(new_n375_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n360_), .A2(KEYINPUT20), .A3(new_n361_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n381_), .B1(new_n236_), .B2(new_n340_), .ZN(new_n382_));
  AOI22_X1  g181(.A1(new_n379_), .A2(new_n380_), .B1(new_n382_), .B2(new_n354_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n377_), .B1(new_n378_), .B2(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n368_), .B1(new_n383_), .B2(KEYINPUT93), .ZN(new_n385_));
  OAI211_X1 g184(.A(new_n315_), .B(new_n317_), .C1(new_n384_), .C2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n380_), .A2(new_n379_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n382_), .A2(new_n354_), .ZN(new_n388_));
  AND3_X1   g187(.A1(new_n387_), .A2(new_n367_), .A3(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n367_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n309_), .A2(new_n310_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT92), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT33), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n392_), .A2(new_n263_), .A3(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n314_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n263_), .B1(new_n308_), .B2(new_n294_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n292_), .A2(new_n293_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n398_), .B1(new_n313_), .B2(new_n399_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n391_), .A2(new_n396_), .A3(new_n397_), .A4(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n386_), .A2(new_n401_), .ZN(new_n402_));
  AOI22_X1  g201(.A1(new_n340_), .A2(KEYINPUT83), .B1(G228gat), .B2(G233gat), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n300_), .A2(new_n301_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT29), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n340_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  XOR2_X1   g205(.A(new_n403_), .B(new_n406_), .Z(new_n407_));
  XOR2_X1   g206(.A(G22gat), .B(G50gat), .Z(new_n408_));
  OR3_X1    g207(.A1(new_n290_), .A2(KEYINPUT29), .A3(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n408_), .B1(new_n290_), .B2(KEYINPUT29), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(KEYINPUT82), .B(KEYINPUT28), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G78gat), .B(G106gat), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  OR2_X1    g214(.A1(new_n415_), .A2(KEYINPUT86), .ZN(new_n416_));
  INV_X1    g215(.A(new_n412_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n409_), .A2(new_n417_), .A3(new_n410_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n413_), .A2(new_n416_), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n415_), .B1(new_n413_), .B2(new_n418_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n407_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n421_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n407_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n423_), .A2(new_n424_), .A3(new_n419_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n422_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n402_), .A2(KEYINPUT96), .A3(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n391_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT27), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n387_), .A2(new_n388_), .A3(new_n367_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(KEYINPUT99), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT99), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n383_), .A2(new_n434_), .A3(new_n367_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n363_), .A2(new_n376_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n367_), .B(KEYINPUT98), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n430_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n436_), .A2(KEYINPUT100), .A3(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(KEYINPUT100), .B1(new_n436_), .B2(new_n439_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n431_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n315_), .A2(new_n317_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT97), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n315_), .A2(KEYINPUT97), .A3(new_n317_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n446_), .A2(new_n426_), .A3(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n428_), .B1(new_n443_), .B2(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(KEYINPUT96), .B1(new_n402_), .B2(new_n427_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n259_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT101), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n446_), .A2(new_n447_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n454_), .A2(new_n259_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n436_), .A2(new_n439_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT100), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  AOI22_X1  g257(.A1(new_n458_), .A2(new_n440_), .B1(new_n430_), .B2(new_n429_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n455_), .A2(new_n427_), .A3(new_n459_), .ZN(new_n460_));
  OAI211_X1 g259(.A(KEYINPUT101), .B(new_n259_), .C1(new_n449_), .C2(new_n450_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n453_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT73), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G99gat), .A2(G106gat), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT6), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT65), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n464_), .B(KEYINPUT6), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT65), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  AND2_X1   g269(.A1(new_n467_), .A2(new_n470_), .ZN(new_n471_));
  XOR2_X1   g270(.A(KEYINPUT10), .B(G99gat), .Z(new_n472_));
  INV_X1    g271(.A(G106gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  XOR2_X1   g273(.A(G85gat), .B(G92gat), .Z(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT9), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT9), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n477_), .A2(G85gat), .A3(G92gat), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n474_), .A2(new_n476_), .A3(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n471_), .A2(new_n479_), .A3(KEYINPUT66), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT66), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n467_), .A2(new_n470_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n474_), .A2(new_n476_), .A3(new_n478_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n481_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n480_), .A2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G29gat), .B(G36gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G43gat), .B(G50gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(G99gat), .A2(G106gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT7), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n467_), .A2(new_n470_), .A3(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT8), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n475_), .B(KEYINPUT67), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n491_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  AND2_X1   g293(.A1(new_n490_), .A2(new_n468_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G85gat), .B(G92gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT67), .ZN(new_n497_));
  OAI21_X1  g296(.A(KEYINPUT8), .B1(new_n495_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n494_), .A2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n485_), .A2(new_n488_), .A3(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G232gat), .A2(G233gat), .ZN(new_n501_));
  XOR2_X1   g300(.A(new_n501_), .B(KEYINPUT34), .Z(new_n502_));
  INV_X1    g301(.A(KEYINPUT35), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(KEYINPUT72), .B(KEYINPUT15), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n488_), .B(new_n505_), .ZN(new_n506_));
  AOI22_X1  g305(.A1(new_n480_), .A2(new_n484_), .B1(new_n494_), .B2(new_n498_), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n500_), .B(new_n504_), .C1(new_n506_), .C2(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n463_), .B1(new_n508_), .B2(KEYINPUT75), .ZN(new_n509_));
  OR2_X1    g308(.A1(new_n507_), .A2(new_n506_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n510_), .A2(KEYINPUT73), .A3(new_n500_), .A4(new_n504_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n502_), .A2(new_n503_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n509_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n513_));
  OAI221_X1 g312(.A(new_n463_), .B1(new_n503_), .B2(new_n502_), .C1(new_n508_), .C2(KEYINPUT75), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT74), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT36), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G190gat), .B(G218gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G134gat), .B(G162gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n517_), .A2(new_n518_), .A3(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(KEYINPUT74), .B1(new_n513_), .B2(new_n514_), .ZN(new_n524_));
  OAI21_X1  g323(.A(KEYINPUT36), .B1(new_n524_), .B2(new_n521_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n515_), .A2(new_n521_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n523_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  AND2_X1   g327(.A1(new_n462_), .A2(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G113gat), .B(G141gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G169gat), .B(G197gat), .ZN(new_n531_));
  XOR2_X1   g330(.A(new_n530_), .B(new_n531_), .Z(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G15gat), .B(G22gat), .ZN(new_n534_));
  INV_X1    g333(.A(G8gat), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G1gat), .B(G8gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(new_n539_), .B(new_n488_), .Z(new_n540_));
  NAND2_X1  g339(.A1(G229gat), .A2(G233gat), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n539_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n506_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n488_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(new_n541_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n543_), .B1(new_n545_), .B2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT77), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(KEYINPUT78), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n549_), .A2(KEYINPUT78), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n533_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n552_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n554_), .A2(new_n550_), .A3(new_n532_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  XOR2_X1   g355(.A(G176gat), .B(G204gat), .Z(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT70), .ZN(new_n558_));
  XOR2_X1   g357(.A(G120gat), .B(G148gat), .Z(new_n559_));
  XOR2_X1   g358(.A(new_n558_), .B(new_n559_), .Z(new_n560_));
  XNOR2_X1  g359(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n562_), .B(KEYINPUT71), .Z(new_n563_));
  NAND2_X1  g362(.A1(new_n485_), .A2(new_n499_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G57gat), .B(G64gat), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n565_), .A2(KEYINPUT11), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(KEYINPUT11), .ZN(new_n567_));
  XOR2_X1   g366(.A(G71gat), .B(G78gat), .Z(new_n568_));
  NAND3_X1  g367(.A1(new_n566_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n569_));
  OR2_X1    g368(.A1(new_n567_), .A2(new_n568_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n564_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n507_), .A2(new_n571_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n573_), .A2(KEYINPUT68), .A3(new_n574_), .ZN(new_n575_));
  OR3_X1    g374(.A1(new_n564_), .A2(KEYINPUT68), .A3(new_n572_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G230gat), .A2(G233gat), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n577_), .B(KEYINPUT64), .Z(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  AND3_X1   g378(.A1(new_n575_), .A2(new_n576_), .A3(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n573_), .A2(KEYINPUT12), .A3(new_n574_), .ZN(new_n581_));
  OR3_X1    g380(.A1(new_n507_), .A2(KEYINPUT12), .A3(new_n571_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n579_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n563_), .B1(new_n580_), .B2(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n580_), .A2(new_n583_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(new_n562_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT13), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n584_), .A2(new_n586_), .A3(KEYINPUT13), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G231gat), .A2(G233gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n539_), .B(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(new_n572_), .ZN(new_n595_));
  XOR2_X1   g394(.A(G127gat), .B(G155gat), .Z(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT16), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G183gat), .B(G211gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT17), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  AND2_X1   g400(.A1(new_n599_), .A2(new_n600_), .ZN(new_n602_));
  NOR3_X1   g401(.A1(new_n595_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n603_), .B1(new_n601_), .B2(new_n595_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT76), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n603_), .A2(KEYINPUT76), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n529_), .A2(new_n556_), .A3(new_n592_), .A4(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT103), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n202_), .B1(new_n612_), .B2(new_n454_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT38), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n462_), .A2(new_n556_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT37), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n527_), .A2(new_n616_), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n523_), .A2(new_n525_), .A3(KEYINPUT37), .A4(new_n526_), .ZN(new_n618_));
  AOI211_X1 g417(.A(new_n608_), .B(new_n591_), .C1(new_n617_), .C2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n615_), .A2(new_n619_), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n620_), .B(KEYINPUT102), .Z(new_n621_));
  NAND3_X1  g420(.A1(new_n621_), .A2(new_n202_), .A3(new_n454_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n613_), .B1(new_n614_), .B2(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n623_), .B1(new_n614_), .B2(new_n622_), .ZN(G1324gat));
  OAI21_X1  g423(.A(G8gat), .B1(new_n610_), .B2(new_n459_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT39), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n621_), .A2(new_n535_), .A3(new_n443_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n628_), .B(KEYINPUT40), .Z(G1325gat));
  XNOR2_X1  g428(.A(new_n610_), .B(KEYINPUT103), .ZN(new_n630_));
  OAI21_X1  g429(.A(G15gat), .B1(new_n630_), .B2(new_n259_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(KEYINPUT104), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT104), .ZN(new_n633_));
  OAI211_X1 g432(.A(new_n633_), .B(G15gat), .C1(new_n630_), .C2(new_n259_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT41), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n621_), .A2(new_n244_), .A3(new_n258_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n632_), .A2(new_n634_), .A3(KEYINPUT41), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n637_), .A2(new_n638_), .A3(new_n639_), .ZN(G1326gat));
  OAI21_X1  g439(.A(G22gat), .B1(new_n630_), .B2(new_n427_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT42), .ZN(new_n642_));
  INV_X1    g441(.A(G22gat), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n621_), .A2(new_n643_), .A3(new_n426_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n644_), .ZN(G1327gat));
  NAND2_X1  g444(.A1(new_n527_), .A2(new_n608_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n646_), .A2(new_n591_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n615_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(G29gat), .B1(new_n649_), .B2(new_n454_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT106), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT43), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n617_), .A2(new_n618_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n461_), .A2(new_n460_), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n446_), .A2(new_n426_), .A3(new_n447_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n459_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n402_), .A2(new_n427_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT96), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n656_), .A2(new_n659_), .A3(new_n428_), .ZN(new_n660_));
  AOI21_X1  g459(.A(KEYINPUT101), .B1(new_n660_), .B2(new_n259_), .ZN(new_n661_));
  OAI211_X1 g460(.A(new_n652_), .B(new_n653_), .C1(new_n654_), .C2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT105), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n462_), .A2(KEYINPUT105), .A3(new_n652_), .A4(new_n653_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n653_), .B1(new_n654_), .B2(new_n661_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(KEYINPUT43), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n664_), .A2(new_n665_), .A3(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n556_), .ZN(new_n669_));
  NOR3_X1   g468(.A1(new_n591_), .A2(new_n609_), .A3(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT44), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n651_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  AOI211_X1 g472(.A(KEYINPUT106), .B(KEYINPUT44), .C1(new_n668_), .C2(new_n670_), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n668_), .A2(KEYINPUT44), .A3(new_n670_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n454_), .A2(G29gat), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n650_), .B1(new_n677_), .B2(new_n678_), .ZN(G1328gat));
  OAI211_X1 g478(.A(new_n676_), .B(new_n443_), .C1(new_n673_), .C2(new_n674_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(G36gat), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n648_), .A2(G36gat), .A3(new_n459_), .ZN(new_n682_));
  XOR2_X1   g481(.A(new_n682_), .B(KEYINPUT45), .Z(new_n683_));
  NAND2_X1  g482(.A1(new_n681_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT46), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n681_), .A2(KEYINPUT46), .A3(new_n683_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(G1329gat));
  NOR2_X1   g487(.A1(new_n259_), .A2(new_n238_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n675_), .A2(new_n676_), .A3(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n238_), .B1(new_n648_), .B2(new_n259_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n692_));
  AND3_X1   g491(.A1(new_n690_), .A2(new_n691_), .A3(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n692_), .B1(new_n690_), .B2(new_n691_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n693_), .A2(new_n694_), .ZN(G1330gat));
  AOI21_X1  g494(.A(G50gat), .B1(new_n649_), .B2(new_n426_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n426_), .A2(G50gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n696_), .B1(new_n677_), .B2(new_n697_), .ZN(G1331gat));
  NOR3_X1   g497(.A1(new_n592_), .A2(new_n556_), .A3(new_n608_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n529_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n454_), .ZN(new_n701_));
  OAI21_X1  g500(.A(G57gat), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n617_), .A2(new_n618_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n703_), .A2(new_n591_), .A3(new_n609_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT108), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n462_), .A2(new_n669_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  OR2_X1    g506(.A1(new_n701_), .A2(G57gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n702_), .B1(new_n707_), .B2(new_n708_), .ZN(G1332gat));
  OAI21_X1  g508(.A(G64gat), .B1(new_n700_), .B2(new_n459_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT48), .ZN(new_n711_));
  OR2_X1    g510(.A1(new_n459_), .A2(G64gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n711_), .B1(new_n707_), .B2(new_n712_), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n713_), .B(KEYINPUT109), .Z(G1333gat));
  OAI21_X1  g513(.A(G71gat), .B1(new_n700_), .B2(new_n259_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT49), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n259_), .A2(G71gat), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT110), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n716_), .B1(new_n707_), .B2(new_n718_), .ZN(G1334gat));
  OAI21_X1  g518(.A(G78gat), .B1(new_n700_), .B2(new_n427_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT50), .ZN(new_n721_));
  OR2_X1    g520(.A1(new_n427_), .A2(G78gat), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n721_), .B1(new_n707_), .B2(new_n722_), .ZN(G1335gat));
  NOR3_X1   g522(.A1(new_n592_), .A2(new_n556_), .A3(new_n609_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n668_), .A2(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(G85gat), .B1(new_n725_), .B2(new_n701_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n592_), .A2(new_n646_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n706_), .A2(new_n727_), .ZN(new_n728_));
  OR2_X1    g527(.A1(new_n701_), .A2(G85gat), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n726_), .B1(new_n728_), .B2(new_n729_), .ZN(G1336gat));
  OAI21_X1  g529(.A(G92gat), .B1(new_n725_), .B2(new_n459_), .ZN(new_n731_));
  OR2_X1    g530(.A1(new_n459_), .A2(G92gat), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n731_), .B1(new_n728_), .B2(new_n732_), .ZN(G1337gat));
  OAI21_X1  g532(.A(G99gat), .B1(new_n725_), .B2(new_n259_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n728_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n735_), .A2(new_n258_), .A3(new_n472_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g537(.A(KEYINPUT112), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n668_), .A2(new_n426_), .A3(new_n724_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n740_), .A2(KEYINPUT111), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT111), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n668_), .A2(new_n742_), .A3(new_n426_), .A4(new_n724_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(G106gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n739_), .B1(new_n741_), .B2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n740_), .A2(KEYINPUT111), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n746_), .A2(KEYINPUT112), .A3(G106gat), .A4(new_n743_), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n745_), .A2(KEYINPUT52), .A3(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT52), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n739_), .B(new_n749_), .C1(new_n741_), .C2(new_n744_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n735_), .A2(new_n473_), .A3(new_n426_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(KEYINPUT53), .B1(new_n748_), .B2(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n745_), .A2(KEYINPUT52), .A3(new_n747_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT53), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n754_), .A2(new_n755_), .A3(new_n750_), .A4(new_n751_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n753_), .A2(new_n756_), .ZN(G1339gat));
  NAND2_X1  g556(.A1(new_n556_), .A2(new_n586_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n581_), .A2(new_n579_), .A3(new_n582_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n583_), .B1(KEYINPUT55), .B2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n581_), .A2(new_n582_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n761_), .A2(KEYINPUT55), .A3(new_n578_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n563_), .B1(new_n760_), .B2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT56), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n759_), .A2(KEYINPUT55), .ZN(new_n767_));
  INV_X1    g566(.A(new_n583_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(new_n762_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n770_), .A2(KEYINPUT56), .A3(new_n563_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n758_), .B1(new_n766_), .B2(new_n771_), .ZN(new_n772_));
  AOI211_X1 g571(.A(new_n541_), .B(new_n545_), .C1(new_n544_), .C2(new_n488_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n540_), .A2(new_n541_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n533_), .B1(new_n773_), .B2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n548_), .A2(new_n532_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n587_), .A2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n528_), .B(KEYINPUT57), .C1(new_n772_), .C2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT115), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n766_), .A2(new_n771_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n783_), .A2(new_n556_), .A3(new_n586_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n527_), .B1(new_n784_), .B2(new_n779_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT115), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n785_), .A2(new_n786_), .A3(KEYINPUT57), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n782_), .A2(new_n787_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n586_), .A2(new_n778_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n783_), .A2(KEYINPUT58), .A3(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(KEYINPUT58), .B1(new_n783_), .B2(new_n789_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n528_), .B1(new_n772_), .B2(new_n780_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT57), .ZN(new_n795_));
  AOI22_X1  g594(.A1(new_n793_), .A2(new_n653_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n788_), .A2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n608_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n703_), .A2(new_n669_), .A3(new_n592_), .A4(new_n609_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT113), .ZN(new_n800_));
  OAI21_X1  g599(.A(KEYINPUT114), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT54), .B1(new_n799_), .B2(new_n800_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT114), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n619_), .A2(KEYINPUT113), .A3(new_n803_), .A4(new_n669_), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n801_), .A2(new_n802_), .A3(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n802_), .B1(new_n804_), .B2(new_n801_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n798_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  NOR4_X1   g606(.A1(new_n443_), .A2(new_n701_), .A3(new_n259_), .A4(new_n426_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n810_), .A2(new_n250_), .A3(new_n556_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n792_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n653_), .A2(new_n812_), .A3(new_n790_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n794_), .A2(new_n795_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(KEYINPUT116), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT116), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n813_), .A2(new_n814_), .A3(new_n817_), .ZN(new_n818_));
  AND3_X1   g617(.A1(new_n816_), .A2(new_n788_), .A3(new_n818_), .ZN(new_n819_));
  OAI22_X1  g618(.A1(new_n819_), .A2(new_n609_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT59), .ZN(new_n821_));
  AND2_X1   g620(.A1(new_n808_), .A2(new_n821_), .ZN(new_n822_));
  AOI22_X1  g621(.A1(KEYINPUT59), .A2(new_n809_), .B1(new_n820_), .B2(new_n822_), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n823_), .A2(new_n556_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n811_), .B1(new_n824_), .B2(new_n250_), .ZN(G1340gat));
  OAI21_X1  g624(.A(new_n248_), .B1(new_n592_), .B2(KEYINPUT60), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n810_), .B(new_n826_), .C1(KEYINPUT60), .C2(new_n248_), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n823_), .A2(new_n591_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n827_), .B1(new_n828_), .B2(new_n248_), .ZN(G1341gat));
  INV_X1    g628(.A(G127gat), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n810_), .A2(new_n830_), .A3(new_n609_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n823_), .A2(new_n609_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n831_), .B1(new_n832_), .B2(new_n830_), .ZN(G1342gat));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n834_));
  INV_X1    g633(.A(G134gat), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n835_), .B1(new_n823_), .B2(new_n653_), .ZN(new_n836_));
  NOR3_X1   g635(.A1(new_n809_), .A2(G134gat), .A3(new_n528_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n834_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n837_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n809_), .A2(KEYINPUT59), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n820_), .A2(new_n822_), .ZN(new_n841_));
  AND3_X1   g640(.A1(new_n840_), .A2(new_n653_), .A3(new_n841_), .ZN(new_n842_));
  OAI211_X1 g641(.A(KEYINPUT117), .B(new_n839_), .C1(new_n842_), .C2(new_n835_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n838_), .A2(new_n843_), .ZN(G1343gat));
  NOR4_X1   g643(.A1(new_n443_), .A2(new_n701_), .A3(new_n258_), .A4(new_n427_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n807_), .A2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n556_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n848_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g648(.A1(new_n847_), .A2(new_n591_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g650(.A1(new_n846_), .A2(new_n608_), .ZN(new_n852_));
  XOR2_X1   g651(.A(KEYINPUT61), .B(G155gat), .Z(new_n853_));
  XNOR2_X1  g652(.A(new_n852_), .B(new_n853_), .ZN(G1346gat));
  NOR3_X1   g653(.A1(new_n846_), .A2(G162gat), .A3(new_n528_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n847_), .A2(new_n653_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n855_), .B1(G162gat), .B2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT118), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n857_), .B(new_n858_), .ZN(G1347gat));
  NAND2_X1  g658(.A1(new_n455_), .A2(new_n443_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n860_), .A2(new_n669_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(KEYINPUT119), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n862_), .A2(new_n426_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n213_), .B1(new_n820_), .B2(new_n863_), .ZN(new_n864_));
  XOR2_X1   g663(.A(new_n864_), .B(KEYINPUT62), .Z(new_n865_));
  NOR2_X1   g664(.A1(new_n860_), .A2(new_n426_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n820_), .A2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n868_), .A2(new_n348_), .A3(new_n556_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n865_), .A2(new_n869_), .ZN(G1348gat));
  AOI21_X1  g669(.A(new_n609_), .B1(new_n788_), .B2(new_n796_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n801_), .A2(new_n804_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n802_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n801_), .A2(new_n802_), .A3(new_n804_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n871_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(KEYINPUT121), .B1(new_n876_), .B2(new_n426_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n860_), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n807_), .A2(new_n880_), .A3(new_n427_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n592_), .A2(new_n214_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n879_), .A2(new_n881_), .A3(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT122), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  NAND4_X1  g684(.A1(new_n879_), .A2(KEYINPUT122), .A3(new_n881_), .A4(new_n882_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n214_), .B1(new_n867_), .B2(new_n592_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(KEYINPUT120), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT120), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n889_), .B(new_n214_), .C1(new_n867_), .C2(new_n592_), .ZN(new_n890_));
  AOI22_X1  g689(.A1(new_n885_), .A2(new_n886_), .B1(new_n888_), .B2(new_n890_), .ZN(G1349gat));
  NAND4_X1  g690(.A1(new_n877_), .A2(new_n881_), .A3(new_n609_), .A4(new_n878_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n203_), .ZN(new_n893_));
  AND2_X1   g692(.A1(new_n204_), .A2(new_n206_), .ZN(new_n894_));
  OR3_X1    g693(.A1(new_n867_), .A2(new_n894_), .A3(new_n608_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n893_), .A2(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT123), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n893_), .A2(new_n895_), .A3(KEYINPUT123), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(G1350gat));
  OAI21_X1  g699(.A(G190gat), .B1(new_n867_), .B2(new_n703_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n527_), .A2(new_n208_), .A3(new_n210_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n867_), .B2(new_n902_), .ZN(G1351gat));
  NAND4_X1  g702(.A1(new_n807_), .A2(new_n259_), .A3(new_n443_), .A4(new_n655_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT124), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n904_), .B(new_n905_), .ZN(new_n906_));
  NOR3_X1   g705(.A1(new_n906_), .A2(new_n323_), .A3(new_n669_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n904_), .B(KEYINPUT124), .ZN(new_n908_));
  AOI21_X1  g707(.A(G197gat), .B1(new_n908_), .B2(new_n556_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n907_), .A2(new_n909_), .ZN(G1352gat));
  AND2_X1   g709(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n911_));
  NOR2_X1   g710(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n912_));
  OAI211_X1 g711(.A(new_n908_), .B(new_n591_), .C1(new_n911_), .C2(new_n912_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n906_), .A2(new_n592_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n913_), .B1(new_n914_), .B2(new_n912_), .ZN(G1353gat));
  INV_X1    g714(.A(KEYINPUT126), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n916_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n917_));
  AOI211_X1 g716(.A(new_n917_), .B(new_n608_), .C1(KEYINPUT63), .C2(G211gat), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n908_), .A2(new_n918_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n916_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n920_));
  INV_X1    g719(.A(new_n920_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n919_), .A2(new_n921_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n908_), .A2(new_n920_), .A3(new_n918_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(G1354gat));
  NAND2_X1  g723(.A1(new_n908_), .A2(new_n527_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n653_), .A2(G218gat), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(KEYINPUT127), .ZN(new_n927_));
  AOI22_X1  g726(.A1(new_n925_), .A2(new_n318_), .B1(new_n908_), .B2(new_n927_), .ZN(G1355gat));
endmodule


