//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1 0 1 1 1 0 1 1 1 1 0 0 1 0 0 1 1 0 1 0 0 0 1 1 1 1 1 0 1 1 0 0 1 1 0 0 1 0 0 0 1 0 1 0 0 1 0 0 0 0 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n655_, new_n656_, new_n657_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n668_, new_n669_, new_n670_, new_n671_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n678_, new_n679_, new_n680_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n694_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n819_,
    new_n820_, new_n822_, new_n823_, new_n825_, new_n826_, new_n827_,
    new_n829_, new_n830_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n859_, new_n860_, new_n861_, new_n863_,
    new_n864_, new_n866_, new_n867_, new_n868_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G57gat), .B(G64gat), .ZN(new_n203_));
  OR2_X1    g002(.A1(new_n203_), .A2(KEYINPUT11), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(KEYINPUT11), .ZN(new_n205_));
  XOR2_X1   g004(.A(G71gat), .B(G78gat), .Z(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  OR2_X1    g006(.A1(new_n205_), .A2(new_n206_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G99gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT10), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT10), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(G99gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT64), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT64), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n212_), .A2(new_n214_), .A3(new_n217_), .ZN(new_n218_));
  AOI21_X1  g017(.A(G106gat), .B1(new_n216_), .B2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G99gat), .A2(G106gat), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT65), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n222_), .A2(KEYINPUT6), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT6), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n224_), .A2(KEYINPUT65), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n221_), .B1(new_n223_), .B2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(KEYINPUT65), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n222_), .A2(KEYINPUT6), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(new_n228_), .A3(new_n220_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G85gat), .A2(G92gat), .ZN(new_n230_));
  OR2_X1    g029(.A1(new_n230_), .A2(KEYINPUT9), .ZN(new_n231_));
  INV_X1    g030(.A(G85gat), .ZN(new_n232_));
  INV_X1    g031(.A(G92gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n234_), .A2(KEYINPUT9), .A3(new_n230_), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n226_), .A2(new_n229_), .A3(new_n231_), .A4(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT66), .B1(new_n219_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(G106gat), .ZN(new_n238_));
  AND3_X1   g037(.A1(new_n212_), .A2(new_n214_), .A3(new_n217_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n217_), .B1(new_n212_), .B2(new_n214_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n238_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n229_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n220_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n235_), .A2(new_n231_), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n241_), .A2(new_n244_), .A3(new_n245_), .A4(new_n246_), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n237_), .A2(new_n247_), .ZN(new_n248_));
  AND2_X1   g047(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n249_));
  NOR2_X1   g048(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n250_));
  OAI22_X1  g049(.A1(new_n249_), .A2(new_n250_), .B1(G99gat), .B2(G106gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n252_), .A2(new_n211_), .A3(new_n238_), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n226_), .A2(new_n229_), .A3(new_n251_), .A4(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT8), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n234_), .A2(new_n230_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n256_), .A2(KEYINPUT68), .ZN(new_n257_));
  AND3_X1   g056(.A1(new_n254_), .A2(new_n255_), .A3(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n255_), .B1(new_n254_), .B2(new_n257_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n210_), .B1(new_n248_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT69), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n254_), .A2(new_n257_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT8), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n254_), .A2(new_n257_), .A3(new_n255_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n237_), .A2(new_n247_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n266_), .A2(new_n267_), .A3(new_n209_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n261_), .A2(new_n262_), .A3(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G230gat), .A2(G233gat), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n248_), .A2(new_n260_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n272_), .A2(KEYINPUT69), .A3(new_n209_), .ZN(new_n273_));
  AND3_X1   g072(.A1(new_n269_), .A2(new_n271_), .A3(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n261_), .A2(KEYINPUT12), .A3(new_n268_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n266_), .A2(new_n267_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT12), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n276_), .A2(new_n277_), .A3(new_n210_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n271_), .B1(new_n275_), .B2(new_n278_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n274_), .A2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G120gat), .B(G148gat), .ZN(new_n281_));
  INV_X1    g080(.A(G204gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT5), .B(G176gat), .ZN(new_n284_));
  XOR2_X1   g083(.A(new_n283_), .B(new_n284_), .Z(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT70), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n280_), .B(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT71), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n288_), .B1(new_n289_), .B2(KEYINPUT13), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n289_), .A2(KEYINPUT13), .ZN(new_n291_));
  OR2_X1    g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n291_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G229gat), .A2(G233gat), .ZN(new_n295_));
  OR2_X1    g094(.A1(KEYINPUT75), .A2(G15gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(KEYINPUT75), .A2(G15gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(G22gat), .ZN(new_n299_));
  INV_X1    g098(.A(G22gat), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n296_), .A2(new_n300_), .A3(new_n297_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT76), .B(G8gat), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT14), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  OAI21_X1  g104(.A(G1gat), .B1(new_n302_), .B2(new_n305_), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n299_), .A2(new_n304_), .A3(new_n202_), .A4(new_n301_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(G8gat), .ZN(new_n309_));
  INV_X1    g108(.A(G8gat), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n306_), .A2(new_n310_), .A3(new_n307_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G29gat), .B(G36gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G43gat), .B(G50gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT15), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n312_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT78), .ZN(new_n318_));
  AND3_X1   g117(.A1(new_n306_), .A2(new_n310_), .A3(new_n307_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n310_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n318_), .B1(new_n321_), .B2(new_n315_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n315_), .ZN(new_n323_));
  NOR4_X1   g122(.A1(new_n319_), .A2(new_n320_), .A3(KEYINPUT78), .A4(new_n323_), .ZN(new_n324_));
  OAI211_X1 g123(.A(new_n295_), .B(new_n317_), .C1(new_n322_), .C2(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n321_), .A2(new_n318_), .A3(new_n315_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n309_), .A2(new_n311_), .A3(new_n315_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT78), .ZN(new_n328_));
  AOI22_X1  g127(.A1(new_n326_), .A2(new_n328_), .B1(new_n312_), .B2(new_n323_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n325_), .B1(new_n329_), .B2(new_n295_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G113gat), .B(G141gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G169gat), .B(G197gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n330_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n333_), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n325_), .B(new_n335_), .C1(new_n329_), .C2(new_n295_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n294_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(G183gat), .ZN(new_n341_));
  OR3_X1    g140(.A1(new_n341_), .A2(KEYINPUT80), .A3(KEYINPUT25), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT26), .B(G190gat), .ZN(new_n343_));
  OAI21_X1  g142(.A(KEYINPUT80), .B1(new_n341_), .B2(KEYINPUT25), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n342_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT79), .B(G183gat), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n345_), .B1(KEYINPUT25), .B2(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(G169gat), .A2(G176gat), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  OR2_X1    g149(.A1(new_n350_), .A2(KEYINPUT24), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G183gat), .A2(G190gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT23), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G169gat), .A2(G176gat), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n350_), .A2(KEYINPUT24), .A3(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n351_), .A2(new_n353_), .A3(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n348_), .A2(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n353_), .B1(G190gat), .B2(new_n346_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT82), .ZN(new_n359_));
  INV_X1    g158(.A(G169gat), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT81), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT22), .ZN(new_n362_));
  INV_X1    g161(.A(G176gat), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n360_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n364_), .B1(new_n362_), .B2(new_n349_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n357_), .B1(new_n359_), .B2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G71gat), .B(G99gat), .ZN(new_n367_));
  INV_X1    g166(.A(G43gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n366_), .B(new_n369_), .ZN(new_n370_));
  XOR2_X1   g169(.A(G113gat), .B(G120gat), .Z(new_n371_));
  XNOR2_X1  g170(.A(G127gat), .B(G134gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n371_), .B(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G227gat), .A2(G233gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT30), .B(G15gat), .ZN(new_n376_));
  XOR2_X1   g175(.A(new_n376_), .B(KEYINPUT31), .Z(new_n377_));
  XNOR2_X1  g176(.A(new_n375_), .B(new_n377_), .ZN(new_n378_));
  OR2_X1    g177(.A1(new_n370_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n370_), .A2(new_n378_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(G78gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G228gat), .A2(G233gat), .ZN(new_n384_));
  INV_X1    g183(.A(G141gat), .ZN(new_n385_));
  INV_X1    g184(.A(G148gat), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n385_), .A2(new_n386_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n387_), .B1(KEYINPUT83), .B2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G155gat), .A2(G162gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(KEYINPUT1), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT1), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n392_), .A2(G155gat), .A3(G162gat), .ZN(new_n393_));
  OR2_X1    g192(.A1(G155gat), .A2(G162gat), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n391_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n389_), .B(new_n395_), .C1(KEYINPUT83), .C2(new_n388_), .ZN(new_n396_));
  OR3_X1    g195(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT2), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n398_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n399_));
  OAI21_X1  g198(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n400_));
  NAND3_X1  g199(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n397_), .A2(new_n399_), .A3(new_n400_), .A4(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n402_), .A2(new_n390_), .A3(new_n394_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n396_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(KEYINPUT29), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G197gat), .B(G204gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(KEYINPUT85), .ZN(new_n407_));
  INV_X1    g206(.A(G197gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(G204gat), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n407_), .B(KEYINPUT21), .C1(KEYINPUT85), .C2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT21), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n406_), .A2(KEYINPUT86), .A3(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G211gat), .B(G218gat), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT86), .ZN(new_n414_));
  INV_X1    g213(.A(new_n406_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n414_), .B1(new_n415_), .B2(KEYINPUT21), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n410_), .A2(new_n412_), .A3(new_n413_), .A4(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT88), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT87), .ZN(new_n419_));
  OR2_X1    g218(.A1(new_n413_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n413_), .A2(new_n419_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n420_), .A2(KEYINPUT21), .A3(new_n415_), .A4(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n417_), .A2(new_n418_), .A3(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n418_), .B1(new_n417_), .B2(new_n422_), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n384_), .B(new_n405_), .C1(new_n424_), .C2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n417_), .A2(new_n422_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n384_), .B1(new_n427_), .B2(new_n405_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n383_), .B1(new_n426_), .B2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n405_), .A2(new_n384_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n427_), .A2(KEYINPUT88), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n431_), .B1(new_n432_), .B2(new_n423_), .ZN(new_n433_));
  NOR3_X1   g232(.A1(new_n433_), .A2(G78gat), .A3(new_n428_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n238_), .B1(new_n430_), .B2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT84), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n426_), .A2(new_n383_), .A3(new_n429_), .ZN(new_n437_));
  OAI21_X1  g236(.A(G78gat), .B1(new_n433_), .B2(new_n428_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n437_), .A2(new_n438_), .A3(G106gat), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n435_), .A2(new_n436_), .A3(new_n439_), .ZN(new_n440_));
  OR2_X1    g239(.A1(new_n404_), .A2(KEYINPUT29), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(KEYINPUT28), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n440_), .A2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G22gat), .B(G50gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n445_), .B(KEYINPUT89), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n435_), .A2(new_n436_), .A3(new_n442_), .A4(new_n439_), .ZN(new_n447_));
  AND3_X1   g246(.A1(new_n444_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n446_), .B1(new_n444_), .B2(new_n447_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n382_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n444_), .A2(new_n447_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n446_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n444_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n453_), .A2(new_n454_), .A3(new_n381_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n450_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT95), .ZN(new_n457_));
  XNOR2_X1  g256(.A(KEYINPUT25), .B(G183gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(KEYINPUT92), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n356_), .B1(new_n459_), .B2(new_n343_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n353_), .B1(G183gat), .B2(G190gat), .ZN(new_n461_));
  INV_X1    g260(.A(new_n354_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(KEYINPUT22), .B(G169gat), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n462_), .B1(new_n463_), .B2(new_n363_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n460_), .B1(new_n461_), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n427_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n366_), .A2(new_n432_), .A3(new_n423_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(KEYINPUT20), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT91), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n467_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n468_), .A2(KEYINPUT91), .A3(KEYINPUT20), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G226gat), .A2(G233gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n457_), .B1(new_n473_), .B2(new_n477_), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n471_), .A2(KEYINPUT95), .A3(new_n476_), .A4(new_n472_), .ZN(new_n479_));
  AND2_X1   g278(.A1(new_n359_), .A2(new_n365_), .ZN(new_n480_));
  OAI22_X1  g279(.A1(new_n480_), .A2(new_n357_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT20), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n482_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n481_), .A2(new_n483_), .ZN(new_n484_));
  AND3_X1   g283(.A1(new_n484_), .A2(KEYINPUT94), .A3(new_n477_), .ZN(new_n485_));
  AOI21_X1  g284(.A(KEYINPUT94), .B1(new_n484_), .B2(new_n477_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n478_), .A2(new_n479_), .A3(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G8gat), .B(G36gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(new_n233_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(KEYINPUT18), .B(G64gat), .ZN(new_n491_));
  XOR2_X1   g290(.A(new_n490_), .B(new_n491_), .Z(new_n492_));
  NAND2_X1  g291(.A1(new_n488_), .A2(new_n492_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n484_), .A2(new_n477_), .ZN(new_n494_));
  AOI211_X1 g293(.A(new_n492_), .B(new_n494_), .C1(new_n473_), .C2(new_n477_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT27), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n493_), .A2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G1gat), .B(G29gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(new_n232_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(KEYINPUT0), .B(G57gat), .ZN(new_n501_));
  XOR2_X1   g300(.A(new_n500_), .B(new_n501_), .Z(new_n502_));
  NAND2_X1  g301(.A1(G225gat), .A2(G233gat), .ZN(new_n503_));
  XOR2_X1   g302(.A(new_n404_), .B(new_n373_), .Z(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT4), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT4), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n404_), .A2(new_n506_), .A3(new_n373_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n503_), .B1(new_n505_), .B2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n503_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n504_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n502_), .B1(new_n509_), .B2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n502_), .ZN(new_n514_));
  NOR3_X1   g313(.A1(new_n508_), .A2(new_n514_), .A3(new_n511_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n494_), .B1(new_n473_), .B2(new_n477_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n492_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n496_), .B1(new_n519_), .B2(new_n495_), .ZN(new_n520_));
  AND3_X1   g319(.A1(new_n498_), .A2(new_n516_), .A3(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n519_), .A2(new_n495_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT93), .ZN(new_n523_));
  NOR3_X1   g322(.A1(new_n513_), .A2(new_n523_), .A3(KEYINPUT33), .ZN(new_n524_));
  OAI221_X1 g323(.A(new_n514_), .B1(new_n523_), .B2(KEYINPUT33), .C1(new_n508_), .C2(new_n511_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n505_), .A2(new_n503_), .A3(new_n507_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n514_), .B1(new_n504_), .B2(new_n510_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n525_), .A2(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n524_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n522_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n518_), .A2(KEYINPUT32), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n488_), .A2(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n516_), .B1(new_n517_), .B2(new_n532_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n531_), .A2(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n382_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n538_));
  AOI22_X1  g337(.A1(new_n456_), .A2(new_n521_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n340_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n516_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G231gat), .A2(G233gat), .ZN(new_n542_));
  XOR2_X1   g341(.A(new_n209_), .B(new_n542_), .Z(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT77), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(new_n321_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G127gat), .B(G155gat), .ZN(new_n546_));
  INV_X1    g345(.A(G211gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(KEYINPUT16), .B(G183gat), .Z(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(KEYINPUT17), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n550_), .A2(KEYINPUT17), .ZN(new_n552_));
  AND3_X1   g351(.A1(new_n545_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n545_), .A2(new_n551_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  OR2_X1    g355(.A1(KEYINPUT74), .A2(KEYINPUT37), .ZN(new_n557_));
  NAND2_X1  g356(.A1(KEYINPUT74), .A2(KEYINPUT37), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n276_), .A2(new_n316_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G232gat), .A2(G233gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT73), .ZN(new_n561_));
  XNOR2_X1  g360(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n563_), .A2(KEYINPUT35), .ZN(new_n564_));
  OAI211_X1 g363(.A(new_n559_), .B(new_n564_), .C1(new_n323_), .C2(new_n276_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(KEYINPUT35), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  OR2_X1    g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G190gat), .B(G218gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G134gat), .B(G162gat), .ZN(new_n570_));
  XOR2_X1   g369(.A(new_n569_), .B(new_n570_), .Z(new_n571_));
  INV_X1    g370(.A(KEYINPUT36), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n565_), .A2(new_n567_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n568_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n571_), .B(KEYINPUT36), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n579_), .B1(new_n568_), .B2(new_n575_), .ZN(new_n580_));
  OAI211_X1 g379(.A(new_n557_), .B(new_n558_), .C1(new_n577_), .C2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n580_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n582_), .A2(KEYINPUT74), .A3(KEYINPUT37), .A4(new_n576_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n556_), .A2(new_n584_), .ZN(new_n585_));
  AND4_X1   g384(.A1(new_n202_), .A2(new_n540_), .A3(new_n541_), .A4(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  XOR2_X1   g387(.A(new_n588_), .B(KEYINPUT98), .Z(new_n589_));
  NAND2_X1  g388(.A1(new_n582_), .A2(new_n576_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n556_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n540_), .A2(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(G1gat), .B1(new_n593_), .B2(new_n516_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n586_), .A2(new_n587_), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n595_), .B(KEYINPUT97), .Z(new_n596_));
  NAND3_X1  g395(.A1(new_n589_), .A2(new_n594_), .A3(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(KEYINPUT99), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT99), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n589_), .A2(new_n596_), .A3(new_n599_), .A4(new_n594_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(G1324gat));
  AND2_X1   g400(.A1(new_n498_), .A2(new_n520_), .ZN(new_n602_));
  OAI21_X1  g401(.A(G8gat), .B1(new_n593_), .B2(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT39), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n540_), .A2(new_n585_), .ZN(new_n605_));
  OR2_X1    g404(.A1(new_n602_), .A2(new_n303_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n604_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n607_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g407(.A(G15gat), .B1(new_n593_), .B2(new_n381_), .ZN(new_n609_));
  XOR2_X1   g408(.A(KEYINPUT100), .B(KEYINPUT41), .Z(new_n610_));
  OR2_X1    g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(new_n610_), .ZN(new_n612_));
  OR3_X1    g411(.A1(new_n605_), .A2(G15gat), .A3(new_n381_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n611_), .A2(new_n612_), .A3(new_n613_), .ZN(G1326gat));
  NAND2_X1  g413(.A1(new_n453_), .A2(new_n454_), .ZN(new_n615_));
  OAI21_X1  g414(.A(G22gat), .B1(new_n593_), .B2(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT42), .ZN(new_n617_));
  INV_X1    g416(.A(new_n615_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(new_n300_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n617_), .B1(new_n605_), .B2(new_n619_), .ZN(G1327gat));
  INV_X1    g419(.A(new_n584_), .ZN(new_n621_));
  OAI21_X1  g420(.A(KEYINPUT43), .B1(new_n539_), .B2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT43), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n498_), .A2(new_n516_), .A3(new_n520_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n624_), .B1(new_n455_), .B2(new_n450_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n537_), .A2(new_n538_), .ZN(new_n626_));
  OAI211_X1 g425(.A(new_n623_), .B(new_n584_), .C1(new_n625_), .C2(new_n626_), .ZN(new_n627_));
  AOI211_X1 g426(.A(new_n340_), .B(new_n555_), .C1(new_n622_), .C2(new_n627_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n628_), .A2(KEYINPUT44), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n628_), .A2(KEYINPUT44), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(G29gat), .B1(new_n632_), .B2(new_n516_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n555_), .A2(new_n590_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n540_), .A2(new_n634_), .ZN(new_n635_));
  OR3_X1    g434(.A1(new_n635_), .A2(G29gat), .A3(new_n516_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n633_), .A2(new_n636_), .ZN(G1328gat));
  INV_X1    g436(.A(G36gat), .ZN(new_n638_));
  INV_X1    g437(.A(new_n602_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n638_), .B1(new_n631_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT46), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n635_), .A2(G36gat), .A3(new_n602_), .ZN(new_n642_));
  XOR2_X1   g441(.A(KEYINPUT101), .B(KEYINPUT45), .Z(new_n643_));
  XNOR2_X1  g442(.A(new_n642_), .B(new_n643_), .ZN(new_n644_));
  OR3_X1    g443(.A1(new_n640_), .A2(new_n641_), .A3(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n641_), .B1(new_n640_), .B2(new_n644_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(G1329gat));
  AOI21_X1  g446(.A(new_n368_), .B1(new_n631_), .B2(new_n382_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n635_), .A2(G43gat), .A3(new_n381_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(KEYINPUT102), .B(KEYINPUT47), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  OR3_X1    g450(.A1(new_n648_), .A2(new_n649_), .A3(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n651_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1330gat));
  OAI21_X1  g453(.A(G50gat), .B1(new_n632_), .B2(new_n615_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n615_), .A2(G50gat), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n656_), .B(KEYINPUT103), .Z(new_n657_));
  OAI21_X1  g456(.A(new_n655_), .B1(new_n635_), .B2(new_n657_), .ZN(G1331gat));
  NAND2_X1  g457(.A1(new_n294_), .A2(new_n338_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n539_), .A2(new_n659_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n660_), .A2(new_n585_), .ZN(new_n661_));
  AOI21_X1  g460(.A(G57gat), .B1(new_n661_), .B2(new_n541_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n592_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n516_), .A2(KEYINPUT104), .ZN(new_n665_));
  MUX2_X1   g464(.A(KEYINPUT104), .B(new_n665_), .S(G57gat), .Z(new_n666_));
  AOI21_X1  g465(.A(new_n662_), .B1(new_n664_), .B2(new_n666_), .ZN(G1332gat));
  OAI21_X1  g466(.A(G64gat), .B1(new_n663_), .B2(new_n602_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT48), .ZN(new_n669_));
  INV_X1    g468(.A(G64gat), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n661_), .A2(new_n670_), .A3(new_n639_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(G1333gat));
  OAI21_X1  g471(.A(G71gat), .B1(new_n663_), .B2(new_n381_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT49), .ZN(new_n674_));
  INV_X1    g473(.A(G71gat), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n661_), .A2(new_n675_), .A3(new_n382_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n676_), .ZN(G1334gat));
  OAI21_X1  g476(.A(G78gat), .B1(new_n663_), .B2(new_n615_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT50), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n661_), .A2(new_n383_), .A3(new_n618_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(G1335gat));
  NAND2_X1  g480(.A1(new_n660_), .A2(new_n634_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(G85gat), .B1(new_n683_), .B2(new_n541_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n622_), .A2(new_n627_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n294_), .A2(new_n338_), .A3(new_n556_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(KEYINPUT105), .B1(new_n685_), .B2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT105), .ZN(new_n689_));
  AOI211_X1 g488(.A(new_n689_), .B(new_n686_), .C1(new_n622_), .C2(new_n627_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n688_), .A2(new_n690_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n516_), .A2(new_n232_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n684_), .B1(new_n691_), .B2(new_n692_), .ZN(G1336gat));
  AOI21_X1  g492(.A(G92gat), .B1(new_n683_), .B2(new_n639_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n602_), .A2(new_n233_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n691_), .B2(new_n695_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT106), .ZN(G1337gat));
  INV_X1    g496(.A(KEYINPUT107), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n382_), .B1(new_n240_), .B2(new_n239_), .ZN(new_n699_));
  OR3_X1    g498(.A1(new_n682_), .A2(new_n698_), .A3(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n698_), .B1(new_n682_), .B2(new_n699_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(KEYINPUT108), .B(KEYINPUT51), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n688_), .A2(new_n690_), .A3(new_n381_), .ZN(new_n704_));
  OAI211_X1 g503(.A(new_n702_), .B(new_n703_), .C1(new_n704_), .C2(new_n211_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(KEYINPUT109), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n622_), .A2(new_n627_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n689_), .B1(new_n707_), .B2(new_n686_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n685_), .A2(KEYINPUT105), .A3(new_n687_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n708_), .A2(new_n382_), .A3(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(G99gat), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n712_));
  NAND4_X1  g511(.A1(new_n711_), .A2(new_n712_), .A3(new_n702_), .A4(new_n703_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n211_), .B1(new_n691_), .B2(new_n382_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n702_), .ZN(new_n715_));
  OAI21_X1  g514(.A(KEYINPUT51), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n706_), .A2(new_n713_), .A3(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(KEYINPUT110), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT110), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n706_), .A2(new_n713_), .A3(new_n716_), .A4(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(G1338gat));
  NAND3_X1  g520(.A1(new_n683_), .A2(new_n238_), .A3(new_n618_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT52), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n707_), .A2(new_n686_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(new_n618_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n723_), .B1(new_n725_), .B2(G106gat), .ZN(new_n726_));
  AOI211_X1 g525(.A(KEYINPUT52), .B(new_n238_), .C1(new_n724_), .C2(new_n618_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n722_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n728_), .B(new_n729_), .Z(G1339gat));
  INV_X1    g529(.A(KEYINPUT113), .ZN(new_n731_));
  NOR3_X1   g530(.A1(new_n274_), .A2(new_n279_), .A3(new_n286_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n732_), .B1(new_n334_), .B2(new_n336_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n275_), .A2(new_n271_), .A3(new_n278_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT55), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n275_), .A2(new_n278_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n736_), .B2(new_n270_), .ZN(new_n737_));
  AOI211_X1 g536(.A(KEYINPUT55), .B(new_n271_), .C1(new_n275_), .C2(new_n278_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n734_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n739_), .A2(KEYINPUT56), .A3(new_n286_), .ZN(new_n740_));
  AOI21_X1  g539(.A(KEYINPUT56), .B1(new_n739_), .B2(new_n286_), .ZN(new_n741_));
  OAI211_X1 g540(.A(new_n731_), .B(new_n733_), .C1(new_n740_), .C2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n295_), .ZN(new_n743_));
  OAI211_X1 g542(.A(new_n743_), .B(new_n317_), .C1(new_n322_), .C2(new_n324_), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n744_), .B(new_n333_), .C1(new_n329_), .C2(new_n743_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n288_), .A2(new_n336_), .A3(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n742_), .A2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT56), .ZN(new_n748_));
  INV_X1    g547(.A(new_n734_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n268_), .A2(KEYINPUT12), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n209_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n278_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n270_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(KEYINPUT55), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n279_), .A2(new_n735_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n749_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n748_), .B1(new_n757_), .B2(new_n285_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n739_), .A2(KEYINPUT56), .A3(new_n286_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n731_), .B1(new_n760_), .B2(new_n733_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n590_), .B1(new_n747_), .B2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT57), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT114), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n758_), .A2(new_n765_), .A3(new_n759_), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n739_), .A2(KEYINPUT114), .A3(KEYINPUT56), .A4(new_n286_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n336_), .A2(new_n745_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n768_), .A2(new_n732_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n767_), .A2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n766_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT58), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n621_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n766_), .A2(new_n770_), .A3(KEYINPUT58), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT115), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n766_), .A2(new_n770_), .A3(KEYINPUT115), .A4(KEYINPUT58), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n773_), .A2(new_n776_), .A3(new_n777_), .ZN(new_n778_));
  OAI211_X1 g577(.A(KEYINPUT57), .B(new_n590_), .C1(new_n747_), .C2(new_n761_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n764_), .A2(new_n778_), .A3(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT116), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT116), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n764_), .A2(new_n778_), .A3(new_n782_), .A4(new_n779_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n781_), .A2(new_n556_), .A3(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n294_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n785_), .A2(new_n338_), .A3(new_n585_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n786_), .B(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n784_), .A2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT117), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT117), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n784_), .A2(new_n788_), .A3(new_n791_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n639_), .A2(new_n516_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n794_), .A2(new_n450_), .ZN(new_n795_));
  AND3_X1   g594(.A1(new_n790_), .A2(new_n792_), .A3(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(G113gat), .B1(new_n796_), .B2(new_n337_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT59), .ZN(new_n798_));
  AOI21_X1  g597(.A(KEYINPUT118), .B1(new_n764_), .B2(new_n778_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n779_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n764_), .A2(new_n778_), .A3(KEYINPUT118), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n555_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n788_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n795_), .A2(new_n798_), .ZN(new_n806_));
  OAI22_X1  g605(.A1(new_n796_), .A2(new_n798_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n337_), .A2(G113gat), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n797_), .B1(new_n808_), .B2(new_n809_), .ZN(G1340gat));
  XOR2_X1   g609(.A(KEYINPUT119), .B(G120gat), .Z(new_n811_));
  INV_X1    g610(.A(KEYINPUT60), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n812_), .B1(new_n785_), .B2(new_n811_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n790_), .A2(new_n792_), .A3(new_n795_), .A4(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n294_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n811_), .B1(new_n807_), .B2(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n796_), .A2(new_n812_), .A3(new_n813_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(G1341gat));
  AOI21_X1  g617(.A(G127gat), .B1(new_n796_), .B2(new_n555_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n555_), .A2(G127gat), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n819_), .B1(new_n808_), .B2(new_n820_), .ZN(G1342gat));
  AOI21_X1  g620(.A(G134gat), .B1(new_n796_), .B2(new_n591_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n584_), .A2(G134gat), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n822_), .B1(new_n808_), .B2(new_n823_), .ZN(G1343gat));
  INV_X1    g623(.A(new_n455_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n790_), .A2(new_n825_), .A3(new_n792_), .A4(new_n793_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n826_), .A2(new_n338_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(new_n385_), .ZN(G1344gat));
  NOR2_X1   g627(.A1(new_n826_), .A2(new_n785_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(KEYINPUT120), .B(G148gat), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n829_), .B(new_n830_), .ZN(G1345gat));
  AND3_X1   g630(.A1(new_n784_), .A2(new_n788_), .A3(new_n791_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n791_), .B1(new_n784_), .B2(new_n788_), .ZN(new_n833_));
  NOR3_X1   g632(.A1(new_n832_), .A2(new_n833_), .A3(new_n455_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT121), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n834_), .A2(new_n835_), .A3(new_n555_), .A4(new_n793_), .ZN(new_n836_));
  OAI21_X1  g635(.A(KEYINPUT121), .B1(new_n826_), .B2(new_n556_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(KEYINPUT61), .B(G155gat), .ZN(new_n838_));
  AND3_X1   g637(.A1(new_n836_), .A2(new_n837_), .A3(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n838_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n839_), .A2(new_n840_), .ZN(G1346gat));
  INV_X1    g640(.A(new_n826_), .ZN(new_n842_));
  AOI21_X1  g641(.A(G162gat), .B1(new_n842_), .B2(new_n591_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n584_), .A2(G162gat), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(KEYINPUT122), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n843_), .B1(new_n842_), .B2(new_n845_), .ZN(G1347gat));
  NOR2_X1   g645(.A1(new_n602_), .A2(new_n541_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n382_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n848_), .A2(new_n618_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n851_), .A2(new_n337_), .A3(new_n463_), .ZN(new_n852_));
  OAI21_X1  g651(.A(G169gat), .B1(new_n850_), .B2(new_n338_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT123), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(new_n854_), .A3(KEYINPUT62), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n855_), .B1(KEYINPUT62), .B2(new_n853_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n854_), .B1(new_n853_), .B2(KEYINPUT62), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n852_), .B1(new_n856_), .B2(new_n857_), .ZN(G1348gat));
  AOI21_X1  g657(.A(G176gat), .B1(new_n851_), .B2(new_n294_), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n832_), .A2(new_n833_), .A3(new_n618_), .ZN(new_n860_));
  NOR3_X1   g659(.A1(new_n848_), .A2(new_n785_), .A3(new_n363_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n859_), .B1(new_n860_), .B2(new_n861_), .ZN(G1349gat));
  NOR3_X1   g661(.A1(new_n850_), .A2(new_n459_), .A3(new_n556_), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n860_), .A2(new_n382_), .A3(new_n555_), .A4(new_n847_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n863_), .B1(new_n864_), .B2(new_n347_), .ZN(G1350gat));
  NAND3_X1  g664(.A1(new_n851_), .A2(new_n343_), .A3(new_n591_), .ZN(new_n866_));
  OAI21_X1  g665(.A(G190gat), .B1(new_n850_), .B2(new_n621_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(KEYINPUT124), .ZN(G1351gat));
  NAND4_X1  g668(.A1(new_n790_), .A2(new_n825_), .A3(new_n792_), .A4(new_n847_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n870_), .A2(new_n338_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(new_n408_), .ZN(G1352gat));
  NOR2_X1   g671(.A1(new_n870_), .A2(new_n785_), .ZN(new_n873_));
  OR2_X1    g672(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  XOR2_X1   g674(.A(KEYINPUT125), .B(G204gat), .Z(new_n876_));
  AOI21_X1  g675(.A(new_n875_), .B1(new_n873_), .B2(new_n876_), .ZN(G1353gat));
  INV_X1    g676(.A(KEYINPUT63), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n878_), .A2(new_n547_), .A3(KEYINPUT126), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n555_), .B(new_n879_), .C1(new_n878_), .C2(new_n547_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n870_), .A2(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(KEYINPUT126), .B1(new_n878_), .B2(new_n547_), .ZN(new_n882_));
  XOR2_X1   g681(.A(new_n881_), .B(new_n882_), .Z(G1354gat));
  NAND4_X1  g682(.A1(new_n834_), .A2(G218gat), .A3(new_n584_), .A4(new_n847_), .ZN(new_n884_));
  INV_X1    g683(.A(G218gat), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n885_), .B1(new_n870_), .B2(new_n590_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n884_), .A2(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT127), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n884_), .A2(new_n886_), .A3(KEYINPUT127), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(G1355gat));
endmodule


