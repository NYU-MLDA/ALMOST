//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 1 0 1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 1 1 0 1 1 1 0 1 0 0 0 1 0 1 0 0 0 0 0 0 0 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n681_, new_n682_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n830_, new_n831_,
    new_n832_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n841_, new_n842_, new_n843_, new_n845_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n869_,
    new_n870_, new_n871_, new_n873_, new_n874_, new_n875_, new_n876_,
    new_n877_, new_n878_, new_n879_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT65), .ZN(new_n204_));
  XOR2_X1   g003(.A(G71gat), .B(G78gat), .Z(new_n205_));
  OAI21_X1  g004(.A(new_n205_), .B1(KEYINPUT11), .B2(new_n202_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n204_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  XOR2_X1   g007(.A(G85gat), .B(G92gat), .Z(new_n209_));
  NAND2_X1  g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  XOR2_X1   g009(.A(new_n210_), .B(KEYINPUT6), .Z(new_n211_));
  OR3_X1    g010(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n209_), .B1(new_n211_), .B2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n215_), .B(KEYINPUT8), .ZN(new_n216_));
  INV_X1    g015(.A(G106gat), .ZN(new_n217_));
  XOR2_X1   g016(.A(KEYINPUT10), .B(G99gat), .Z(new_n218_));
  AOI21_X1  g017(.A(new_n211_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n220_));
  XOR2_X1   g019(.A(KEYINPUT64), .B(G85gat), .Z(new_n221_));
  INV_X1    g020(.A(G92gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n220_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n219_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n216_), .A2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n208_), .B(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT12), .ZN(new_n229_));
  AND2_X1   g028(.A1(new_n216_), .A2(new_n226_), .ZN(new_n230_));
  OR3_X1    g029(.A1(new_n230_), .A2(new_n208_), .A3(KEYINPUT12), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G230gat), .A2(G233gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n234_), .B1(new_n233_), .B2(new_n228_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G120gat), .B(G148gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(G204gat), .ZN(new_n237_));
  XOR2_X1   g036(.A(KEYINPUT5), .B(G176gat), .Z(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  XOR2_X1   g038(.A(new_n235_), .B(new_n239_), .Z(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(KEYINPUT13), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT72), .B(G22gat), .ZN(new_n242_));
  INV_X1    g041(.A(G15gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT14), .ZN(new_n245_));
  XOR2_X1   g044(.A(KEYINPUT73), .B(G1gat), .Z(new_n246_));
  AOI21_X1  g045(.A(new_n245_), .B1(new_n246_), .B2(G8gat), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n244_), .A2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT74), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(G1gat), .ZN(new_n250_));
  INV_X1    g049(.A(G8gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  OR2_X1    g051(.A1(new_n249_), .A2(G1gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n249_), .A2(G1gat), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n253_), .A2(G8gat), .A3(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n252_), .A2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G29gat), .B(G36gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G43gat), .B(G50gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n256_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT77), .ZN(new_n261_));
  INV_X1    g060(.A(new_n259_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n252_), .A2(new_n255_), .A3(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n260_), .A2(new_n261_), .A3(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G229gat), .A2(G233gat), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n256_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n267_), .A2(KEYINPUT77), .A3(new_n262_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n264_), .A2(new_n266_), .A3(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n259_), .B(KEYINPUT15), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n267_), .A2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n271_), .A2(new_n265_), .A3(new_n260_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n269_), .A2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G113gat), .B(G141gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(G169gat), .ZN(new_n275_));
  INV_X1    g074(.A(G197gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n273_), .A2(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n269_), .A2(new_n272_), .A3(new_n277_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n241_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n230_), .A2(new_n259_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n227_), .A2(new_n270_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G232gat), .A2(G233gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT34), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT66), .B(KEYINPUT35), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n284_), .A2(new_n285_), .A3(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n288_), .A2(new_n289_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n292_), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n284_), .A2(new_n294_), .A3(new_n285_), .A4(new_n290_), .ZN(new_n295_));
  AND2_X1   g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G190gat), .B(G218gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT67), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(G134gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(G162gat), .ZN(new_n300_));
  INV_X1    g099(.A(G134gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n298_), .B(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(G162gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n300_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(KEYINPUT36), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n296_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT36), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n300_), .A2(new_n304_), .A3(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT68), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n293_), .A2(new_n312_), .A3(new_n295_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT69), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT69), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n293_), .A2(new_n312_), .A3(new_n315_), .A4(new_n295_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n308_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT37), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT70), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n307_), .B1(new_n317_), .B2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n314_), .A2(KEYINPUT70), .A3(new_n316_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n320_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT71), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n321_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n327_), .B1(new_n326_), .B2(new_n325_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G231gat), .A2(G233gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n256_), .B(new_n329_), .ZN(new_n330_));
  OR2_X1    g129(.A1(new_n330_), .A2(new_n207_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n207_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT17), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G183gat), .B(G211gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G127gat), .B(G155gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  NOR3_X1   g138(.A1(new_n333_), .A2(new_n334_), .A3(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(KEYINPUT17), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n342_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n343_));
  OR2_X1    g142(.A1(new_n340_), .A2(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(KEYINPUT76), .B1(new_n328_), .B2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT27), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT89), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G197gat), .B(G204gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(KEYINPUT85), .ZN(new_n349_));
  INV_X1    g148(.A(G218gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(G211gat), .ZN(new_n351_));
  INV_X1    g150(.A(G211gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(G218gat), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT86), .ZN(new_n354_));
  AND3_X1   g153(.A1(new_n351_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n354_), .B1(new_n351_), .B2(new_n353_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n349_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n352_), .A2(G218gat), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n350_), .A2(G211gat), .ZN(new_n359_));
  OAI21_X1  g158(.A(KEYINPUT86), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n351_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n360_), .A2(new_n361_), .A3(new_n348_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n357_), .A2(new_n362_), .A3(KEYINPUT21), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT21), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n349_), .B(new_n364_), .C1(new_n355_), .C2(new_n356_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  NOR3_X1   g165(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT24), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n368_), .B1(G169gat), .B2(G176gat), .ZN(new_n369_));
  OR2_X1    g168(.A1(G169gat), .A2(G176gat), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n367_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(G183gat), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT25), .B1(new_n372_), .B2(KEYINPUT78), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT78), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT25), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n374_), .A2(new_n375_), .A3(G183gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(KEYINPUT79), .A2(G190gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(KEYINPUT26), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT26), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n379_), .A2(KEYINPUT79), .A3(G190gat), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n373_), .A2(new_n376_), .A3(new_n378_), .A4(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G183gat), .A2(G190gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(KEYINPUT80), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT80), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n384_), .A2(G183gat), .A3(G190gat), .ZN(new_n385_));
  AOI21_X1  g184(.A(KEYINPUT23), .B1(new_n383_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT23), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n387_), .B1(G183gat), .B2(G190gat), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n371_), .B(new_n381_), .C1(new_n386_), .C2(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(G183gat), .A2(G190gat), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT81), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n391_), .B1(new_n382_), .B2(KEYINPUT23), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n387_), .A2(KEYINPUT81), .A3(G183gat), .A4(G190gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n383_), .A2(new_n385_), .A3(KEYINPUT23), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n390_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G169gat), .A2(G176gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT22), .B(G169gat), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n397_), .B1(new_n399_), .B2(G176gat), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n389_), .B1(new_n396_), .B2(new_n400_), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n347_), .B(KEYINPUT20), .C1(new_n366_), .C2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n397_), .B(KEYINPUT91), .ZN(new_n403_));
  INV_X1    g202(.A(G176gat), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n403_), .B1(new_n404_), .B2(new_n398_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n386_), .A2(new_n388_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n405_), .B1(new_n390_), .B2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(KEYINPUT25), .B(G183gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n379_), .A2(G190gat), .ZN(new_n409_));
  INV_X1    g208(.A(G190gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT26), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT90), .ZN(new_n412_));
  AND3_X1   g211(.A1(new_n409_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n412_), .B1(new_n409_), .B2(new_n411_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n408_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n394_), .A2(new_n395_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n415_), .A2(new_n416_), .A3(new_n371_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n407_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(new_n366_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n402_), .A2(new_n419_), .ZN(new_n420_));
  OR2_X1    g219(.A1(new_n396_), .A2(new_n400_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n421_), .A2(new_n363_), .A3(new_n365_), .A4(new_n389_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n347_), .B1(new_n422_), .B2(KEYINPUT20), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n420_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n366_), .A2(new_n401_), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n425_), .B(KEYINPUT20), .C1(new_n366_), .C2(new_n418_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G226gat), .A2(G233gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(KEYINPUT19), .ZN(new_n428_));
  MUX2_X1   g227(.A(new_n424_), .B(new_n426_), .S(new_n428_), .Z(new_n429_));
  XNOR2_X1  g228(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G8gat), .B(G36gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n430_), .B(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G64gat), .B(G92gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n432_), .B(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n346_), .B1(new_n429_), .B2(new_n434_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n426_), .A2(new_n428_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n428_), .B1(new_n420_), .B2(new_n423_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT92), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n436_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n434_), .ZN(new_n440_));
  OAI211_X1 g239(.A(KEYINPUT92), .B(new_n428_), .C1(new_n420_), .C2(new_n423_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n439_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n435_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT100), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n439_), .A2(new_n441_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(new_n434_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(KEYINPUT94), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n440_), .B1(new_n439_), .B2(new_n441_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT94), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n447_), .A2(new_n450_), .A3(new_n442_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n444_), .B1(new_n451_), .B2(new_n346_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n442_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n453_));
  AOI211_X1 g252(.A(KEYINPUT94), .B(new_n440_), .C1(new_n439_), .C2(new_n441_), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n444_), .B(new_n346_), .C1(new_n453_), .C2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n443_), .B1(new_n452_), .B2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT101), .ZN(new_n458_));
  INV_X1    g257(.A(new_n443_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n346_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT100), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n459_), .B1(new_n461_), .B2(new_n455_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT101), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT88), .ZN(new_n465_));
  AND2_X1   g264(.A1(G228gat), .A2(G233gat), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT84), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n466_), .B1(new_n366_), .B2(new_n467_), .ZN(new_n468_));
  NOR3_X1   g267(.A1(KEYINPUT83), .A2(G155gat), .A3(G162gat), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(KEYINPUT83), .B1(G155gat), .B2(G162gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G155gat), .A2(G162gat), .ZN(new_n473_));
  NOR2_X1   g272(.A1(G141gat), .A2(G148gat), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT3), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G141gat), .A2(G148gat), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT2), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n472_), .B(new_n473_), .C1(new_n476_), .C2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n474_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n471_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n482_), .A2(new_n469_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n473_), .B(KEYINPUT1), .ZN(new_n484_));
  OAI211_X1 g283(.A(new_n477_), .B(new_n481_), .C1(new_n483_), .C2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n480_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT29), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(new_n366_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n468_), .A2(new_n488_), .ZN(new_n489_));
  OAI211_X1 g288(.A(new_n487_), .B(new_n366_), .C1(new_n467_), .C2(new_n466_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G78gat), .B(G106gat), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n491_), .A2(KEYINPUT87), .A3(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n489_), .A2(new_n492_), .A3(new_n490_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n486_), .A2(KEYINPUT29), .ZN(new_n496_));
  XOR2_X1   g295(.A(G22gat), .B(G50gat), .Z(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT28), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n496_), .B(new_n498_), .ZN(new_n499_));
  AND3_X1   g298(.A1(new_n494_), .A2(new_n495_), .A3(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(KEYINPUT87), .B1(new_n491_), .B2(new_n493_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n465_), .B1(new_n500_), .B2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n494_), .A2(new_n495_), .A3(new_n499_), .ZN(new_n504_));
  NOR3_X1   g303(.A1(new_n504_), .A2(KEYINPUT88), .A3(new_n501_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n491_), .A2(new_n493_), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n506_), .A2(new_n495_), .ZN(new_n507_));
  OAI22_X1  g306(.A1(new_n503_), .A2(new_n505_), .B1(new_n507_), .B2(new_n499_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  XOR2_X1   g308(.A(new_n401_), .B(KEYINPUT30), .Z(new_n510_));
  XOR2_X1   g309(.A(G71gat), .B(G99gat), .Z(new_n511_));
  NAND2_X1  g310(.A1(G227gat), .A2(G233gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n510_), .B(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G127gat), .B(G134gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G113gat), .B(G120gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n514_), .B(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G15gat), .B(G43gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT31), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n518_), .B(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G225gat), .A2(G233gat), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n517_), .B1(new_n480_), .B2(new_n485_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n480_), .A2(new_n485_), .A3(new_n517_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n523_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n525_), .A2(KEYINPUT4), .A3(new_n526_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT4), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n524_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n527_), .B1(new_n531_), .B2(new_n523_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G1gat), .B(G29gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT0), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(G57gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(G85gat), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n532_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT98), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT98), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n532_), .A2(new_n539_), .A3(new_n536_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n531_), .A2(new_n523_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n527_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n536_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n538_), .A2(new_n540_), .A3(new_n544_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n521_), .A2(new_n545_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n458_), .A2(new_n464_), .A3(new_n509_), .A4(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n521_), .B(KEYINPUT82), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT95), .ZN(new_n549_));
  OAI21_X1  g348(.A(KEYINPUT33), .B1(new_n543_), .B2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n525_), .A2(new_n526_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n536_), .B1(new_n522_), .B2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT96), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT96), .ZN(new_n554_));
  OAI211_X1 g353(.A(new_n536_), .B(new_n554_), .C1(new_n522_), .C2(new_n551_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n528_), .A2(new_n522_), .A3(new_n530_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n553_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT33), .ZN(new_n558_));
  OAI211_X1 g357(.A(KEYINPUT95), .B(new_n558_), .C1(new_n532_), .C2(new_n536_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n550_), .A2(new_n557_), .A3(new_n559_), .ZN(new_n560_));
  NOR3_X1   g359(.A1(new_n453_), .A2(new_n454_), .A3(new_n560_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n440_), .A2(KEYINPUT32), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n562_), .B(KEYINPUT97), .Z(new_n563_));
  NAND3_X1  g362(.A1(new_n563_), .A2(new_n441_), .A3(new_n439_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n429_), .A2(new_n562_), .ZN(new_n565_));
  AND3_X1   g364(.A1(new_n545_), .A2(new_n564_), .A3(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n509_), .B1(new_n561_), .B2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(KEYINPUT99), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT99), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n509_), .B(new_n569_), .C1(new_n561_), .C2(new_n566_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n545_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n508_), .A2(new_n572_), .ZN(new_n573_));
  AOI211_X1 g372(.A(new_n459_), .B(new_n573_), .C1(new_n461_), .C2(new_n455_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n548_), .B1(new_n571_), .B2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n547_), .A2(new_n575_), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n325_), .A2(new_n326_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n325_), .A2(new_n326_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n577_), .A2(new_n578_), .A3(new_n321_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT76), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n340_), .A2(new_n343_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n579_), .A2(new_n580_), .A3(new_n581_), .ZN(new_n582_));
  AND4_X1   g381(.A1(new_n283_), .A2(new_n345_), .A3(new_n576_), .A4(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT102), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n585_), .A2(KEYINPUT38), .ZN(new_n586_));
  NOR4_X1   g385(.A1(new_n584_), .A2(new_n572_), .A3(new_n246_), .A4(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(KEYINPUT38), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n576_), .A2(new_n318_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n344_), .B1(new_n590_), .B2(KEYINPUT103), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT103), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n576_), .A2(new_n592_), .A3(new_n318_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n591_), .A2(new_n283_), .A3(new_n593_), .ZN(new_n594_));
  OAI21_X1  g393(.A(G1gat), .B1(new_n594_), .B2(new_n572_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n589_), .A2(new_n595_), .ZN(G1324gat));
  INV_X1    g395(.A(KEYINPUT40), .ZN(new_n597_));
  INV_X1    g396(.A(new_n464_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n462_), .A2(new_n463_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  OAI21_X1  g399(.A(G8gat), .B1(new_n594_), .B2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT39), .ZN(new_n602_));
  INV_X1    g401(.A(new_n600_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(new_n251_), .ZN(new_n604_));
  OAI21_X1  g403(.A(KEYINPUT104), .B1(new_n584_), .B2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT104), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n583_), .A2(new_n606_), .A3(new_n251_), .A4(new_n603_), .ZN(new_n607_));
  AOI22_X1  g406(.A1(new_n601_), .A2(new_n602_), .B1(new_n605_), .B2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT105), .ZN(new_n609_));
  OAI211_X1 g408(.A(KEYINPUT39), .B(G8gat), .C1(new_n594_), .C2(new_n600_), .ZN(new_n610_));
  AND3_X1   g409(.A1(new_n608_), .A2(new_n609_), .A3(new_n610_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n609_), .B1(new_n608_), .B2(new_n610_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n597_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n601_), .A2(new_n602_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n605_), .A2(new_n607_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n614_), .A2(new_n615_), .A3(new_n610_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(KEYINPUT105), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n608_), .A2(new_n609_), .A3(new_n610_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n617_), .A2(KEYINPUT40), .A3(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n613_), .A2(new_n619_), .ZN(G1325gat));
  OAI21_X1  g419(.A(G15gat), .B1(new_n594_), .B2(new_n548_), .ZN(new_n621_));
  XOR2_X1   g420(.A(new_n621_), .B(KEYINPUT41), .Z(new_n622_));
  INV_X1    g421(.A(new_n548_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n583_), .A2(new_n243_), .A3(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n622_), .A2(new_n624_), .ZN(G1326gat));
  OR3_X1    g424(.A1(new_n584_), .A2(G22gat), .A3(new_n509_), .ZN(new_n626_));
  OAI21_X1  g425(.A(G22gat), .B1(new_n594_), .B2(new_n509_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT106), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n629_), .A2(KEYINPUT42), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n629_), .A2(KEYINPUT42), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n626_), .B1(new_n630_), .B2(new_n631_), .ZN(G1327gat));
  NAND2_X1  g431(.A1(new_n283_), .A2(new_n344_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n318_), .B1(new_n547_), .B2(new_n575_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(G29gat), .B1(new_n637_), .B2(new_n545_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT43), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n639_), .B1(new_n576_), .B2(new_n328_), .ZN(new_n640_));
  AOI211_X1 g439(.A(KEYINPUT43), .B(new_n579_), .C1(new_n547_), .C2(new_n575_), .ZN(new_n641_));
  OAI211_X1 g440(.A(KEYINPUT44), .B(new_n634_), .C1(new_n640_), .C2(new_n641_), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n642_), .A2(G29gat), .A3(new_n545_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n634_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT44), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n638_), .B1(new_n643_), .B2(new_n646_), .ZN(G1328gat));
  INV_X1    g446(.A(KEYINPUT46), .ZN(new_n648_));
  XOR2_X1   g447(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n600_), .A2(KEYINPUT107), .ZN(new_n651_));
  INV_X1    g450(.A(G36gat), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT107), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n653_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n651_), .A2(new_n652_), .A3(new_n654_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n650_), .B1(new_n636_), .B2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n655_), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n657_), .A2(new_n634_), .A3(new_n635_), .A4(new_n649_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n646_), .A2(new_n603_), .A3(new_n642_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n659_), .B1(new_n660_), .B2(G36gat), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT109), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n648_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n642_), .A2(new_n603_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n652_), .B1(new_n664_), .B2(new_n646_), .ZN(new_n665_));
  NOR3_X1   g464(.A1(new_n665_), .A2(KEYINPUT109), .A3(new_n659_), .ZN(new_n666_));
  OAI21_X1  g465(.A(KEYINPUT110), .B1(new_n663_), .B2(new_n666_), .ZN(new_n667_));
  OAI21_X1  g466(.A(KEYINPUT109), .B1(new_n665_), .B2(new_n659_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n661_), .A2(new_n662_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT110), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n668_), .A2(new_n669_), .A3(new_n670_), .A4(new_n648_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n661_), .A2(KEYINPUT46), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n667_), .A2(new_n671_), .A3(new_n672_), .ZN(G1329gat));
  XOR2_X1   g472(.A(KEYINPUT111), .B(G43gat), .Z(new_n674_));
  OAI21_X1  g473(.A(new_n674_), .B1(new_n636_), .B2(new_n548_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n646_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n521_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n642_), .A2(G43gat), .A3(new_n677_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n675_), .B1(new_n676_), .B2(new_n678_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g479(.A(G50gat), .B1(new_n637_), .B2(new_n508_), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n642_), .A2(G50gat), .A3(new_n508_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n681_), .B1(new_n682_), .B2(new_n646_), .ZN(G1331gat));
  INV_X1    g482(.A(KEYINPUT13), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n240_), .B(new_n684_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n685_), .A2(new_n281_), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n591_), .A2(new_n593_), .A3(new_n686_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n545_), .A2(G57gat), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n687_), .B1(KEYINPUT112), .B2(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(G57gat), .B1(new_n689_), .B2(KEYINPUT112), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n345_), .A2(new_n582_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n691_), .A2(new_n576_), .A3(new_n686_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n689_), .A2(new_n545_), .A3(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n690_), .A2(new_n694_), .ZN(G1332gat));
  NAND2_X1  g494(.A1(new_n651_), .A2(new_n654_), .ZN(new_n696_));
  OR3_X1    g495(.A1(new_n692_), .A2(G64gat), .A3(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n696_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n687_), .A2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(G64gat), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n700_), .A2(KEYINPUT48), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n700_), .A2(KEYINPUT48), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n697_), .B1(new_n701_), .B2(new_n702_), .ZN(G1333gat));
  OR3_X1    g502(.A1(new_n692_), .A2(G71gat), .A3(new_n548_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n687_), .A2(new_n623_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(G71gat), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n706_), .A2(KEYINPUT49), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n706_), .A2(KEYINPUT49), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n704_), .B1(new_n707_), .B2(new_n708_), .ZN(G1334gat));
  OR3_X1    g508(.A1(new_n692_), .A2(G78gat), .A3(new_n509_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n687_), .A2(new_n508_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT50), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n711_), .A2(new_n712_), .A3(G78gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n711_), .B2(G78gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n710_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT113), .ZN(G1335gat));
  NOR3_X1   g515(.A1(new_n685_), .A2(new_n281_), .A3(new_n581_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n635_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(G85gat), .B1(new_n719_), .B2(new_n545_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n576_), .A2(new_n328_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(KEYINPUT43), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n576_), .A2(new_n639_), .A3(new_n328_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(new_n717_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT114), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n572_), .A2(new_n221_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n720_), .B1(new_n726_), .B2(new_n727_), .ZN(G1336gat));
  NAND3_X1  g527(.A1(new_n719_), .A2(new_n222_), .A3(new_n603_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n726_), .A2(new_n698_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n729_), .B1(new_n730_), .B2(new_n222_), .ZN(G1337gat));
  OAI21_X1  g530(.A(G99gat), .B1(new_n725_), .B2(new_n548_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n719_), .A2(new_n218_), .A3(new_n677_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g534(.A1(new_n719_), .A2(new_n217_), .A3(new_n508_), .ZN(new_n736_));
  OAI21_X1  g535(.A(G106gat), .B1(new_n725_), .B2(new_n509_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n737_), .A2(KEYINPUT52), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n737_), .A2(KEYINPUT52), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n736_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g540(.A(G113gat), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT57), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n264_), .A2(new_n265_), .A3(new_n268_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n271_), .A2(new_n266_), .A3(new_n260_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n744_), .A2(new_n278_), .A3(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n280_), .A2(new_n746_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n240_), .A2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n233_), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n229_), .A2(new_n749_), .A3(new_n231_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n229_), .B2(new_n231_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(KEYINPUT55), .B2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT55), .ZN(new_n753_));
  AOI21_X1  g552(.A(KEYINPUT115), .B1(new_n234_), .B2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT115), .ZN(new_n755_));
  NOR3_X1   g554(.A1(new_n751_), .A2(new_n755_), .A3(KEYINPUT55), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n752_), .B1(new_n754_), .B2(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(KEYINPUT56), .B1(new_n757_), .B2(new_n239_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n757_), .A2(KEYINPUT56), .A3(new_n239_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n235_), .A2(new_n239_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n762_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n748_), .B1(new_n761_), .B2(new_n763_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n743_), .B1(new_n764_), .B2(new_n319_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n760_), .B1(new_n758_), .B2(KEYINPUT117), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT117), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n757_), .A2(new_n767_), .A3(KEYINPUT56), .A4(new_n239_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n762_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n769_), .A2(new_n280_), .A3(new_n746_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT116), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT116), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n769_), .A2(new_n280_), .A3(new_n746_), .A4(new_n772_), .ZN(new_n773_));
  AOI22_X1  g572(.A1(new_n766_), .A2(new_n768_), .B1(new_n771_), .B2(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n328_), .B1(new_n774_), .B2(KEYINPUT58), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n766_), .A2(new_n768_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n771_), .A2(new_n773_), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n776_), .A2(KEYINPUT58), .A3(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n765_), .B1(new_n775_), .B2(new_n778_), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n764_), .A2(new_n743_), .A3(new_n319_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n344_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n579_), .A2(new_n685_), .A3(new_n282_), .A4(new_n581_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT54), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n782_), .B(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n781_), .A2(new_n785_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n603_), .A2(new_n508_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n521_), .A2(new_n572_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n786_), .A2(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n742_), .B1(new_n791_), .B2(new_n282_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT118), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT118), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n794_), .B(new_n742_), .C1(new_n791_), .C2(new_n282_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n793_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT59), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n790_), .A2(new_n797_), .ZN(new_n798_));
  OAI211_X1 g597(.A(new_n765_), .B(KEYINPUT119), .C1(new_n775_), .C2(new_n778_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n780_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n776_), .A2(new_n777_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT58), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n774_), .A2(KEYINPUT58), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n804_), .A2(new_n805_), .A3(new_n328_), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT119), .B1(new_n806_), .B2(new_n765_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n344_), .B1(new_n801_), .B2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n798_), .B1(new_n808_), .B2(new_n785_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n797_), .B1(new_n786_), .B2(new_n790_), .ZN(new_n810_));
  OAI21_X1  g609(.A(KEYINPUT120), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n806_), .A2(new_n800_), .A3(new_n765_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n784_), .B1(new_n812_), .B2(new_n344_), .ZN(new_n813_));
  OAI21_X1  g612(.A(KEYINPUT59), .B1(new_n813_), .B2(new_n789_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT120), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT119), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n779_), .A2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n817_), .A2(new_n800_), .A3(new_n799_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n784_), .B1(new_n818_), .B2(new_n344_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n814_), .B(new_n815_), .C1(new_n819_), .C2(new_n798_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n811_), .A2(new_n820_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n282_), .A2(new_n742_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n796_), .B1(new_n821_), .B2(new_n822_), .ZN(G1340gat));
  OAI21_X1  g622(.A(new_n814_), .B1(new_n819_), .B2(new_n798_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n685_), .A2(G120gat), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n786_), .B(new_n790_), .C1(KEYINPUT60), .C2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n241_), .ZN(new_n827_));
  OAI21_X1  g626(.A(G120gat), .B1(new_n824_), .B2(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n828_), .B1(KEYINPUT60), .B2(new_n826_), .ZN(G1341gat));
  AOI21_X1  g628(.A(new_n344_), .B1(new_n811_), .B2(new_n820_), .ZN(new_n830_));
  INV_X1    g629(.A(G127gat), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n581_), .A2(new_n831_), .ZN(new_n832_));
  OAI22_X1  g631(.A1(new_n830_), .A2(new_n831_), .B1(new_n791_), .B2(new_n832_), .ZN(G1342gat));
  OAI21_X1  g632(.A(new_n301_), .B1(new_n791_), .B2(new_n318_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(KEYINPUT121), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT121), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n836_), .B(new_n301_), .C1(new_n791_), .C2(new_n318_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n835_), .A2(new_n837_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n579_), .A2(new_n301_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n838_), .B1(new_n821_), .B2(new_n839_), .ZN(G1343gat));
  NOR2_X1   g639(.A1(new_n623_), .A2(new_n509_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n786_), .A2(new_n545_), .A3(new_n696_), .A4(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n842_), .A2(new_n282_), .ZN(new_n843_));
  XOR2_X1   g642(.A(new_n843_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g643(.A1(new_n842_), .A2(new_n685_), .ZN(new_n845_));
  XOR2_X1   g644(.A(new_n845_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g645(.A1(new_n842_), .A2(new_n344_), .ZN(new_n847_));
  XOR2_X1   g646(.A(KEYINPUT61), .B(G155gat), .Z(new_n848_));
  XNOR2_X1  g647(.A(new_n847_), .B(new_n848_), .ZN(G1346gat));
  OAI21_X1  g648(.A(G162gat), .B1(new_n842_), .B2(new_n579_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n319_), .A2(new_n303_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n850_), .B1(new_n842_), .B2(new_n851_), .ZN(G1347gat));
  NAND2_X1  g651(.A1(new_n808_), .A2(new_n785_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n696_), .A2(new_n545_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n855_), .A2(new_n548_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n853_), .A2(new_n281_), .A3(new_n509_), .A4(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(G169gat), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT62), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n857_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n860_), .B(new_n861_), .C1(new_n399_), .C2(new_n857_), .ZN(G1348gat));
  NOR2_X1   g661(.A1(new_n819_), .A2(new_n508_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n863_), .A2(new_n241_), .A3(new_n856_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n813_), .A2(new_n508_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n856_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n866_), .A2(new_n404_), .A3(new_n685_), .ZN(new_n867_));
  AOI22_X1  g666(.A1(new_n864_), .A2(new_n404_), .B1(new_n865_), .B2(new_n867_), .ZN(G1349gat));
  NOR2_X1   g667(.A1(new_n866_), .A2(new_n344_), .ZN(new_n869_));
  AOI21_X1  g668(.A(G183gat), .B1(new_n869_), .B2(new_n865_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n866_), .A2(new_n408_), .A3(new_n344_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n870_), .B1(new_n863_), .B2(new_n871_), .ZN(G1350gat));
  NAND4_X1  g671(.A1(new_n853_), .A2(new_n509_), .A3(new_n328_), .A4(new_n856_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT122), .ZN(new_n874_));
  AND3_X1   g673(.A1(new_n873_), .A2(new_n874_), .A3(G190gat), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n874_), .B1(new_n873_), .B2(G190gat), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n863_), .A2(new_n856_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n319_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n878_));
  XOR2_X1   g677(.A(new_n878_), .B(KEYINPUT123), .Z(new_n879_));
  OAI22_X1  g678(.A1(new_n875_), .A2(new_n876_), .B1(new_n877_), .B2(new_n879_), .ZN(G1351gat));
  INV_X1    g679(.A(KEYINPUT124), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n786_), .A2(new_n841_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n882_), .A2(new_n855_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(new_n281_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n881_), .B1(new_n884_), .B2(new_n276_), .ZN(new_n885_));
  NAND4_X1  g684(.A1(new_n883_), .A2(KEYINPUT124), .A3(G197gat), .A4(new_n281_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n884_), .A2(new_n276_), .ZN(new_n887_));
  AND3_X1   g686(.A1(new_n885_), .A2(new_n886_), .A3(new_n887_), .ZN(G1352gat));
  NAND2_X1  g687(.A1(new_n883_), .A2(new_n241_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g689(.A(new_n344_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n786_), .A2(new_n841_), .A3(new_n854_), .A4(new_n891_), .ZN(new_n892_));
  AND2_X1   g691(.A1(new_n892_), .A2(KEYINPUT125), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n892_), .A2(KEYINPUT125), .ZN(new_n894_));
  OR2_X1    g693(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n895_));
  OR3_X1    g694(.A1(new_n893_), .A2(new_n894_), .A3(new_n895_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n893_), .B2(new_n894_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(G1354gat));
  NOR2_X1   g697(.A1(new_n579_), .A2(new_n350_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(KEYINPUT126), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n883_), .A2(new_n900_), .ZN(new_n901_));
  NOR3_X1   g700(.A1(new_n882_), .A2(new_n318_), .A3(new_n855_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(G218gat), .B2(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT127), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n901_), .B(KEYINPUT127), .C1(G218gat), .C2(new_n902_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(G1355gat));
endmodule


