//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 1 1 0 0 0 1 1 1 1 1 1 1 0 0 1 0 1 0 1 1 1 1 1 0 1 0 1 1 1 0 1 0 0 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n669_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n692_,
    new_n693_, new_n694_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n845_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n873_, new_n874_, new_n875_,
    new_n877_, new_n878_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_;
  XOR2_X1   g000(.A(G22gat), .B(G50gat), .Z(new_n202_));
  INV_X1    g001(.A(KEYINPUT85), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G141gat), .A2(G148gat), .ZN(new_n209_));
  AND2_X1   g008(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n210_));
  NOR2_X1   g009(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n209_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT82), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n212_), .B(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT3), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G141gat), .A2(G148gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT2), .ZN(new_n217_));
  OAI22_X1  g016(.A1(new_n209_), .A2(new_n215_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT83), .ZN(new_n219_));
  INV_X1    g018(.A(new_n216_), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n219_), .B1(new_n220_), .B2(KEYINPUT2), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n216_), .A2(KEYINPUT83), .A3(new_n217_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n218_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n214_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT84), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n214_), .A2(KEYINPUT84), .A3(new_n223_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n208_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n206_), .B1(KEYINPUT1), .B2(new_n204_), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n204_), .A2(KEYINPUT1), .ZN(new_n230_));
  AOI211_X1 g029(.A(new_n209_), .B(new_n220_), .C1(new_n229_), .C2(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n203_), .B1(new_n228_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n227_), .ZN(new_n233_));
  AOI21_X1  g032(.A(KEYINPUT84), .B1(new_n214_), .B2(new_n223_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n207_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n231_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(KEYINPUT85), .A3(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n232_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT29), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT86), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT28), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT86), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n238_), .A2(new_n243_), .A3(new_n239_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n241_), .A2(new_n242_), .A3(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n242_), .B1(new_n241_), .B2(new_n244_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n202_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n241_), .A2(new_n244_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT28), .ZN(new_n250_));
  INV_X1    g049(.A(new_n202_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n250_), .A2(new_n245_), .A3(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT87), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n253_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G228gat), .A2(G233gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G211gat), .B(G218gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G197gat), .B(G204gat), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT21), .ZN(new_n258_));
  NOR4_X1   g057(.A1(new_n256_), .A2(new_n257_), .A3(KEYINPUT88), .A4(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT88), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n257_), .A2(new_n258_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n256_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n260_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  AND2_X1   g062(.A1(new_n257_), .A2(new_n258_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n256_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n265_));
  OAI22_X1  g064(.A1(new_n259_), .A2(new_n263_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n232_), .A2(new_n237_), .A3(KEYINPUT87), .A4(KEYINPUT29), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n254_), .A2(new_n255_), .A3(new_n266_), .A4(new_n267_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n228_), .A2(new_n231_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(KEYINPUT89), .B(KEYINPUT29), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n266_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n271_), .A2(G228gat), .A3(G233gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G78gat), .B(G106gat), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n268_), .A2(new_n272_), .A3(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(KEYINPUT90), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n248_), .A2(new_n252_), .A3(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n268_), .A2(new_n272_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(new_n273_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(new_n275_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n277_), .A2(new_n281_), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n280_), .A2(new_n276_), .A3(new_n252_), .A4(new_n248_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(KEYINPUT25), .B(G183gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT26), .B(G190gat), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT24), .ZN(new_n287_));
  NOR2_X1   g086(.A1(G169gat), .A2(G176gat), .ZN(new_n288_));
  AOI22_X1  g087(.A1(new_n285_), .A2(new_n286_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G169gat), .A2(G176gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(KEYINPUT24), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n289_), .B1(new_n288_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(G183gat), .ZN(new_n293_));
  INV_X1    g092(.A(G190gat), .ZN(new_n294_));
  OAI21_X1  g093(.A(KEYINPUT78), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT78), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n296_), .A2(G183gat), .A3(G190gat), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT23), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n295_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n292_), .A2(new_n301_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(G183gat), .A2(G190gat), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n295_), .A2(new_n297_), .A3(KEYINPUT23), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n298_), .A2(G183gat), .A3(G190gat), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n303_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT79), .ZN(new_n307_));
  OR2_X1    g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  XOR2_X1   g107(.A(KEYINPUT22), .B(G169gat), .Z(new_n309_));
  OAI21_X1  g108(.A(new_n290_), .B1(new_n309_), .B2(G176gat), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n310_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n302_), .B1(new_n308_), .B2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT30), .ZN(new_n313_));
  XOR2_X1   g112(.A(G71gat), .B(G99gat), .Z(new_n314_));
  NAND2_X1  g113(.A1(G227gat), .A2(G233gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G15gat), .B(G43gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT80), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n316_), .B(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n313_), .B(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT31), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G127gat), .B(G134gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G113gat), .B(G120gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n321_), .B(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n232_), .A2(new_n237_), .A3(new_n325_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n269_), .A2(new_n324_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G225gat), .A2(G233gat), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n327_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT95), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT95), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n327_), .A2(new_n328_), .A3(new_n332_), .A4(new_n329_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n238_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n324_), .A2(KEYINPUT4), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n329_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n327_), .A2(KEYINPUT4), .A3(new_n328_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n337_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n334_), .A2(new_n340_), .ZN(new_n341_));
  XOR2_X1   g140(.A(G1gat), .B(G29gat), .Z(new_n342_));
  XNOR2_X1  g141(.A(G57gat), .B(G85gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n345_));
  XOR2_X1   g144(.A(new_n344_), .B(new_n345_), .Z(new_n346_));
  NAND2_X1  g145(.A1(new_n341_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n346_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n334_), .A2(new_n348_), .A3(new_n340_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n347_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n326_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT27), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G226gat), .A2(G233gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT19), .ZN(new_n355_));
  OAI221_X1 g154(.A(new_n290_), .B1(G176gat), .B2(new_n309_), .C1(new_n301_), .C2(new_n303_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n304_), .A2(new_n305_), .ZN(new_n357_));
  XOR2_X1   g156(.A(new_n291_), .B(KEYINPUT91), .Z(new_n358_));
  OAI211_X1 g157(.A(new_n357_), .B(new_n289_), .C1(new_n358_), .C2(new_n288_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n356_), .A2(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT97), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n361_), .A2(new_n266_), .ZN(new_n362_));
  AND2_X1   g161(.A1(new_n308_), .A2(new_n311_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n266_), .B1(new_n363_), .B2(new_n302_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(KEYINPUT20), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n355_), .B1(new_n362_), .B2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n266_), .A2(new_n356_), .A3(new_n359_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n367_), .B1(new_n312_), .B2(new_n266_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT20), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n366_), .B1(new_n355_), .B2(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G8gat), .B(G36gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT18), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G64gat), .B(G92gat), .ZN(new_n373_));
  XOR2_X1   g172(.A(new_n372_), .B(new_n373_), .Z(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n353_), .B1(new_n370_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n355_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n377_), .B1(new_n360_), .B2(new_n266_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n365_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT92), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n381_), .B1(new_n369_), .B2(new_n355_), .ZN(new_n382_));
  AOI211_X1 g181(.A(KEYINPUT92), .B(new_n377_), .C1(new_n368_), .C2(KEYINPUT20), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n374_), .B(new_n380_), .C1(new_n382_), .C2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n376_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT93), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n369_), .A2(new_n355_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT92), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n369_), .A2(new_n381_), .A3(new_n355_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n379_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(KEYINPUT93), .B1(new_n391_), .B2(new_n374_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n387_), .B1(new_n392_), .B2(new_n384_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n385_), .B1(new_n393_), .B2(KEYINPUT27), .ZN(new_n394_));
  NOR3_X1   g193(.A1(new_n284_), .A2(new_n352_), .A3(new_n394_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n282_), .A2(new_n283_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n327_), .A2(new_n328_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n346_), .B1(new_n397_), .B2(new_n329_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n338_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n398_), .B1(new_n339_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT33), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n400_), .B1(new_n349_), .B2(new_n401_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n334_), .A2(KEYINPUT33), .A3(new_n348_), .A4(new_n340_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n402_), .A2(new_n393_), .A3(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT96), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n402_), .A2(new_n393_), .A3(KEYINPUT96), .A4(new_n403_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n370_), .A2(KEYINPUT32), .A3(new_n374_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT32), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n391_), .B1(new_n409_), .B2(new_n375_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n350_), .A2(new_n408_), .A3(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n407_), .A2(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n396_), .B1(new_n406_), .B2(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n394_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(new_n351_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n326_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n395_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT72), .B(G1gat), .ZN(new_n419_));
  INV_X1    g218(.A(G8gat), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT14), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G15gat), .B(G22gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G1gat), .B(G8gat), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n423_), .A2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n421_), .A2(new_n422_), .A3(new_n424_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G29gat), .B(G36gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G43gat), .B(G50gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n429_), .B(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n428_), .B(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n432_), .A2(G229gat), .A3(G233gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n431_), .B(KEYINPUT15), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n434_), .A2(new_n427_), .A3(new_n426_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n428_), .A2(new_n431_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G229gat), .A2(G233gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(KEYINPUT76), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n435_), .A2(new_n436_), .A3(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n433_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G113gat), .B(G141gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G169gat), .B(G197gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n441_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n440_), .A2(new_n444_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT77), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n446_), .A2(KEYINPUT77), .A3(new_n447_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT12), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT9), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G85gat), .B(G92gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(KEYINPUT10), .B(G99gat), .ZN(new_n457_));
  OAI22_X1  g256(.A1(new_n455_), .A2(new_n456_), .B1(new_n457_), .B2(G106gat), .ZN(new_n458_));
  AND3_X1   g257(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n459_));
  AOI21_X1  g258(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  AND2_X1   g260(.A1(G85gat), .A2(G92gat), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n461_), .B1(KEYINPUT9), .B2(new_n463_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n458_), .A2(new_n464_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(G85gat), .A2(G92gat), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n462_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT65), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT7), .ZN(new_n469_));
  INV_X1    g268(.A(G99gat), .ZN(new_n470_));
  INV_X1    g269(.A(G106gat), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n468_), .A2(new_n469_), .A3(new_n470_), .A4(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G99gat), .A2(G106gat), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT6), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n472_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(KEYINPUT65), .A2(G99gat), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n469_), .B1(new_n478_), .B2(new_n471_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n467_), .B1(new_n477_), .B2(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(KEYINPUT8), .B1(new_n467_), .B2(KEYINPUT66), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n468_), .A2(new_n470_), .A3(new_n471_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT7), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n485_), .A2(new_n461_), .A3(new_n472_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n486_), .A2(new_n467_), .A3(new_n481_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n465_), .B1(new_n483_), .B2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G57gat), .B(G64gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(KEYINPUT11), .ZN(new_n490_));
  XOR2_X1   g289(.A(G71gat), .B(G78gat), .Z(new_n491_));
  NOR2_X1   g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n490_), .A2(new_n491_), .ZN(new_n493_));
  OR2_X1    g292(.A1(new_n489_), .A2(KEYINPUT11), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n492_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n454_), .B1(new_n488_), .B2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT68), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  OR2_X1    g298(.A1(new_n458_), .A2(new_n464_), .ZN(new_n500_));
  AND3_X1   g299(.A1(new_n486_), .A2(new_n467_), .A3(new_n481_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n481_), .B1(new_n486_), .B2(new_n467_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n500_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(new_n495_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n504_), .A2(KEYINPUT68), .A3(new_n454_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n499_), .A2(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n503_), .A2(KEYINPUT12), .A3(new_n495_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT67), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n503_), .A2(KEYINPUT67), .A3(KEYINPUT12), .A4(new_n495_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G230gat), .A2(G233gat), .ZN(new_n512_));
  XOR2_X1   g311(.A(new_n512_), .B(KEYINPUT64), .Z(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n488_), .A2(new_n496_), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n506_), .A2(new_n511_), .A3(new_n514_), .A4(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n504_), .A2(new_n515_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(new_n513_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  XOR2_X1   g318(.A(G120gat), .B(G148gat), .Z(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT5), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G176gat), .B(G204gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n519_), .B(new_n523_), .ZN(new_n524_));
  OR2_X1    g323(.A1(new_n524_), .A2(KEYINPUT13), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(KEYINPUT13), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G232gat), .A2(G233gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT34), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT35), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT70), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n434_), .A2(new_n503_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT69), .ZN(new_n536_));
  AOI22_X1  g335(.A1(new_n488_), .A2(new_n431_), .B1(new_n531_), .B2(new_n530_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n534_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n532_), .A2(new_n533_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n536_), .A2(new_n533_), .A3(new_n537_), .A4(new_n532_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  XOR2_X1   g341(.A(G190gat), .B(G218gat), .Z(new_n543_));
  XNOR2_X1  g342(.A(G134gat), .B(G162gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n546_), .A2(KEYINPUT36), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n542_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT71), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n545_), .B(KEYINPUT36), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n540_), .A2(new_n541_), .A3(new_n550_), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n548_), .A2(new_n549_), .A3(KEYINPUT37), .A4(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT37), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n548_), .A2(new_n551_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n553_), .B1(new_n554_), .B2(KEYINPUT71), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G231gat), .A2(G233gat), .ZN(new_n556_));
  XOR2_X1   g355(.A(new_n556_), .B(KEYINPUT73), .Z(new_n557_));
  XNOR2_X1  g356(.A(new_n495_), .B(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(new_n428_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G127gat), .B(G155gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT16), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G183gat), .B(G211gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(KEYINPUT17), .B1(new_n559_), .B2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT74), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n563_), .B1(new_n559_), .B2(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n564_), .B(new_n566_), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n527_), .A2(new_n552_), .A3(new_n555_), .A4(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n568_), .B(KEYINPUT75), .Z(new_n569_));
  NOR3_X1   g368(.A1(new_n418_), .A2(new_n453_), .A3(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n570_), .A2(new_n350_), .A3(new_n419_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT38), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n573_), .B(KEYINPUT98), .Z(new_n574_));
  NAND2_X1  g373(.A1(new_n571_), .A2(new_n572_), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n575_), .B(KEYINPUT99), .Z(new_n576_));
  INV_X1    g375(.A(new_n395_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n404_), .A2(new_n405_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n578_), .A2(new_n407_), .A3(new_n411_), .ZN(new_n579_));
  AOI22_X1  g378(.A1(new_n579_), .A2(new_n396_), .B1(new_n414_), .B2(new_n351_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n577_), .B1(new_n580_), .B2(new_n326_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n527_), .A2(new_n452_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n567_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n581_), .A2(new_n554_), .A3(new_n584_), .ZN(new_n585_));
  OAI21_X1  g384(.A(G1gat), .B1(new_n585_), .B2(new_n351_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n574_), .A2(new_n576_), .A3(new_n586_), .ZN(G1324gat));
  INV_X1    g386(.A(KEYINPUT40), .ZN(new_n588_));
  INV_X1    g387(.A(new_n394_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n589_), .A2(G8gat), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n570_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT100), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n585_), .A2(new_n589_), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n594_), .A2(KEYINPUT101), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n420_), .B1(new_n594_), .B2(KEYINPUT101), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n595_), .A2(KEYINPUT39), .A3(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n593_), .A2(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(KEYINPUT39), .B1(new_n595_), .B2(new_n596_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n588_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n599_), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n601_), .A2(KEYINPUT40), .A3(new_n597_), .A4(new_n593_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(G1325gat));
  OAI21_X1  g402(.A(G15gat), .B1(new_n585_), .B2(new_n417_), .ZN(new_n604_));
  OR2_X1    g403(.A1(new_n604_), .A2(KEYINPUT41), .ZN(new_n605_));
  INV_X1    g404(.A(G15gat), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n570_), .A2(new_n606_), .A3(new_n326_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n604_), .A2(KEYINPUT41), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n605_), .A2(new_n607_), .A3(new_n608_), .ZN(G1326gat));
  XNOR2_X1  g408(.A(new_n396_), .B(KEYINPUT102), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  OAI21_X1  g410(.A(G22gat), .B1(new_n585_), .B2(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT42), .ZN(new_n613_));
  INV_X1    g412(.A(G22gat), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n570_), .A2(new_n614_), .A3(new_n610_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n613_), .A2(new_n615_), .ZN(G1327gat));
  NOR3_X1   g415(.A1(new_n582_), .A2(new_n554_), .A3(new_n567_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n581_), .A2(new_n617_), .ZN(new_n618_));
  OR3_X1    g417(.A1(new_n618_), .A2(G29gat), .A3(new_n351_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n582_), .A2(new_n567_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT43), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n555_), .A2(new_n552_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n326_), .B1(new_n413_), .B2(new_n415_), .ZN(new_n623_));
  OAI211_X1 g422(.A(new_n621_), .B(new_n622_), .C1(new_n623_), .C2(new_n395_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n621_), .B1(new_n581_), .B2(new_n622_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n620_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT44), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n622_), .ZN(new_n630_));
  OAI21_X1  g429(.A(KEYINPUT43), .B1(new_n418_), .B2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(new_n624_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n632_), .A2(KEYINPUT44), .A3(new_n620_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n629_), .A2(new_n350_), .A3(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT103), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n634_), .A2(new_n635_), .A3(G29gat), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n635_), .B1(new_n634_), .B2(G29gat), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n619_), .B1(new_n636_), .B2(new_n637_), .ZN(G1328gat));
  INV_X1    g437(.A(KEYINPUT105), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT46), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  XOR2_X1   g440(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n642_));
  NOR2_X1   g441(.A1(new_n589_), .A2(G36gat), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n642_), .B1(new_n618_), .B2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n642_), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n581_), .A2(new_n617_), .A3(new_n643_), .A4(new_n646_), .ZN(new_n647_));
  AOI22_X1  g446(.A1(new_n645_), .A2(new_n647_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n629_), .A2(new_n394_), .A3(new_n633_), .ZN(new_n650_));
  AOI211_X1 g449(.A(new_n641_), .B(new_n649_), .C1(new_n650_), .C2(G36gat), .ZN(new_n651_));
  INV_X1    g450(.A(new_n641_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n620_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n653_), .B1(new_n631_), .B2(new_n624_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n394_), .B1(new_n654_), .B2(KEYINPUT44), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n627_), .A2(new_n628_), .ZN(new_n656_));
  OAI21_X1  g455(.A(G36gat), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n652_), .B1(new_n657_), .B2(new_n648_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n651_), .A2(new_n658_), .ZN(G1329gat));
  INV_X1    g458(.A(G43gat), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n660_), .B1(new_n618_), .B2(new_n417_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT106), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n629_), .A2(G43gat), .A3(new_n326_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n662_), .B1(new_n663_), .B2(new_n656_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(KEYINPUT47), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT47), .ZN(new_n666_));
  OAI211_X1 g465(.A(new_n662_), .B(new_n666_), .C1(new_n663_), .C2(new_n656_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(G1330gat));
  INV_X1    g467(.A(new_n618_), .ZN(new_n669_));
  AOI21_X1  g468(.A(G50gat), .B1(new_n669_), .B2(new_n610_), .ZN(new_n670_));
  AND3_X1   g469(.A1(new_n629_), .A2(G50gat), .A3(new_n284_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n670_), .B1(new_n671_), .B2(new_n633_), .ZN(G1331gat));
  NOR2_X1   g471(.A1(new_n527_), .A2(new_n452_), .ZN(new_n673_));
  NAND4_X1  g472(.A1(new_n581_), .A2(new_n554_), .A3(new_n567_), .A4(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(G57gat), .B1(new_n674_), .B2(new_n351_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n673_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n418_), .A2(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n622_), .A2(new_n583_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  OR2_X1    g478(.A1(new_n351_), .A2(G57gat), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n675_), .B1(new_n679_), .B2(new_n680_), .ZN(G1332gat));
  OAI21_X1  g480(.A(G64gat), .B1(new_n674_), .B2(new_n589_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT48), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n589_), .A2(G64gat), .ZN(new_n684_));
  XOR2_X1   g483(.A(new_n684_), .B(KEYINPUT107), .Z(new_n685_));
  OAI21_X1  g484(.A(new_n683_), .B1(new_n679_), .B2(new_n685_), .ZN(G1333gat));
  OAI21_X1  g485(.A(G71gat), .B1(new_n674_), .B2(new_n417_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT49), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n417_), .A2(G71gat), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n689_), .B(KEYINPUT108), .Z(new_n690_));
  OAI21_X1  g489(.A(new_n688_), .B1(new_n679_), .B2(new_n690_), .ZN(G1334gat));
  OAI21_X1  g490(.A(G78gat), .B1(new_n674_), .B2(new_n611_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT50), .ZN(new_n693_));
  OR2_X1    g492(.A1(new_n611_), .A2(G78gat), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n693_), .B1(new_n679_), .B2(new_n694_), .ZN(G1335gat));
  NOR2_X1   g494(.A1(new_n676_), .A2(new_n567_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n632_), .A2(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(G85gat), .B1(new_n697_), .B2(new_n351_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n554_), .A2(new_n567_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n677_), .A2(new_n699_), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n351_), .A2(G85gat), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n698_), .B1(new_n700_), .B2(new_n701_), .ZN(G1336gat));
  OAI21_X1  g501(.A(G92gat), .B1(new_n697_), .B2(new_n589_), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n589_), .A2(G92gat), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n703_), .B1(new_n700_), .B2(new_n704_), .ZN(G1337gat));
  NOR3_X1   g504(.A1(new_n700_), .A2(new_n417_), .A3(new_n457_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n706_), .A2(KEYINPUT110), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n326_), .B(new_n696_), .C1(new_n625_), .C2(new_n626_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT109), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n708_), .A2(new_n709_), .A3(G99gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n709_), .B1(new_n708_), .B2(G99gat), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n707_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT51), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT51), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n707_), .B(new_n714_), .C1(new_n710_), .C2(new_n711_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(G1338gat));
  NAND4_X1  g515(.A1(new_n677_), .A2(new_n471_), .A3(new_n284_), .A4(new_n699_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT111), .ZN(new_n718_));
  OAI211_X1 g517(.A(new_n284_), .B(new_n696_), .C1(new_n625_), .C2(new_n626_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(G106gat), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT52), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n719_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n718_), .A2(new_n722_), .A3(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(KEYINPUT53), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT53), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n718_), .A2(new_n722_), .A3(new_n726_), .A4(new_n723_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(G1339gat));
  INV_X1    g527(.A(KEYINPUT112), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n729_), .B(KEYINPUT54), .C1(new_n568_), .C2(new_n452_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n678_), .A2(new_n453_), .A3(new_n527_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n730_), .B1(new_n731_), .B2(KEYINPUT54), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n729_), .B1(new_n731_), .B2(KEYINPUT54), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n519_), .A2(new_n523_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n435_), .A2(new_n436_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT114), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n737_), .A2(new_n438_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n445_), .B1(new_n432_), .B2(new_n438_), .ZN(new_n739_));
  AOI22_X1  g538(.A1(new_n738_), .A2(new_n739_), .B1(new_n441_), .B2(new_n445_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT55), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n516_), .A2(new_n741_), .ZN(new_n742_));
  AOI22_X1  g541(.A1(new_n499_), .A2(new_n505_), .B1(new_n488_), .B2(new_n496_), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n743_), .A2(KEYINPUT55), .A3(new_n514_), .A4(new_n511_), .ZN(new_n744_));
  AOI21_X1  g543(.A(KEYINPUT68), .B1(new_n504_), .B2(new_n454_), .ZN(new_n745_));
  AOI211_X1 g544(.A(new_n498_), .B(KEYINPUT12), .C1(new_n503_), .C2(new_n495_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n515_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n509_), .A2(new_n510_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n513_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n742_), .A2(new_n744_), .A3(new_n749_), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n750_), .A2(KEYINPUT56), .A3(new_n523_), .ZN(new_n751_));
  AOI21_X1  g550(.A(KEYINPUT56), .B1(new_n750_), .B2(new_n523_), .ZN(new_n752_));
  OAI211_X1 g551(.A(new_n735_), .B(new_n740_), .C1(new_n751_), .C2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT58), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n753_), .A2(KEYINPUT115), .A3(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n750_), .A2(new_n523_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT56), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n750_), .A2(KEYINPUT56), .A3(new_n523_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n754_), .A2(KEYINPUT115), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n760_), .A2(new_n735_), .A3(new_n740_), .A4(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n755_), .A2(new_n622_), .A3(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n554_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n524_), .A2(new_n740_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  OAI211_X1 g565(.A(new_n452_), .B(new_n735_), .C1(new_n751_), .C2(new_n752_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT113), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n766_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n760_), .A2(KEYINPUT113), .A3(new_n452_), .A4(new_n735_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n764_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n763_), .B1(new_n771_), .B2(KEYINPUT57), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n767_), .A2(new_n768_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n773_), .A2(new_n770_), .A3(new_n765_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n774_), .A2(KEYINPUT57), .A3(new_n554_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT116), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n771_), .A2(KEYINPUT116), .A3(KEYINPUT57), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n772_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n734_), .B1(new_n567_), .B2(new_n779_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n284_), .A2(new_n394_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n781_), .A2(new_n326_), .A3(new_n350_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n780_), .A2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT59), .ZN(new_n785_));
  OAI21_X1  g584(.A(KEYINPUT118), .B1(new_n779_), .B2(new_n567_), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n755_), .A2(new_n622_), .A3(new_n762_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n774_), .A2(new_n554_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT57), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n787_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  AND4_X1   g589(.A1(KEYINPUT116), .A2(new_n774_), .A3(KEYINPUT57), .A4(new_n554_), .ZN(new_n791_));
  AOI21_X1  g590(.A(KEYINPUT116), .B1(new_n771_), .B2(KEYINPUT57), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n790_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT118), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n793_), .A2(new_n794_), .A3(new_n583_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n786_), .A2(new_n734_), .A3(new_n795_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n782_), .A2(KEYINPUT59), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n785_), .A2(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(G113gat), .B1(new_n799_), .B2(new_n453_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n732_), .A2(new_n733_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n801_), .B1(new_n583_), .B2(new_n793_), .ZN(new_n802_));
  OAI21_X1  g601(.A(KEYINPUT117), .B1(new_n802_), .B2(new_n782_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT117), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n780_), .A2(new_n804_), .A3(new_n783_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n805_), .ZN(new_n806_));
  OR2_X1    g605(.A1(new_n453_), .A2(G113gat), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n800_), .B1(new_n806_), .B2(new_n807_), .ZN(G1340gat));
  OAI21_X1  g607(.A(G120gat), .B1(new_n799_), .B2(new_n527_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n527_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT60), .ZN(new_n811_));
  INV_X1    g610(.A(G120gat), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n810_), .A2(new_n811_), .A3(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n813_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n803_), .A2(new_n805_), .A3(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n809_), .A2(KEYINPUT119), .A3(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT119), .ZN(new_n817_));
  AOI22_X1  g616(.A1(new_n784_), .A2(KEYINPUT59), .B1(new_n796_), .B2(new_n797_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n812_), .B1(new_n818_), .B2(new_n810_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n815_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n817_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n816_), .A2(new_n821_), .ZN(G1341gat));
  INV_X1    g621(.A(G127gat), .ZN(new_n823_));
  NOR3_X1   g622(.A1(new_n799_), .A2(new_n823_), .A3(new_n583_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n803_), .A2(new_n805_), .A3(new_n567_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT120), .ZN(new_n826_));
  AND3_X1   g625(.A1(new_n825_), .A2(new_n826_), .A3(new_n823_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n826_), .B1(new_n825_), .B2(new_n823_), .ZN(new_n828_));
  NOR3_X1   g627(.A1(new_n824_), .A2(new_n827_), .A3(new_n828_), .ZN(G1342gat));
  INV_X1    g628(.A(G134gat), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n830_), .B1(new_n806_), .B2(new_n554_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n622_), .A2(G134gat), .ZN(new_n832_));
  XOR2_X1   g631(.A(new_n832_), .B(KEYINPUT121), .Z(new_n833_));
  NAND2_X1  g632(.A1(new_n818_), .A2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n831_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT122), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n831_), .A2(new_n834_), .A3(KEYINPUT122), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(G1343gat));
  AND3_X1   g638(.A1(new_n414_), .A2(new_n417_), .A3(new_n350_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n780_), .A2(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n841_), .A2(new_n453_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(KEYINPUT123), .B(G141gat), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n842_), .B(new_n843_), .ZN(G1344gat));
  NOR2_X1   g643(.A1(new_n841_), .A2(new_n527_), .ZN(new_n845_));
  XOR2_X1   g644(.A(new_n845_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g645(.A1(new_n841_), .A2(new_n583_), .ZN(new_n847_));
  XOR2_X1   g646(.A(KEYINPUT61), .B(G155gat), .Z(new_n848_));
  XNOR2_X1  g647(.A(new_n847_), .B(new_n848_), .ZN(G1346gat));
  OAI21_X1  g648(.A(G162gat), .B1(new_n841_), .B2(new_n630_), .ZN(new_n850_));
  OR2_X1    g649(.A1(new_n554_), .A2(G162gat), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n850_), .B1(new_n841_), .B2(new_n851_), .ZN(G1347gat));
  NOR2_X1   g651(.A1(new_n352_), .A2(new_n589_), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n796_), .A2(new_n853_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n453_), .A2(new_n309_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(KEYINPUT125), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n854_), .A2(new_n611_), .A3(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT62), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n610_), .A2(new_n453_), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n796_), .A2(KEYINPUT124), .A3(new_n853_), .A4(new_n859_), .ZN(new_n860_));
  AND2_X1   g659(.A1(new_n860_), .A2(G169gat), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n796_), .A2(new_n853_), .A3(new_n859_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT124), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n858_), .B1(new_n861_), .B2(new_n864_), .ZN(new_n865_));
  AND4_X1   g664(.A1(new_n858_), .A2(new_n864_), .A3(G169gat), .A4(new_n860_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n857_), .B1(new_n865_), .B2(new_n866_), .ZN(G1348gat));
  NOR2_X1   g666(.A1(new_n802_), .A2(new_n284_), .ZN(new_n868_));
  AND4_X1   g667(.A1(G176gat), .A2(new_n868_), .A3(new_n810_), .A4(new_n853_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n854_), .A2(new_n810_), .A3(new_n611_), .ZN(new_n870_));
  INV_X1    g669(.A(G176gat), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n869_), .B1(new_n870_), .B2(new_n871_), .ZN(G1349gat));
  NAND2_X1  g671(.A1(new_n854_), .A2(new_n611_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n873_), .A2(new_n285_), .A3(new_n583_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n868_), .A2(new_n567_), .A3(new_n853_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n874_), .B1(new_n293_), .B2(new_n875_), .ZN(G1350gat));
  OAI21_X1  g675(.A(G190gat), .B1(new_n873_), .B2(new_n630_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n764_), .A2(new_n286_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n873_), .B2(new_n878_), .ZN(G1351gat));
  INV_X1    g678(.A(KEYINPUT126), .ZN(new_n880_));
  NOR4_X1   g679(.A1(new_n396_), .A2(new_n589_), .A3(new_n326_), .A4(new_n350_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n880_), .B1(new_n802_), .B2(new_n882_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n780_), .A2(KEYINPUT126), .A3(new_n881_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n452_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g686(.A1(new_n885_), .A2(new_n810_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g688(.A(new_n583_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n891_));
  AND2_X1   g690(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n890_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n893_), .B1(new_n890_), .B2(new_n891_), .ZN(G1354gat));
  AND2_X1   g693(.A1(new_n622_), .A2(G218gat), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n885_), .A2(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n554_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(G218gat), .B2(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT127), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  OAI211_X1 g699(.A(new_n896_), .B(KEYINPUT127), .C1(G218gat), .C2(new_n897_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(G1355gat));
endmodule


