//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 0 1 0 1 1 1 0 1 1 1 0 0 1 1 1 1 1 0 1 0 1 0 0 1 0 0 0 1 0 1 0 0 1 1 1 0 0 1 0 1 0 0 1 0 1 1 1 1 0 1 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n637_, new_n638_, new_n639_, new_n640_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n749_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n872_, new_n873_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n881_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n916_, new_n917_,
    new_n918_, new_n920_, new_n921_, new_n923_, new_n924_, new_n925_,
    new_n927_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_;
  XNOR2_X1  g000(.A(G71gat), .B(G99gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G15gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT80), .B(G43gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G227gat), .A2(G233gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT26), .B(G190gat), .ZN(new_n208_));
  INV_X1    g007(.A(G183gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT25), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT76), .B1(new_n209_), .B2(KEYINPUT25), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT76), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT25), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n212_), .A2(new_n213_), .A3(G183gat), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n208_), .A2(new_n210_), .A3(new_n211_), .A4(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT77), .ZN(new_n216_));
  OR2_X1    g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(new_n216_), .ZN(new_n218_));
  OR2_X1    g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n219_), .A2(KEYINPUT24), .ZN(new_n220_));
  INV_X1    g019(.A(G190gat), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT23), .B1(new_n209_), .B2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT23), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(G183gat), .A3(G190gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n222_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n219_), .A2(KEYINPUT24), .A3(new_n226_), .ZN(new_n227_));
  AND3_X1   g026(.A1(new_n220_), .A2(new_n225_), .A3(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n217_), .A2(new_n218_), .A3(new_n228_), .ZN(new_n229_));
  XOR2_X1   g028(.A(KEYINPUT78), .B(G176gat), .Z(new_n230_));
  XNOR2_X1  g029(.A(KEYINPUT22), .B(G169gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n222_), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n224_), .A2(KEYINPUT79), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n224_), .A2(KEYINPUT79), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n233_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(G183gat), .A2(G190gat), .ZN(new_n237_));
  OAI211_X1 g036(.A(new_n226_), .B(new_n232_), .C1(new_n236_), .C2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n229_), .A2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT30), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT81), .ZN(new_n241_));
  AND2_X1   g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n240_), .A2(new_n241_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n207_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n244_), .B1(new_n242_), .B2(new_n207_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G127gat), .B(G134gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G113gat), .B(G120gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  XOR2_X1   g047(.A(KEYINPUT82), .B(KEYINPUT31), .Z(new_n249_));
  XOR2_X1   g048(.A(new_n248_), .B(new_n249_), .Z(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n245_), .B(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT91), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G228gat), .A2(G233gat), .ZN(new_n254_));
  NOR2_X1   g053(.A1(G155gat), .A2(G162gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G155gat), .A2(G162gat), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n255_), .B1(KEYINPUT1), .B2(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n257_), .B1(KEYINPUT1), .B2(new_n256_), .ZN(new_n258_));
  XOR2_X1   g057(.A(G141gat), .B(G148gat), .Z(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  AND3_X1   g059(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n261_));
  AOI21_X1  g060(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  OAI22_X1  g062(.A1(KEYINPUT83), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(KEYINPUT83), .A2(KEYINPUT3), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  OAI211_X1 g065(.A(KEYINPUT83), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n263_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT84), .ZN(new_n269_));
  XOR2_X1   g068(.A(G155gat), .B(G162gat), .Z(new_n270_));
  AND3_X1   g069(.A1(new_n268_), .A2(new_n269_), .A3(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n269_), .B1(new_n268_), .B2(new_n270_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n260_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT29), .ZN(new_n274_));
  INV_X1    g073(.A(G197gat), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n275_), .A2(G204gat), .ZN(new_n276_));
  INV_X1    g075(.A(G204gat), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n277_), .A2(G197gat), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT21), .B1(new_n276_), .B2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT89), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G211gat), .B(G218gat), .ZN(new_n281_));
  OR3_X1    g080(.A1(new_n279_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n280_), .B1(new_n279_), .B2(new_n281_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G197gat), .B(G204gat), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT21), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n287_), .A2(new_n279_), .A3(new_n281_), .ZN(new_n288_));
  AND2_X1   g087(.A1(new_n288_), .A2(KEYINPUT88), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n288_), .A2(KEYINPUT88), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n284_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n254_), .B1(new_n274_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT85), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n268_), .A2(new_n270_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(KEYINPUT84), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n268_), .A2(new_n269_), .A3(new_n270_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n293_), .B1(new_n297_), .B2(new_n260_), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n293_), .B(new_n260_), .C1(new_n271_), .C2(new_n272_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT29), .B1(new_n298_), .B2(new_n300_), .ZN(new_n301_));
  XOR2_X1   g100(.A(new_n254_), .B(KEYINPUT87), .Z(new_n302_));
  NAND2_X1  g101(.A1(new_n291_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n292_), .B1(new_n301_), .B2(new_n304_), .ZN(new_n305_));
  XOR2_X1   g104(.A(G78gat), .B(G106gat), .Z(new_n306_));
  OAI21_X1  g105(.A(new_n253_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n292_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT29), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n273_), .A2(KEYINPUT85), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n309_), .B1(new_n310_), .B2(new_n299_), .ZN(new_n311_));
  OAI211_X1 g110(.A(new_n308_), .B(new_n306_), .C1(new_n311_), .C2(new_n303_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n310_), .A2(new_n309_), .A3(new_n299_), .ZN(new_n313_));
  XOR2_X1   g112(.A(KEYINPUT86), .B(KEYINPUT28), .Z(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n314_), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n310_), .A2(new_n309_), .A3(new_n299_), .A4(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G22gat), .B(G50gat), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n315_), .A2(new_n319_), .A3(new_n317_), .ZN(new_n322_));
  AOI22_X1  g121(.A1(new_n307_), .A2(new_n312_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n305_), .A2(new_n253_), .A3(new_n306_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n306_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n310_), .A2(new_n299_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n303_), .B1(new_n327_), .B2(KEYINPUT29), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n326_), .B1(new_n328_), .B2(new_n292_), .ZN(new_n329_));
  AND2_X1   g128(.A1(new_n329_), .A2(new_n312_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n321_), .A2(new_n322_), .ZN(new_n331_));
  NOR3_X1   g130(.A1(new_n330_), .A2(new_n331_), .A3(KEYINPUT90), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT90), .ZN(new_n333_));
  INV_X1    g132(.A(new_n322_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n319_), .B1(new_n315_), .B2(new_n317_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n329_), .A2(new_n312_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n333_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n325_), .B1(new_n332_), .B2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G1gat), .B(G29gat), .ZN(new_n340_));
  INV_X1    g139(.A(G85gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT0), .B(G57gat), .ZN(new_n343_));
  XOR2_X1   g142(.A(new_n342_), .B(new_n343_), .Z(new_n344_));
  NAND2_X1  g143(.A1(G225gat), .A2(G233gat), .ZN(new_n345_));
  AOI22_X1  g144(.A1(new_n295_), .A2(new_n296_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n346_));
  AOI21_X1  g145(.A(KEYINPUT94), .B1(new_n346_), .B2(new_n248_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n248_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n347_), .B1(new_n327_), .B2(new_n348_), .ZN(new_n349_));
  AOI211_X1 g148(.A(KEYINPUT94), .B(new_n248_), .C1(new_n310_), .C2(new_n299_), .ZN(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT4), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n248_), .B1(new_n310_), .B2(new_n299_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n352_), .A2(KEYINPUT4), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n345_), .B1(new_n351_), .B2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n327_), .A2(new_n348_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n347_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT94), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n359_), .B(new_n348_), .C1(new_n298_), .C2(new_n300_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n358_), .A2(new_n345_), .A3(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n344_), .B1(new_n355_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n344_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n360_), .B1(new_n352_), .B2(new_n347_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n353_), .B1(new_n365_), .B2(KEYINPUT4), .ZN(new_n366_));
  OAI211_X1 g165(.A(new_n364_), .B(new_n361_), .C1(new_n366_), .C2(new_n345_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n363_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G226gat), .A2(G233gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT19), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT20), .ZN(new_n372_));
  INV_X1    g171(.A(new_n291_), .ZN(new_n373_));
  AND2_X1   g172(.A1(new_n229_), .A2(new_n238_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n372_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n288_), .B(KEYINPUT88), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n231_), .B(KEYINPUT93), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(new_n230_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n225_), .B1(G183gat), .B2(G190gat), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n378_), .A2(new_n226_), .A3(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n213_), .A2(G183gat), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n208_), .A2(new_n210_), .A3(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(new_n227_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT92), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n234_), .A2(new_n235_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(new_n222_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n382_), .A2(KEYINPUT92), .A3(new_n227_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n385_), .A2(new_n387_), .A3(new_n220_), .A4(new_n388_), .ZN(new_n389_));
  AOI22_X1  g188(.A1(new_n376_), .A2(new_n284_), .B1(new_n380_), .B2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n371_), .B1(new_n375_), .B2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n239_), .A2(new_n291_), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n376_), .A2(new_n380_), .A3(new_n389_), .A4(new_n284_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n393_), .A2(new_n394_), .A3(KEYINPUT20), .A4(new_n371_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n392_), .A2(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G8gat), .B(G36gat), .ZN(new_n398_));
  INV_X1    g197(.A(G92gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(KEYINPUT18), .B(G64gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n400_), .B(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT32), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(KEYINPUT95), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n397_), .A2(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT20), .B1(new_n239_), .B2(new_n291_), .ZN(new_n407_));
  NOR3_X1   g206(.A1(new_n407_), .A2(new_n390_), .A3(new_n370_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n393_), .A2(new_n394_), .A3(KEYINPUT20), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n408_), .B1(new_n370_), .B2(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n406_), .B1(new_n403_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n368_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT33), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n367_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n402_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n416_), .B1(new_n392_), .B2(new_n396_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n370_), .B1(new_n407_), .B2(new_n390_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n418_), .A2(new_n402_), .A3(new_n395_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT4), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n421_), .B1(new_n358_), .B2(new_n360_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n345_), .B1(new_n422_), .B2(new_n353_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n345_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n358_), .A2(new_n424_), .A3(new_n360_), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n425_), .A2(new_n344_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n420_), .B1(new_n423_), .B2(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n424_), .B1(new_n422_), .B2(new_n353_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n428_), .A2(KEYINPUT33), .A3(new_n364_), .A4(new_n361_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n415_), .A2(new_n427_), .A3(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n339_), .B1(new_n413_), .B2(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT90), .B1(new_n330_), .B2(new_n331_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n336_), .A2(new_n333_), .A3(new_n337_), .ZN(new_n433_));
  AOI22_X1  g232(.A1(new_n432_), .A2(new_n433_), .B1(new_n324_), .B2(new_n323_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT27), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n420_), .A2(new_n435_), .ZN(new_n436_));
  OAI211_X1 g235(.A(KEYINPUT27), .B(new_n419_), .C1(new_n410_), .C2(new_n402_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NOR3_X1   g237(.A1(new_n434_), .A2(new_n368_), .A3(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n252_), .B1(new_n431_), .B2(new_n439_), .ZN(new_n440_));
  NOR3_X1   g239(.A1(new_n252_), .A2(new_n339_), .A3(new_n368_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n438_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n440_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(G230gat), .A2(G233gat), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G99gat), .A2(G106gat), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT6), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n450_));
  AND2_X1   g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(KEYINPUT10), .B(G99gat), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n451_), .B1(G106gat), .B2(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(G85gat), .A2(G92gat), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT64), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G85gat), .A2(G92gat), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n455_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  OR2_X1    g257(.A1(new_n458_), .A2(KEYINPUT9), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n454_), .B1(new_n458_), .B2(KEYINPUT9), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n453_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT66), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NOR3_X1   g263(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n462_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT7), .ZN(new_n467_));
  INV_X1    g266(.A(G99gat), .ZN(new_n468_));
  INV_X1    g267(.A(G106gat), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n467_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n470_), .A2(KEYINPUT66), .A3(new_n463_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n466_), .A2(new_n451_), .A3(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n457_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n473_), .A2(new_n454_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT8), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n470_), .A2(new_n449_), .A3(new_n450_), .A4(new_n463_), .ZN(new_n477_));
  NOR3_X1   g276(.A1(new_n473_), .A2(new_n454_), .A3(KEYINPUT8), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n477_), .A2(KEYINPUT65), .A3(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(KEYINPUT65), .B1(new_n477_), .B2(new_n478_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n461_), .B1(new_n476_), .B2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G71gat), .B(G78gat), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G57gat), .A2(G64gat), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(G57gat), .A2(G64gat), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT11), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(G57gat), .ZN(new_n490_));
  INV_X1    g289(.A(G64gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT11), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n492_), .A2(new_n493_), .A3(new_n486_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n485_), .A2(new_n489_), .A3(new_n494_), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n484_), .B(KEYINPUT11), .C1(new_n488_), .C2(new_n487_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n483_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n459_), .A2(new_n460_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n453_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n481_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(new_n479_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT8), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n504_), .B1(new_n472_), .B2(new_n474_), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n501_), .B(new_n497_), .C1(new_n503_), .C2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n446_), .B1(new_n498_), .B2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT68), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n497_), .A2(KEYINPUT67), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT67), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n495_), .A2(new_n496_), .A3(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n510_), .A2(KEYINPUT12), .A3(new_n512_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n506_), .B1(new_n483_), .B2(new_n513_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n501_), .B1(new_n503_), .B2(new_n505_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n497_), .ZN(new_n516_));
  AOI21_X1  g315(.A(KEYINPUT12), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n514_), .A2(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n509_), .B1(new_n518_), .B2(new_n445_), .ZN(new_n519_));
  NOR4_X1   g318(.A1(new_n514_), .A2(new_n517_), .A3(KEYINPUT68), .A4(new_n446_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n508_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G120gat), .B(G148gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(new_n277_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(KEYINPUT5), .B(G176gat), .ZN(new_n524_));
  XOR2_X1   g323(.A(new_n523_), .B(new_n524_), .Z(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n521_), .A2(new_n526_), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n508_), .B(new_n525_), .C1(new_n519_), .C2(new_n520_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n529_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n527_), .A2(new_n528_), .A3(new_n530_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  XOR2_X1   g335(.A(G43gat), .B(G50gat), .Z(new_n537_));
  XNOR2_X1  g336(.A(G29gat), .B(G36gat), .ZN(new_n538_));
  OR2_X1    g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n537_), .A2(new_n538_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT73), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G15gat), .B(G22gat), .ZN(new_n543_));
  INV_X1    g342(.A(G1gat), .ZN(new_n544_));
  INV_X1    g343(.A(G8gat), .ZN(new_n545_));
  OAI21_X1  g344(.A(KEYINPUT14), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n543_), .A2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G1gat), .B(G8gat), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n547_), .B(new_n548_), .Z(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n542_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT15), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n541_), .B(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(new_n550_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n551_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G229gat), .A2(G233gat), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n542_), .A2(new_n550_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n556_), .B1(new_n551_), .B2(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G169gat), .B(G197gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT75), .ZN(new_n563_));
  XOR2_X1   g362(.A(G113gat), .B(G141gat), .Z(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT74), .ZN(new_n566_));
  OR2_X1    g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n561_), .B(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n536_), .A2(new_n569_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n444_), .A2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n483_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n553_), .A2(new_n515_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(G232gat), .A2(G233gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT34), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n575_), .A2(KEYINPUT35), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n575_), .A2(KEYINPUT35), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n572_), .A2(new_n573_), .A3(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n572_), .A2(new_n573_), .ZN(new_n580_));
  AOI22_X1  g379(.A1(new_n579_), .A2(KEYINPUT70), .B1(new_n580_), .B2(new_n576_), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n579_), .A2(KEYINPUT70), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  XOR2_X1   g382(.A(G190gat), .B(G218gat), .Z(new_n584_));
  XNOR2_X1  g383(.A(G134gat), .B(G162gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT36), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n586_), .A2(new_n587_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n583_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n581_), .A2(new_n582_), .A3(new_n587_), .A4(new_n586_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT71), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT37), .ZN(new_n594_));
  NOR3_X1   g393(.A1(new_n592_), .A2(new_n593_), .A3(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n593_), .A2(new_n594_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(KEYINPUT71), .A2(KEYINPUT37), .ZN(new_n597_));
  AOI211_X1 g396(.A(new_n596_), .B(new_n597_), .C1(new_n590_), .C2(new_n591_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n595_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G231gat), .A2(G233gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n549_), .B(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(new_n516_), .ZN(new_n603_));
  XOR2_X1   g402(.A(G183gat), .B(G211gat), .Z(new_n604_));
  XNOR2_X1  g403(.A(G127gat), .B(G155gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n606_), .B(new_n607_), .Z(new_n608_));
  INV_X1    g407(.A(KEYINPUT17), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n608_), .A2(new_n511_), .A3(new_n609_), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n603_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n608_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n612_), .A2(KEYINPUT17), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n603_), .B1(new_n613_), .B2(new_n610_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n611_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n600_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n571_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n619_), .A2(new_n544_), .A3(new_n368_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT38), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n592_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n623_), .A2(new_n616_), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n571_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n368_), .ZN(new_n627_));
  OAI21_X1  g426(.A(G1gat), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n620_), .A2(new_n621_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n622_), .A2(new_n628_), .A3(new_n629_), .ZN(G1324gat));
  AOI21_X1  g429(.A(new_n545_), .B1(new_n625_), .B2(new_n438_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT39), .Z(new_n632_));
  NAND3_X1  g431(.A1(new_n619_), .A2(new_n545_), .A3(new_n438_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(KEYINPUT96), .B(KEYINPUT40), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(G1325gat));
  OAI21_X1  g435(.A(G15gat), .B1(new_n626_), .B2(new_n252_), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n637_), .A2(KEYINPUT41), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(KEYINPUT41), .ZN(new_n639_));
  OR3_X1    g438(.A1(new_n618_), .A2(G15gat), .A3(new_n252_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n638_), .A2(new_n639_), .A3(new_n640_), .ZN(G1326gat));
  INV_X1    g440(.A(G22gat), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n642_), .B1(new_n625_), .B2(new_n339_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT42), .Z(new_n644_));
  NAND2_X1  g443(.A1(new_n339_), .A2(new_n642_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT97), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n644_), .B1(new_n618_), .B2(new_n646_), .ZN(G1327gat));
  NOR2_X1   g446(.A1(new_n592_), .A2(new_n615_), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n444_), .A2(new_n570_), .A3(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(G29gat), .B1(new_n649_), .B2(new_n368_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT43), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n651_), .B1(new_n444_), .B2(new_n600_), .ZN(new_n652_));
  AOI211_X1 g451(.A(KEYINPUT43), .B(new_n599_), .C1(new_n440_), .C2(new_n443_), .ZN(new_n653_));
  OAI211_X1 g452(.A(new_n570_), .B(new_n616_), .C1(new_n652_), .C2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT44), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n656_), .A2(G29gat), .A3(new_n368_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT98), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n658_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n659_));
  NOR4_X1   g458(.A1(new_n252_), .A2(new_n339_), .A3(new_n368_), .A4(new_n438_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n627_), .A2(new_n339_), .A3(new_n442_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n411_), .B1(new_n363_), .B2(new_n367_), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n418_), .A2(new_n402_), .A3(new_n395_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n402_), .B1(new_n418_), .B2(new_n395_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n424_), .B1(new_n351_), .B2(new_n354_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n425_), .A2(new_n344_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n665_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n668_), .B1(new_n414_), .B2(new_n367_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n662_), .B1(new_n669_), .B2(new_n429_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n661_), .B1(new_n670_), .B2(new_n339_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n660_), .B1(new_n671_), .B2(new_n252_), .ZN(new_n672_));
  OAI21_X1  g471(.A(KEYINPUT43), .B1(new_n672_), .B2(new_n599_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n444_), .A2(new_n651_), .A3(new_n600_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n615_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n675_), .A2(KEYINPUT98), .A3(KEYINPUT44), .A4(new_n570_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n659_), .A2(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n650_), .B1(new_n657_), .B2(new_n677_), .ZN(G1328gat));
  INV_X1    g477(.A(KEYINPUT101), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT99), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n442_), .A2(G36gat), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n649_), .A2(new_n680_), .A3(new_n681_), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n444_), .A2(new_n570_), .A3(new_n648_), .A4(new_n681_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(KEYINPUT99), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n682_), .A2(KEYINPUT45), .A3(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT46), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(KEYINPUT100), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n685_), .A2(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(KEYINPUT45), .B1(new_n682_), .B2(new_n684_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n656_), .A2(new_n438_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n691_), .B1(new_n659_), .B2(new_n676_), .ZN(new_n692_));
  INV_X1    g491(.A(G36gat), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n679_), .B(new_n690_), .C1(new_n692_), .C2(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n442_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n693_), .B1(new_n677_), .B2(new_n695_), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n688_), .A2(new_n689_), .ZN(new_n697_));
  OAI21_X1  g496(.A(KEYINPUT101), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n686_), .A2(KEYINPUT100), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n694_), .A2(new_n698_), .A3(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n694_), .B2(new_n698_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n700_), .A2(new_n701_), .ZN(G1329gat));
  INV_X1    g501(.A(G43gat), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n252_), .A2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n677_), .A2(new_n656_), .A3(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n649_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n703_), .B1(new_n706_), .B2(new_n252_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n707_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g508(.A(G50gat), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n649_), .A2(new_n710_), .A3(new_n339_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT102), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n434_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n677_), .A2(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n712_), .B1(new_n714_), .B2(G50gat), .ZN(new_n715_));
  AOI211_X1 g514(.A(KEYINPUT102), .B(new_n710_), .C1(new_n677_), .C2(new_n713_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n711_), .B1(new_n715_), .B2(new_n716_), .ZN(G1331gat));
  NOR2_X1   g516(.A1(new_n535_), .A2(new_n568_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n444_), .A2(new_n624_), .A3(new_n718_), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n719_), .A2(new_n490_), .A3(new_n627_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n444_), .A2(new_n569_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n721_), .A2(KEYINPUT103), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n721_), .A2(KEYINPUT103), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n722_), .A2(new_n723_), .A3(new_n535_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(new_n617_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n627_), .B1(new_n725_), .B2(KEYINPUT104), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n726_), .B1(KEYINPUT104), .B2(new_n725_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n720_), .B1(new_n727_), .B2(new_n490_), .ZN(G1332gat));
  OAI21_X1  g527(.A(G64gat), .B1(new_n719_), .B2(new_n442_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT48), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n438_), .A2(new_n491_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n730_), .B1(new_n725_), .B2(new_n731_), .ZN(G1333gat));
  OAI21_X1  g531(.A(G71gat), .B1(new_n719_), .B2(new_n252_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT49), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n252_), .A2(G71gat), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n734_), .B1(new_n725_), .B2(new_n735_), .ZN(G1334gat));
  OAI21_X1  g535(.A(G78gat), .B1(new_n719_), .B2(new_n434_), .ZN(new_n737_));
  XOR2_X1   g536(.A(KEYINPUT105), .B(KEYINPUT50), .Z(new_n738_));
  XNOR2_X1  g537(.A(new_n737_), .B(new_n738_), .ZN(new_n739_));
  OR2_X1    g538(.A1(new_n434_), .A2(G78gat), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n739_), .B1(new_n725_), .B2(new_n740_), .ZN(G1335gat));
  NAND2_X1  g540(.A1(new_n724_), .A2(new_n648_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n341_), .B1(new_n742_), .B2(new_n627_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n675_), .A2(new_n718_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n368_), .A2(G85gat), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n745_), .B(KEYINPUT106), .Z(new_n746_));
  OAI21_X1  g545(.A(new_n743_), .B1(new_n744_), .B2(new_n746_), .ZN(new_n747_));
  XOR2_X1   g546(.A(new_n747_), .B(KEYINPUT107), .Z(G1336gat));
  NOR3_X1   g547(.A1(new_n744_), .A2(new_n399_), .A3(new_n442_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n742_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(new_n438_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n749_), .B1(new_n751_), .B2(new_n399_), .ZN(G1337gat));
  OAI21_X1  g551(.A(G99gat), .B1(new_n744_), .B2(new_n252_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT108), .ZN(new_n754_));
  OR2_X1    g553(.A1(new_n252_), .A2(new_n452_), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n753_), .B(new_n754_), .C1(new_n742_), .C2(new_n755_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g556(.A1(new_n750_), .A2(new_n469_), .A3(new_n339_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT52), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n675_), .A2(new_n339_), .A3(new_n718_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n760_), .B2(G106gat), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n760_), .A2(new_n759_), .A3(G106gat), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n758_), .B1(new_n761_), .B2(new_n763_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR4_X1   g564(.A1(new_n627_), .A2(new_n252_), .A3(new_n339_), .A4(new_n438_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT117), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n555_), .A2(new_n557_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n551_), .A2(new_n556_), .A3(new_n559_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n565_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n770_), .B1(new_n561_), .B2(new_n565_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n529_), .A2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT113), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT113), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n529_), .A2(new_n774_), .A3(new_n771_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n568_), .A2(new_n528_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n514_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT12), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n779_), .B1(new_n483_), .B2(new_n497_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n445_), .A2(KEYINPUT111), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n778_), .A2(new_n780_), .A3(new_n781_), .ZN(new_n782_));
  OAI22_X1  g581(.A1(new_n514_), .A2(new_n517_), .B1(KEYINPUT111), .B2(new_n445_), .ZN(new_n783_));
  OR2_X1    g582(.A1(new_n446_), .A2(KEYINPUT55), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n782_), .A2(new_n783_), .A3(new_n784_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n512_), .A2(KEYINPUT12), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n515_), .A2(new_n510_), .A3(new_n787_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n780_), .A2(new_n445_), .A3(new_n506_), .A4(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT68), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n778_), .A2(new_n509_), .A3(new_n445_), .A4(new_n780_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n786_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT110), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n785_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  AOI211_X1 g593(.A(KEYINPUT110), .B(new_n786_), .C1(new_n790_), .C2(new_n791_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n526_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(KEYINPUT112), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT56), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n777_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n796_), .A2(KEYINPUT112), .A3(KEYINPUT56), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n776_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT116), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT57), .ZN(new_n803_));
  NOR4_X1   g602(.A1(new_n801_), .A2(new_n802_), .A3(new_n803_), .A4(new_n623_), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n782_), .A2(new_n783_), .A3(new_n784_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n786_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n806_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n805_), .B1(new_n807_), .B2(KEYINPUT110), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n792_), .A2(new_n793_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n525_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT112), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n798_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n777_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n812_), .A2(new_n800_), .A3(new_n813_), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n773_), .A2(new_n775_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n623_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(KEYINPUT116), .B1(new_n816_), .B2(KEYINPUT57), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n804_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT114), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n819_), .B1(new_n796_), .B2(new_n798_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n808_), .A2(new_n809_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n821_), .A2(KEYINPUT114), .A3(KEYINPUT56), .A4(new_n526_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n796_), .A2(new_n798_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n820_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT58), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT115), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n771_), .A2(new_n528_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n824_), .A2(new_n826_), .A3(new_n827_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n828_), .A2(new_n600_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n824_), .A2(new_n827_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n830_), .A2(KEYINPUT115), .A3(new_n825_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n814_), .A2(new_n815_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(new_n592_), .ZN(new_n833_));
  AOI22_X1  g632(.A1(new_n829_), .A2(new_n831_), .B1(new_n833_), .B2(new_n803_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n615_), .B1(new_n818_), .B2(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n617_), .A2(new_n569_), .A3(new_n535_), .ZN(new_n836_));
  XOR2_X1   g635(.A(new_n836_), .B(KEYINPUT54), .Z(new_n837_));
  OAI21_X1  g636(.A(new_n767_), .B1(new_n835_), .B2(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(KEYINPUT118), .B1(new_n835_), .B2(new_n837_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT59), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n838_), .A2(new_n839_), .A3(new_n840_), .ZN(new_n841_));
  OAI221_X1 g640(.A(new_n767_), .B1(KEYINPUT118), .B2(KEYINPUT59), .C1(new_n835_), .C2(new_n837_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT119), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n841_), .A2(KEYINPUT119), .A3(new_n842_), .ZN(new_n846_));
  INV_X1    g645(.A(G113gat), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n569_), .A2(new_n847_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n845_), .A2(new_n846_), .A3(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n847_), .B1(new_n838_), .B2(new_n569_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n849_), .A2(new_n850_), .ZN(G1340gat));
  INV_X1    g650(.A(G120gat), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n852_), .B1(new_n535_), .B2(KEYINPUT60), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n853_), .A2(KEYINPUT120), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(KEYINPUT120), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n855_), .B1(KEYINPUT60), .B2(new_n852_), .ZN(new_n856_));
  OR3_X1    g655(.A1(new_n838_), .A2(new_n854_), .A3(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n535_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n858_), .B2(new_n852_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(KEYINPUT121), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT121), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n861_), .B(new_n857_), .C1(new_n858_), .C2(new_n852_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n862_), .ZN(G1341gat));
  NAND2_X1  g662(.A1(new_n615_), .A2(G127gat), .ZN(new_n864_));
  XOR2_X1   g663(.A(new_n864_), .B(KEYINPUT122), .Z(new_n865_));
  NAND3_X1  g664(.A1(new_n845_), .A2(new_n846_), .A3(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(G127gat), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n867_), .B1(new_n838_), .B2(new_n616_), .ZN(new_n868_));
  AND2_X1   g667(.A1(new_n866_), .A2(new_n868_), .ZN(G1342gat));
  INV_X1    g668(.A(G134gat), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n599_), .A2(new_n870_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n845_), .A2(new_n846_), .A3(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n870_), .B1(new_n838_), .B2(new_n592_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n872_), .A2(new_n873_), .ZN(G1343gat));
  OR2_X1    g673(.A1(new_n835_), .A2(new_n837_), .ZN(new_n875_));
  AND4_X1   g674(.A1(new_n368_), .A2(new_n252_), .A3(new_n339_), .A4(new_n442_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n568_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g679(.A1(new_n878_), .A2(new_n536_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g681(.A(KEYINPUT123), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n878_), .A2(new_n883_), .A3(new_n615_), .ZN(new_n884_));
  OAI21_X1  g683(.A(KEYINPUT123), .B1(new_n877_), .B2(new_n616_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(KEYINPUT61), .B(G155gat), .ZN(new_n886_));
  AND3_X1   g685(.A1(new_n884_), .A2(new_n885_), .A3(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n886_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n887_), .A2(new_n888_), .ZN(G1346gat));
  AND3_X1   g688(.A1(new_n878_), .A2(G162gat), .A3(new_n600_), .ZN(new_n890_));
  AOI21_X1  g689(.A(G162gat), .B1(new_n878_), .B2(new_n623_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n890_), .A2(new_n891_), .ZN(G1347gat));
  XOR2_X1   g691(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n835_), .A2(new_n837_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n441_), .ZN(new_n896_));
  NOR4_X1   g695(.A1(new_n895_), .A2(new_n569_), .A3(new_n442_), .A4(new_n896_), .ZN(new_n897_));
  OAI21_X1  g696(.A(G169gat), .B1(new_n897_), .B2(KEYINPUT124), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n875_), .A2(new_n438_), .A3(new_n441_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT124), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n899_), .A2(new_n900_), .A3(new_n569_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n894_), .B1(new_n898_), .B2(new_n901_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n900_), .B1(new_n899_), .B2(new_n569_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n897_), .A2(KEYINPUT124), .ZN(new_n904_));
  NAND4_X1  g703(.A1(new_n903_), .A2(new_n904_), .A3(G169gat), .A4(new_n893_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n897_), .A2(new_n377_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n902_), .A2(new_n905_), .A3(new_n906_), .ZN(G1348gat));
  NOR3_X1   g706(.A1(new_n895_), .A2(new_n442_), .A3(new_n896_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(new_n536_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT126), .ZN(new_n910_));
  AND3_X1   g709(.A1(new_n909_), .A2(new_n910_), .A3(new_n230_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n910_), .B1(new_n909_), .B2(new_n230_), .ZN(new_n912_));
  INV_X1    g711(.A(G176gat), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n909_), .A2(new_n913_), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n911_), .A2(new_n912_), .A3(new_n914_), .ZN(G1349gat));
  NOR2_X1   g714(.A1(new_n899_), .A2(new_n616_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n916_), .A2(G183gat), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n210_), .A2(new_n381_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n917_), .B1(new_n918_), .B2(new_n916_), .ZN(G1350gat));
  OAI21_X1  g718(.A(G190gat), .B1(new_n899_), .B2(new_n599_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n908_), .A2(new_n208_), .A3(new_n623_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n920_), .A2(new_n921_), .ZN(G1351gat));
  AND3_X1   g721(.A1(new_n252_), .A2(new_n627_), .A3(new_n339_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n875_), .A2(new_n438_), .A3(new_n923_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n924_), .A2(new_n569_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(new_n275_), .ZN(G1352gat));
  NOR2_X1   g725(.A1(new_n924_), .A2(new_n535_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(new_n277_), .ZN(G1353gat));
  NOR2_X1   g727(.A1(new_n895_), .A2(new_n442_), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n929_), .A2(new_n615_), .A3(new_n923_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n931_));
  AND2_X1   g730(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n932_));
  NOR3_X1   g731(.A1(new_n930_), .A2(new_n931_), .A3(new_n932_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n933_), .B1(new_n930_), .B2(new_n931_), .ZN(G1354gat));
  OAI21_X1  g733(.A(G218gat), .B1(new_n924_), .B2(new_n599_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT127), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n592_), .A2(G218gat), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n929_), .A2(new_n923_), .A3(new_n937_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n935_), .A2(new_n936_), .A3(new_n938_), .ZN(new_n939_));
  INV_X1    g738(.A(new_n939_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n936_), .B1(new_n935_), .B2(new_n938_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n940_), .A2(new_n941_), .ZN(G1355gat));
endmodule


