//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 0 1 0 1 0 0 0 1 1 1 1 1 0 1 1 1 1 0 0 1 1 1 0 1 1 0 1 0 0 0 1 0 0 0 1 1 1 0 1 1 1 0 0 1 1 0 0 1 0 0 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n670_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n841_, new_n842_, new_n843_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n850_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n880_, new_n881_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n889_,
    new_n890_, new_n892_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_;
  XOR2_X1   g000(.A(G71gat), .B(G99gat), .Z(new_n202_));
  NAND2_X1  g001(.A1(G227gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(G15gat), .B(G43gat), .Z(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XOR2_X1   g005(.A(KEYINPUT80), .B(G190gat), .Z(new_n207_));
  INV_X1    g006(.A(G183gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT23), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G169gat), .ZN(new_n213_));
  INV_X1    g012(.A(G176gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT22), .B(G169gat), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n215_), .B1(new_n216_), .B2(new_n214_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n212_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(G190gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n219_), .A2(KEYINPUT26), .ZN(new_n220_));
  XOR2_X1   g019(.A(KEYINPUT25), .B(G183gat), .Z(new_n221_));
  AOI211_X1 g020(.A(new_n220_), .B(new_n221_), .C1(KEYINPUT26), .C2(new_n207_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n215_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n213_), .A2(new_n214_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n223_), .A2(KEYINPUT24), .A3(new_n224_), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n211_), .B(new_n225_), .C1(KEYINPUT24), .C2(new_n224_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n218_), .B1(new_n222_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT30), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n227_), .B(new_n228_), .ZN(new_n229_));
  AND2_X1   g028(.A1(new_n229_), .A2(KEYINPUT81), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n229_), .A2(KEYINPUT81), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n206_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n232_), .B1(new_n230_), .B2(new_n206_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G127gat), .B(G134gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G113gat), .B(G120gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n237_));
  XOR2_X1   g036(.A(new_n236_), .B(new_n237_), .Z(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n233_), .A2(new_n239_), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n232_), .B(new_n238_), .C1(new_n230_), .C2(new_n206_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(G197gat), .ZN(new_n244_));
  AND2_X1   g043(.A1(new_n244_), .A2(G204gat), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n244_), .A2(G204gat), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT21), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G211gat), .B(G218gat), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT94), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n245_), .A2(new_n246_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(KEYINPUT93), .A2(KEYINPUT21), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n246_), .A2(KEYINPUT93), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n254_), .B(new_n248_), .C1(new_n247_), .C2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n251_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT95), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G228gat), .A2(G233gat), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n257_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT1), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G155gat), .A2(G162gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT84), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT84), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n264_), .A2(G155gat), .A3(G162gat), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n261_), .B1(new_n263_), .B2(new_n265_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(G155gat), .A2(G162gat), .ZN(new_n267_));
  OR3_X1    g066(.A1(new_n266_), .A2(KEYINPUT85), .A3(new_n267_), .ZN(new_n268_));
  AND2_X1   g067(.A1(new_n263_), .A2(new_n265_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(new_n261_), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT85), .B1(new_n266_), .B2(new_n267_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n268_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G141gat), .A2(G148gat), .ZN(new_n273_));
  XOR2_X1   g072(.A(new_n273_), .B(KEYINPUT83), .Z(new_n274_));
  NOR2_X1   g073(.A1(G141gat), .A2(G148gat), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n272_), .A2(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n269_), .A2(new_n267_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT89), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT2), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n279_), .B1(new_n273_), .B2(new_n280_), .ZN(new_n281_));
  NAND4_X1  g080(.A1(KEYINPUT89), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT87), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT3), .ZN(new_n284_));
  AOI211_X1 g083(.A(G141gat), .B(G148gat), .C1(new_n284_), .C2(KEYINPUT86), .ZN(new_n285_));
  OAI21_X1  g084(.A(KEYINPUT86), .B1(G141gat), .B2(G148gat), .ZN(new_n286_));
  AOI21_X1  g085(.A(KEYINPUT3), .B1(new_n286_), .B2(new_n283_), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n281_), .B(new_n282_), .C1(new_n285_), .C2(new_n287_), .ZN(new_n288_));
  XOR2_X1   g087(.A(KEYINPUT88), .B(KEYINPUT2), .Z(new_n289_));
  NOR2_X1   g088(.A1(new_n274_), .A2(new_n289_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n278_), .B1(new_n288_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n277_), .A2(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n260_), .B1(KEYINPUT29), .B2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G78gat), .B(G106gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n294_), .ZN(new_n296_));
  AND2_X1   g095(.A1(new_n277_), .A2(new_n291_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT29), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n296_), .B1(new_n299_), .B2(new_n260_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n297_), .A2(new_n298_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G22gat), .B(G50gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  XOR2_X1   g102(.A(KEYINPUT91), .B(KEYINPUT92), .Z(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n292_), .A2(KEYINPUT29), .ZN(new_n306_));
  INV_X1    g105(.A(new_n302_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  AND3_X1   g107(.A1(new_n303_), .A2(new_n305_), .A3(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n305_), .B1(new_n303_), .B2(new_n308_), .ZN(new_n310_));
  OAI211_X1 g109(.A(new_n295_), .B(new_n300_), .C1(new_n309_), .C2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n310_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n295_), .A2(new_n300_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n303_), .A2(new_n305_), .A3(new_n308_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n312_), .A2(new_n313_), .A3(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n259_), .A2(new_n258_), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n316_), .B(new_n317_), .Z(new_n318_));
  NAND3_X1  g117(.A1(new_n311_), .A2(new_n315_), .A3(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n318_), .B1(new_n311_), .B2(new_n315_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n243_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n321_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n323_), .A2(new_n242_), .A3(new_n319_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT20), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n217_), .B(KEYINPUT96), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n211_), .B1(G183gat), .B2(G190gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n221_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT26), .B(G190gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n328_), .B1(new_n226_), .B2(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n325_), .B1(new_n333_), .B2(new_n257_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n334_), .B1(new_n227_), .B2(new_n257_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G226gat), .A2(G233gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT19), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n335_), .A2(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n325_), .B1(new_n257_), .B2(new_n227_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n337_), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n339_), .B(new_n340_), .C1(new_n257_), .C2(new_n333_), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n338_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G8gat), .B(G36gat), .ZN(new_n343_));
  INV_X1    g142(.A(G92gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT18), .B(G64gat), .ZN(new_n346_));
  XOR2_X1   g145(.A(new_n345_), .B(new_n346_), .Z(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n342_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n338_), .A2(new_n341_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(new_n347_), .ZN(new_n351_));
  AOI21_X1  g150(.A(KEYINPUT27), .B1(new_n349_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT98), .ZN(new_n353_));
  OR2_X1    g152(.A1(new_n333_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n257_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n333_), .A2(new_n353_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n354_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n340_), .B1(new_n357_), .B2(new_n339_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n335_), .A2(new_n337_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n347_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  AND2_X1   g159(.A1(new_n349_), .A2(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n352_), .B1(new_n361_), .B2(KEYINPUT27), .ZN(new_n362_));
  INV_X1    g161(.A(new_n236_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n292_), .A2(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n277_), .A2(new_n291_), .A3(new_n236_), .ZN(new_n365_));
  AND2_X1   g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G225gat), .A2(G233gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n364_), .A2(KEYINPUT4), .A3(new_n365_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n367_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT4), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n292_), .A2(new_n371_), .A3(new_n363_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n369_), .A2(new_n370_), .A3(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n368_), .A2(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G1gat), .B(G29gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(G85gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT0), .B(G57gat), .ZN(new_n377_));
  XOR2_X1   g176(.A(new_n376_), .B(new_n377_), .Z(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n374_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT99), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n368_), .A2(new_n373_), .A3(new_n378_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n380_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n368_), .A2(new_n373_), .A3(KEYINPUT99), .A4(new_n378_), .ZN(new_n384_));
  AND2_X1   g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  AOI22_X1  g185(.A1(new_n322_), .A2(new_n324_), .B1(new_n362_), .B2(new_n386_), .ZN(new_n387_));
  AND2_X1   g186(.A1(new_n348_), .A2(KEYINPUT32), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n388_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(KEYINPUT97), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n342_), .A2(new_n390_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n385_), .A2(KEYINPUT100), .A3(new_n389_), .A4(new_n391_), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n383_), .A2(new_n384_), .A3(new_n389_), .A4(new_n391_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT100), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n382_), .B(KEYINPUT33), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n366_), .A2(new_n370_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n369_), .A2(new_n367_), .A3(new_n372_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n397_), .A2(new_n398_), .A3(new_n379_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n396_), .A2(new_n349_), .A3(new_n351_), .A4(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n392_), .A2(new_n395_), .A3(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n323_), .A2(new_n319_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n324_), .A2(new_n322_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n387_), .B1(new_n403_), .B2(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G29gat), .B(G36gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G43gat), .B(G50gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(KEYINPUT15), .ZN(new_n410_));
  AND2_X1   g209(.A1(G99gat), .A2(G106gat), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT67), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n413_), .A2(KEYINPUT6), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT6), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n415_), .A2(KEYINPUT67), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n412_), .B1(new_n414_), .B2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n415_), .A2(KEYINPUT67), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n413_), .A2(KEYINPUT6), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(new_n419_), .A3(new_n411_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n417_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G85gat), .A2(G92gat), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(KEYINPUT65), .B1(new_n423_), .B2(KEYINPUT9), .ZN(new_n424_));
  NOR2_X1   g223(.A1(G85gat), .A2(G92gat), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT65), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT9), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n422_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n424_), .A2(new_n426_), .A3(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n431_), .B(KEYINPUT66), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n421_), .B1(new_n430_), .B2(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(KEYINPUT10), .B(G99gat), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(G106gat), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n435_), .A2(KEYINPUT64), .A3(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT64), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n438_), .B1(new_n434_), .B2(G106gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  OR2_X1    g239(.A1(new_n433_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT8), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n442_), .A2(KEYINPUT69), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT7), .ZN(new_n445_));
  INV_X1    g244(.A(G99gat), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n445_), .A2(new_n446_), .A3(new_n436_), .A4(KEYINPUT68), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT68), .ZN(new_n448_));
  OAI22_X1  g247(.A1(new_n448_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n423_), .B1(new_n421_), .B2(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n444_), .B1(new_n452_), .B2(new_n426_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n450_), .B1(new_n417_), .B2(new_n420_), .ZN(new_n454_));
  NOR4_X1   g253(.A1(new_n454_), .A2(new_n443_), .A3(new_n425_), .A4(new_n423_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n441_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n456_), .A2(KEYINPUT73), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT73), .ZN(new_n458_));
  AND3_X1   g257(.A1(new_n418_), .A2(new_n419_), .A3(new_n411_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n411_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  OAI211_X1 g260(.A(new_n426_), .B(new_n422_), .C1(new_n461_), .C2(new_n450_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(new_n443_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n452_), .A2(new_n444_), .A3(new_n426_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n458_), .B1(new_n465_), .B2(new_n441_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n410_), .B1(new_n457_), .B2(new_n466_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n433_), .A2(new_n440_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n468_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G232gat), .A2(G233gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n470_), .B(KEYINPUT34), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  XOR2_X1   g271(.A(KEYINPUT74), .B(KEYINPUT35), .Z(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  AOI22_X1  g273(.A1(new_n469_), .A2(new_n409_), .B1(new_n472_), .B2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n467_), .A2(new_n475_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n472_), .A2(new_n474_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G190gat), .B(G218gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G134gat), .B(G162gat), .ZN(new_n480_));
  XOR2_X1   g279(.A(new_n479_), .B(new_n480_), .Z(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  OR2_X1    g281(.A1(new_n482_), .A2(KEYINPUT36), .ZN(new_n483_));
  OR2_X1    g282(.A1(new_n478_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n482_), .A2(KEYINPUT36), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n478_), .A2(new_n483_), .A3(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n484_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT37), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT37), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n484_), .A2(new_n486_), .A3(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT77), .ZN(new_n493_));
  XNOR2_X1  g292(.A(KEYINPUT75), .B(G15gat), .ZN(new_n494_));
  INV_X1    g293(.A(G22gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(G1gat), .ZN(new_n497_));
  INV_X1    g296(.A(G8gat), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT14), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n496_), .A2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G1gat), .B(G8gat), .ZN(new_n501_));
  OR2_X1    g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n500_), .A2(new_n501_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(G231gat), .ZN(new_n505_));
  INV_X1    g304(.A(G233gat), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n504_), .B(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G57gat), .A2(G64gat), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(G57gat), .A2(G64gat), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT70), .ZN(new_n513_));
  NOR3_X1   g312(.A1(new_n511_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(G57gat), .ZN(new_n515_));
  INV_X1    g314(.A(G64gat), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(KEYINPUT70), .B1(new_n517_), .B2(new_n510_), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT11), .B1(new_n514_), .B2(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n513_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n517_), .A2(KEYINPUT70), .A3(new_n510_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT11), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n520_), .A2(new_n521_), .A3(new_n522_), .ZN(new_n523_));
  XOR2_X1   g322(.A(G71gat), .B(G78gat), .Z(new_n524_));
  NAND3_X1  g323(.A1(new_n519_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(KEYINPUT71), .B(KEYINPUT72), .ZN(new_n526_));
  INV_X1    g325(.A(new_n524_), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n527_), .B(KEYINPUT11), .C1(new_n518_), .C2(new_n514_), .ZN(new_n528_));
  AND3_X1   g327(.A1(new_n525_), .A2(new_n526_), .A3(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n526_), .B1(new_n525_), .B2(new_n528_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n509_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n525_), .A2(new_n528_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n526_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n525_), .A2(new_n526_), .A3(new_n528_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n504_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n538_), .A2(new_n508_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n504_), .A2(new_n507_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n537_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n493_), .B1(new_n532_), .B2(new_n541_), .ZN(new_n542_));
  XOR2_X1   g341(.A(KEYINPUT76), .B(KEYINPUT16), .Z(new_n543_));
  XNOR2_X1  g342(.A(G127gat), .B(G155gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G183gat), .B(G211gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NOR3_X1   g347(.A1(new_n542_), .A2(KEYINPUT17), .A3(new_n548_), .ZN(new_n549_));
  OR2_X1    g348(.A1(new_n542_), .A2(new_n548_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT17), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n532_), .A2(new_n541_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n551_), .B1(new_n552_), .B2(new_n548_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n549_), .B1(new_n550_), .B2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n492_), .A2(new_n555_), .ZN(new_n556_));
  OAI211_X1 g355(.A(KEYINPUT12), .B(new_n531_), .C1(new_n457_), .C2(new_n466_), .ZN(new_n557_));
  AOI21_X1  g356(.A(KEYINPUT12), .B1(new_n531_), .B2(new_n456_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n531_), .A2(new_n456_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(G230gat), .A2(G233gat), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n557_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n531_), .B(new_n469_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n562_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(KEYINPUT5), .B(G176gat), .Z(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(G204gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G120gat), .B(G148gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  AND2_X1   g367(.A1(new_n564_), .A2(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n564_), .A2(new_n568_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT13), .ZN(new_n571_));
  OR3_X1    g370(.A1(new_n569_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n571_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n538_), .A2(new_n409_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G229gat), .A2(G233gat), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n504_), .A2(new_n410_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n575_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n504_), .B(new_n409_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n578_), .B1(new_n579_), .B2(new_n576_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(KEYINPUT78), .B(G113gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(G141gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G169gat), .B(G197gat), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n582_), .B(new_n583_), .Z(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n580_), .A2(new_n585_), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n578_), .B(new_n584_), .C1(new_n579_), .C2(new_n576_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT79), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n574_), .A2(new_n590_), .ZN(new_n591_));
  AND3_X1   g390(.A1(new_n406_), .A2(new_n556_), .A3(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n592_), .A2(new_n497_), .A3(new_n385_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT38), .ZN(new_n594_));
  INV_X1    g393(.A(new_n588_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n574_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT101), .ZN(new_n597_));
  AND3_X1   g396(.A1(new_n484_), .A2(new_n486_), .A3(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n597_), .B1(new_n484_), .B2(new_n486_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n406_), .A2(new_n554_), .A3(new_n596_), .A4(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(G1gat), .B1(new_n601_), .B2(new_n386_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n594_), .A2(new_n602_), .ZN(G1324gat));
  OAI21_X1  g402(.A(G8gat), .B1(new_n601_), .B2(new_n362_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT102), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  OAI211_X1 g405(.A(KEYINPUT102), .B(G8gat), .C1(new_n601_), .C2(new_n362_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n606_), .A2(KEYINPUT39), .A3(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n362_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n592_), .A2(new_n498_), .A3(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT39), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n604_), .A2(new_n605_), .A3(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n608_), .A2(new_n610_), .A3(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT40), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(G1325gat));
  INV_X1    g414(.A(G15gat), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n592_), .A2(new_n616_), .A3(new_n243_), .ZN(new_n617_));
  OAI21_X1  g416(.A(G15gat), .B1(new_n601_), .B2(new_n242_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT41), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n618_), .A2(new_n619_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n617_), .B1(new_n620_), .B2(new_n621_), .ZN(G1326gat));
  INV_X1    g421(.A(new_n402_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n592_), .A2(new_n495_), .A3(new_n623_), .ZN(new_n624_));
  OAI21_X1  g423(.A(G22gat), .B1(new_n601_), .B2(new_n402_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n625_), .A2(KEYINPUT42), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n625_), .A2(KEYINPUT42), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n624_), .B1(new_n626_), .B2(new_n627_), .ZN(G1327gat));
  NOR3_X1   g427(.A1(new_n574_), .A2(new_n554_), .A3(new_n595_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT43), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n630_), .B1(new_n406_), .B2(new_n492_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n404_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n632_));
  NOR4_X1   g431(.A1(new_n632_), .A2(KEYINPUT43), .A3(new_n387_), .A4(new_n491_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n629_), .B1(new_n631_), .B2(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(KEYINPUT103), .A2(KEYINPUT44), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  OAI221_X1 g435(.A(new_n629_), .B1(KEYINPUT103), .B2(KEYINPUT44), .C1(new_n631_), .C2(new_n633_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n636_), .A2(new_n637_), .A3(new_n385_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT104), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n636_), .A2(new_n637_), .A3(KEYINPUT104), .A4(new_n385_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n640_), .A2(G29gat), .A3(new_n641_), .ZN(new_n642_));
  NOR3_X1   g441(.A1(new_n632_), .A2(new_n600_), .A3(new_n387_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n643_), .A2(new_n555_), .A3(new_n591_), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n386_), .A2(G29gat), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n642_), .B1(new_n644_), .B2(new_n645_), .ZN(G1328gat));
  NAND3_X1  g445(.A1(new_n636_), .A2(new_n637_), .A3(new_n609_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(G36gat), .ZN(new_n648_));
  INV_X1    g447(.A(new_n644_), .ZN(new_n649_));
  INV_X1    g448(.A(G36gat), .ZN(new_n650_));
  XOR2_X1   g449(.A(new_n362_), .B(KEYINPUT105), .Z(new_n651_));
  NAND3_X1  g450(.A1(new_n649_), .A2(new_n650_), .A3(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(KEYINPUT45), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT45), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n649_), .A2(new_n654_), .A3(new_n650_), .A4(new_n651_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n653_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n648_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT46), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n648_), .A2(KEYINPUT46), .A3(new_n656_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(G1329gat));
  NAND4_X1  g460(.A1(new_n636_), .A2(new_n637_), .A3(G43gat), .A4(new_n243_), .ZN(new_n662_));
  INV_X1    g461(.A(G43gat), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n663_), .B1(new_n644_), .B2(new_n242_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(KEYINPUT106), .B(KEYINPUT47), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n665_), .B(new_n666_), .ZN(G1330gat));
  NAND3_X1  g466(.A1(new_n636_), .A2(new_n637_), .A3(new_n623_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(G50gat), .ZN(new_n669_));
  OR2_X1    g468(.A1(new_n644_), .A2(G50gat), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n669_), .B1(new_n402_), .B2(new_n670_), .ZN(G1331gat));
  INV_X1    g470(.A(new_n600_), .ZN(new_n672_));
  NOR3_X1   g471(.A1(new_n632_), .A2(new_n672_), .A3(new_n387_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n588_), .B(KEYINPUT79), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n555_), .A2(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n673_), .A2(new_n574_), .A3(new_n675_), .ZN(new_n676_));
  NOR3_X1   g475(.A1(new_n676_), .A2(new_n515_), .A3(new_n386_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n574_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n678_), .A2(new_n588_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n406_), .A2(new_n556_), .A3(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(G57gat), .B1(new_n681_), .B2(new_n385_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n677_), .A2(new_n682_), .ZN(G1332gat));
  NAND3_X1  g482(.A1(new_n681_), .A2(new_n516_), .A3(new_n651_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n676_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(new_n651_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(KEYINPUT107), .B(KEYINPUT48), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n686_), .A2(G64gat), .A3(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(new_n686_), .B2(G64gat), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n684_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(KEYINPUT108), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT108), .ZN(new_n692_));
  OAI211_X1 g491(.A(new_n692_), .B(new_n684_), .C1(new_n688_), .C2(new_n689_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(G1333gat));
  NAND2_X1  g493(.A1(new_n685_), .A2(new_n243_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(G71gat), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(KEYINPUT109), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT109), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n695_), .A2(new_n698_), .A3(G71gat), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n697_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT49), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  OR3_X1    g501(.A1(new_n680_), .A2(G71gat), .A3(new_n242_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n697_), .A2(KEYINPUT49), .A3(new_n699_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n702_), .A2(new_n703_), .A3(new_n704_), .ZN(G1334gat));
  OR3_X1    g504(.A1(new_n680_), .A2(G78gat), .A3(new_n402_), .ZN(new_n706_));
  OAI21_X1  g505(.A(G78gat), .B1(new_n676_), .B2(new_n402_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n707_), .A2(KEYINPUT50), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n707_), .A2(KEYINPUT50), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n706_), .B1(new_n708_), .B2(new_n709_), .ZN(G1335gat));
  NOR3_X1   g509(.A1(new_n678_), .A2(new_n554_), .A3(new_n588_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n643_), .A2(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(G85gat), .B1(new_n712_), .B2(new_n385_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT110), .ZN(new_n714_));
  OR2_X1    g513(.A1(new_n631_), .A2(new_n633_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(new_n711_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n385_), .A2(G85gat), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT111), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n714_), .B1(new_n717_), .B2(new_n719_), .ZN(G1336gat));
  AOI21_X1  g519(.A(G92gat), .B1(new_n712_), .B2(new_n609_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n716_), .A2(new_n344_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n722_), .B2(new_n651_), .ZN(G1337gat));
  OAI211_X1 g522(.A(new_n243_), .B(new_n711_), .C1(new_n631_), .C2(new_n633_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n242_), .A2(new_n434_), .ZN(new_n725_));
  AOI22_X1  g524(.A1(new_n724_), .A2(G99gat), .B1(new_n712_), .B2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT112), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n727_), .A2(KEYINPUT51), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n726_), .A2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(KEYINPUT51), .ZN(new_n730_));
  XOR2_X1   g529(.A(new_n729_), .B(new_n730_), .Z(G1338gat));
  XNOR2_X1  g530(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT52), .ZN(new_n733_));
  OAI211_X1 g532(.A(new_n623_), .B(new_n711_), .C1(new_n631_), .C2(new_n633_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n734_), .B2(G106gat), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n734_), .A2(new_n733_), .A3(G106gat), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n712_), .A2(new_n436_), .A3(new_n623_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n732_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n737_), .ZN(new_n741_));
  OAI211_X1 g540(.A(new_n739_), .B(new_n732_), .C1(new_n741_), .C2(new_n735_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n740_), .A2(new_n743_), .ZN(G1339gat));
  INV_X1    g543(.A(KEYINPUT121), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT12), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n746_), .B1(new_n537_), .B2(new_n469_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n537_), .A2(new_n469_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n456_), .A2(KEYINPUT73), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n469_), .A2(new_n458_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n537_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n749_), .B1(KEYINPUT12), .B2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT115), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n753_), .A2(new_n754_), .A3(KEYINPUT55), .A4(new_n561_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT55), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n562_), .A2(new_n756_), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n557_), .A2(new_n560_), .A3(KEYINPUT55), .A4(new_n561_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT115), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n557_), .A2(new_n560_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n760_), .A2(G230gat), .A3(G233gat), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n755_), .A2(new_n757_), .A3(new_n759_), .A4(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(new_n568_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT56), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT118), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n762_), .A2(KEYINPUT56), .A3(new_n568_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n765_), .A2(new_n766_), .A3(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n576_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n575_), .A2(new_n769_), .A3(new_n577_), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n770_), .B(new_n585_), .C1(new_n579_), .C2(new_n769_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n771_), .A2(KEYINPUT116), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n771_), .A2(KEYINPUT116), .ZN(new_n773_));
  INV_X1    g572(.A(new_n587_), .ZN(new_n774_));
  NOR3_X1   g573(.A1(new_n772_), .A2(new_n773_), .A3(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(KEYINPUT56), .B1(new_n762_), .B2(new_n568_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n570_), .B1(new_n776_), .B2(KEYINPUT118), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n768_), .A2(new_n775_), .A3(new_n777_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(KEYINPUT119), .A2(KEYINPUT58), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n779_), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n768_), .A2(new_n777_), .A3(new_n781_), .A4(new_n775_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n780_), .A2(new_n492_), .A3(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT120), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT57), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n775_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT117), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n775_), .B(KEYINPUT117), .C1(new_n569_), .C2(new_n570_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n588_), .B1(new_n564_), .B2(new_n568_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n792_), .B1(new_n765_), .B2(new_n767_), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n600_), .B(new_n786_), .C1(new_n791_), .C2(new_n793_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n784_), .A2(new_n785_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n600_), .B(new_n795_), .C1(new_n791_), .C2(new_n793_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n783_), .A2(new_n797_), .A3(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n555_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT114), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n801_), .B1(new_n590_), .B2(new_n554_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n802_), .B1(new_n488_), .B2(new_n490_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT54), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n590_), .A2(new_n801_), .A3(new_n554_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n803_), .A2(new_n804_), .A3(new_n678_), .A4(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(KEYINPUT114), .B1(new_n555_), .B2(new_n674_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n491_), .A2(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n805_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n809_));
  OAI21_X1  g608(.A(KEYINPUT54), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  AND2_X1   g609(.A1(new_n806_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n386_), .B1(new_n800_), .B2(new_n812_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n609_), .A2(new_n322_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n745_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n811_), .B1(new_n799_), .B2(new_n555_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n814_), .ZN(new_n817_));
  NOR4_X1   g616(.A1(new_n816_), .A2(KEYINPUT121), .A3(new_n386_), .A4(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n588_), .B1(new_n815_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(G113gat), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT59), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n821_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n822_));
  NOR4_X1   g621(.A1(new_n816_), .A2(KEYINPUT59), .A3(new_n386_), .A4(new_n817_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(KEYINPUT122), .B(G113gat), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n590_), .A2(new_n825_), .ZN(new_n826_));
  AOI22_X1  g625(.A1(new_n819_), .A2(new_n820_), .B1(new_n824_), .B2(new_n826_), .ZN(G1340gat));
  NOR3_X1   g626(.A1(new_n822_), .A2(new_n823_), .A3(new_n678_), .ZN(new_n828_));
  INV_X1    g627(.A(G120gat), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n829_), .B1(new_n678_), .B2(KEYINPUT60), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n830_), .B1(new_n815_), .B2(new_n818_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n829_), .A2(KEYINPUT60), .ZN(new_n832_));
  OAI22_X1  g631(.A1(new_n828_), .A2(new_n829_), .B1(new_n831_), .B2(new_n832_), .ZN(G1341gat));
  INV_X1    g632(.A(KEYINPUT123), .ZN(new_n834_));
  OAI21_X1  g633(.A(G127gat), .B1(new_n555_), .B2(new_n834_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n834_), .A2(G127gat), .ZN(new_n836_));
  NOR3_X1   g635(.A1(new_n822_), .A2(new_n823_), .A3(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n554_), .B1(new_n815_), .B2(new_n818_), .ZN(new_n838_));
  INV_X1    g637(.A(G127gat), .ZN(new_n839_));
  AOI22_X1  g638(.A1(new_n835_), .A2(new_n837_), .B1(new_n838_), .B2(new_n839_), .ZN(G1342gat));
  INV_X1    g639(.A(G134gat), .ZN(new_n841_));
  NOR3_X1   g640(.A1(new_n822_), .A2(new_n823_), .A3(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n672_), .B1(new_n815_), .B2(new_n818_), .ZN(new_n843_));
  AOI22_X1  g642(.A1(new_n492_), .A2(new_n842_), .B1(new_n843_), .B2(new_n841_), .ZN(G1343gat));
  AOI21_X1  g643(.A(new_n324_), .B1(new_n800_), .B2(new_n812_), .ZN(new_n845_));
  OR2_X1    g644(.A1(new_n651_), .A2(new_n386_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n845_), .A2(new_n588_), .A3(new_n847_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n848_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g648(.A1(new_n845_), .A2(new_n574_), .A3(new_n847_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g650(.A1(new_n845_), .A2(new_n554_), .A3(new_n847_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(KEYINPUT61), .B(G155gat), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n852_), .B(new_n853_), .ZN(G1346gat));
  NAND4_X1  g653(.A1(new_n845_), .A2(G162gat), .A3(new_n492_), .A4(new_n847_), .ZN(new_n855_));
  NOR4_X1   g654(.A1(new_n816_), .A2(new_n600_), .A3(new_n324_), .A4(new_n846_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n855_), .B1(new_n856_), .B2(G162gat), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(KEYINPUT124), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT124), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n855_), .B(new_n859_), .C1(new_n856_), .C2(G162gat), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n858_), .A2(new_n860_), .ZN(G1347gat));
  INV_X1    g660(.A(KEYINPUT62), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n800_), .A2(new_n812_), .ZN(new_n863_));
  AND2_X1   g662(.A1(new_n651_), .A2(new_n386_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n865_), .A2(new_n242_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n863_), .A2(new_n402_), .A3(new_n866_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n867_), .A2(new_n595_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n862_), .B1(new_n868_), .B2(new_n213_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n216_), .ZN(new_n870_));
  OAI211_X1 g669(.A(KEYINPUT62), .B(G169gat), .C1(new_n867_), .C2(new_n595_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n869_), .A2(new_n870_), .A3(new_n871_), .ZN(G1348gat));
  INV_X1    g671(.A(new_n867_), .ZN(new_n873_));
  AOI21_X1  g672(.A(G176gat), .B1(new_n873_), .B2(new_n574_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n863_), .A2(KEYINPUT125), .A3(new_n402_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT125), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n876_), .B1(new_n816_), .B2(new_n623_), .ZN(new_n877_));
  AND4_X1   g676(.A1(new_n574_), .A2(new_n875_), .A3(new_n866_), .A4(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n874_), .B1(new_n878_), .B2(G176gat), .ZN(G1349gat));
  NOR3_X1   g678(.A1(new_n867_), .A2(new_n555_), .A3(new_n329_), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n875_), .A2(new_n877_), .A3(new_n554_), .A4(new_n866_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n880_), .B1(new_n208_), .B2(new_n881_), .ZN(G1350gat));
  NAND3_X1  g681(.A1(new_n873_), .A2(new_n672_), .A3(new_n330_), .ZN(new_n883_));
  NAND4_X1  g682(.A1(new_n863_), .A2(new_n402_), .A3(new_n492_), .A4(new_n866_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT126), .ZN(new_n885_));
  AND3_X1   g684(.A1(new_n884_), .A2(new_n885_), .A3(G190gat), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n885_), .B1(new_n884_), .B2(G190gat), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n883_), .B1(new_n886_), .B2(new_n887_), .ZN(G1351gat));
  NOR3_X1   g687(.A1(new_n816_), .A2(new_n324_), .A3(new_n865_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(new_n588_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n574_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g692(.A1(new_n889_), .A2(new_n554_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(KEYINPUT63), .B(G211gat), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n896_), .B1(new_n894_), .B2(new_n897_), .ZN(G1354gat));
  AOI21_X1  g697(.A(G218gat), .B1(new_n889_), .B2(new_n672_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n492_), .A2(G218gat), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(KEYINPUT127), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n899_), .B1(new_n889_), .B2(new_n901_), .ZN(G1355gat));
endmodule


