//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 1 1 0 1 0 1 1 0 0 1 1 1 1 1 0 1 1 1 1 0 1 0 0 1 0 0 1 0 1 1 1 1 1 0 1 1 0 1 1 1 0 1 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n777_, new_n778_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n829_, new_n830_, new_n831_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n929_, new_n930_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n948_, new_n950_, new_n952_, new_n953_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n970_,
    new_n972_, new_n973_, new_n974_, new_n975_, new_n976_, new_n977_,
    new_n978_, new_n980_, new_n981_, new_n982_, new_n984_, new_n985_,
    new_n986_, new_n987_, new_n988_, new_n990_, new_n991_, new_n992_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1000_, new_n1001_, new_n1003_, new_n1004_, new_n1005_, new_n1006_;
  INV_X1    g000(.A(G8gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT76), .B(G1gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT14), .B1(new_n203_), .B2(new_n202_), .ZN(new_n204_));
  INV_X1    g003(.A(G1gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G15gat), .B(G22gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n205_), .B1(new_n204_), .B2(new_n206_), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n202_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n204_), .A2(new_n206_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G1gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(G8gat), .A3(new_n207_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n210_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G231gat), .A2(G233gat), .ZN(new_n215_));
  XOR2_X1   g014(.A(new_n215_), .B(KEYINPUT77), .Z(new_n216_));
  AND2_X1   g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n214_), .A2(new_n216_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(G71gat), .B(G78gat), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G57gat), .A2(G64gat), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(G57gat), .A2(G64gat), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT68), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G57gat), .ZN(new_n225_));
  INV_X1    g024(.A(G64gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT68), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(new_n228_), .A3(new_n221_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n224_), .A2(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n220_), .B1(new_n230_), .B2(KEYINPUT11), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT11), .ZN(new_n232_));
  AOI211_X1 g031(.A(new_n232_), .B(new_n219_), .C1(new_n224_), .C2(new_n229_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n230_), .A2(KEYINPUT11), .ZN(new_n234_));
  OR3_X1    g033(.A1(new_n231_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  OR3_X1    g034(.A1(new_n217_), .A2(new_n218_), .A3(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT78), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G127gat), .B(G155gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT16), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(G183gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(G211gat), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n237_), .B1(new_n241_), .B2(KEYINPUT17), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n235_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n243_));
  AND3_X1   g042(.A1(new_n236_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n242_), .B1(new_n236_), .B2(new_n243_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n241_), .A2(KEYINPUT17), .ZN(new_n246_));
  NOR3_X1   g045(.A1(new_n244_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G232gat), .A2(G233gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT70), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT34), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT35), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT73), .ZN(new_n253_));
  INV_X1    g052(.A(G85gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT65), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT65), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(G85gat), .ZN(new_n257_));
  INV_X1    g056(.A(G92gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT66), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT66), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(G92gat), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n255_), .A2(new_n257_), .A3(new_n259_), .A4(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT9), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(G85gat), .A2(G92gat), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n264_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G99gat), .A2(G106gat), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT67), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n271_), .A2(KEYINPUT6), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT6), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n273_), .A2(KEYINPUT67), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n270_), .B1(new_n272_), .B2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n273_), .A2(KEYINPUT67), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n271_), .A2(KEYINPUT6), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n276_), .A2(new_n277_), .A3(new_n269_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n275_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(KEYINPUT10), .B(G99gat), .Z(new_n281_));
  INV_X1    g080(.A(G106gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n268_), .A2(new_n280_), .A3(new_n283_), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT7), .ZN(new_n286_));
  INV_X1    g085(.A(G99gat), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n286_), .A2(new_n287_), .A3(new_n282_), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n275_), .A2(new_n278_), .A3(new_n285_), .A4(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT8), .ZN(new_n290_));
  XOR2_X1   g089(.A(G85gat), .B(G92gat), .Z(new_n291_));
  AND3_X1   g090(.A1(new_n289_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n290_), .B1(new_n289_), .B2(new_n291_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n284_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  AND2_X1   g093(.A1(G29gat), .A2(G36gat), .ZN(new_n295_));
  NOR2_X1   g094(.A1(G29gat), .A2(G36gat), .ZN(new_n296_));
  OAI21_X1  g095(.A(KEYINPUT71), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(G29gat), .ZN(new_n298_));
  INV_X1    g097(.A(G36gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT71), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G29gat), .A2(G36gat), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n300_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G43gat), .B(G50gat), .ZN(new_n304_));
  AND3_X1   g103(.A1(new_n297_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n304_), .B1(new_n297_), .B2(new_n303_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT72), .B(KEYINPUT15), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n297_), .A2(new_n303_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n304_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n297_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n308_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n309_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n294_), .A2(new_n317_), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n284_), .B(new_n314_), .C1(new_n292_), .C2(new_n293_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n253_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n253_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n250_), .A2(new_n251_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n252_), .B1(new_n320_), .B2(new_n323_), .ZN(new_n324_));
  AND3_X1   g123(.A1(new_n276_), .A2(new_n277_), .A3(new_n269_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n269_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n288_), .A2(new_n285_), .ZN(new_n327_));
  NOR3_X1   g126(.A1(new_n325_), .A2(new_n326_), .A3(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n291_), .ZN(new_n329_));
  OAI21_X1  g128(.A(KEYINPUT8), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n289_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n265_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n279_), .B1(new_n332_), .B2(new_n267_), .ZN(new_n333_));
  AOI22_X1  g132(.A1(new_n330_), .A2(new_n331_), .B1(new_n333_), .B2(new_n283_), .ZN(new_n334_));
  NOR3_X1   g133(.A1(new_n305_), .A2(new_n306_), .A3(new_n315_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n308_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n319_), .B1(new_n334_), .B2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(KEYINPUT73), .ZN(new_n339_));
  INV_X1    g138(.A(new_n252_), .ZN(new_n340_));
  AOI22_X1  g139(.A1(new_n319_), .A2(new_n253_), .B1(new_n251_), .B2(new_n250_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n339_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n324_), .A2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G190gat), .B(G218gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(G134gat), .ZN(new_n345_));
  INV_X1    g144(.A(G162gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT36), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n343_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT37), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT36), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n324_), .A2(new_n342_), .A3(new_n351_), .A4(new_n347_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n349_), .A2(new_n350_), .A3(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT75), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT74), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n355_), .B1(new_n343_), .B2(new_n348_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n348_), .ZN(new_n357_));
  AOI211_X1 g156(.A(KEYINPUT74), .B(new_n357_), .C1(new_n324_), .C2(new_n342_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n352_), .ZN(new_n359_));
  NOR3_X1   g158(.A1(new_n356_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n354_), .B1(new_n360_), .B2(new_n350_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n349_), .A2(KEYINPUT74), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n343_), .A2(new_n355_), .A3(new_n348_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n362_), .A2(new_n352_), .A3(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n364_), .A2(KEYINPUT75), .A3(KEYINPUT37), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n247_), .B1(new_n361_), .B2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT79), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT93), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT22), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(G169gat), .ZN(new_n370_));
  INV_X1    g169(.A(G169gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(KEYINPUT22), .ZN(new_n372_));
  INV_X1    g171(.A(G176gat), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n370_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n371_), .A2(new_n373_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n368_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n375_), .A2(KEYINPUT93), .ZN(new_n378_));
  OAI21_X1  g177(.A(KEYINPUT94), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT94), .ZN(new_n380_));
  INV_X1    g179(.A(new_n378_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(KEYINPUT22), .B(G169gat), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n375_), .B1(new_n382_), .B2(new_n373_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n380_), .B(new_n381_), .C1(new_n383_), .C2(new_n368_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G183gat), .A2(G190gat), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT82), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(KEYINPUT82), .A2(G183gat), .A3(G190gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n389_), .A2(KEYINPUT23), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT23), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n391_), .B1(G183gat), .B2(G190gat), .ZN(new_n392_));
  OAI22_X1  g191(.A1(new_n390_), .A2(new_n392_), .B1(G183gat), .B2(G190gat), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n379_), .A2(new_n384_), .A3(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT95), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(G204gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(G197gat), .ZN(new_n398_));
  INV_X1    g197(.A(G197gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(G204gat), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n398_), .A2(new_n400_), .A3(KEYINPUT90), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT21), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G211gat), .B(G218gat), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT21), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n398_), .A2(new_n400_), .A3(KEYINPUT90), .A4(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n402_), .A2(new_n403_), .A3(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT91), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n399_), .A2(G204gat), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n397_), .A2(G197gat), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n407_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n398_), .A2(new_n400_), .A3(KEYINPUT91), .ZN(new_n411_));
  XOR2_X1   g210(.A(G211gat), .B(G218gat), .Z(new_n412_));
  NAND4_X1  g211(.A1(new_n410_), .A2(KEYINPUT21), .A3(new_n411_), .A4(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n406_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  XOR2_X1   g214(.A(KEYINPUT25), .B(G183gat), .Z(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT26), .B(G190gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NOR3_X1   g218(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n420_), .B1(new_n376_), .B2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n419_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n385_), .A2(new_n391_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n425_), .B1(new_n389_), .B2(new_n391_), .ZN(new_n426_));
  OR2_X1    g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n379_), .A2(new_n384_), .A3(new_n393_), .A4(KEYINPUT95), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n396_), .A2(new_n415_), .A3(new_n427_), .A4(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G226gat), .A2(G233gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n430_), .B(KEYINPUT19), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT20), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n369_), .B1(KEYINPUT83), .B2(G169gat), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n369_), .A2(KEYINPUT83), .A3(G169gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n373_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(G183gat), .A2(G190gat), .ZN(new_n437_));
  OAI221_X1 g236(.A(new_n376_), .B1(new_n434_), .B2(new_n436_), .C1(new_n426_), .C2(new_n437_), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n419_), .B(new_n423_), .C1(new_n390_), .C2(new_n392_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n433_), .B1(new_n440_), .B2(new_n414_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n429_), .A2(new_n432_), .A3(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT20), .B1(new_n440_), .B2(new_n414_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n396_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n443_), .B1(new_n444_), .B2(new_n414_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n442_), .B1(new_n445_), .B2(new_n432_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G8gat), .B(G36gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(KEYINPUT18), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(G64gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(new_n258_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n446_), .A2(new_n451_), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n450_), .B(new_n442_), .C1(new_n445_), .C2(new_n432_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT96), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G1gat), .B(G29gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(new_n254_), .ZN(new_n457_));
  OR2_X1    g256(.A1(new_n457_), .A2(KEYINPUT0), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(KEYINPUT0), .ZN(new_n459_));
  AND3_X1   g258(.A1(new_n458_), .A2(G57gat), .A3(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(G57gat), .B1(new_n458_), .B2(new_n459_), .ZN(new_n461_));
  OR2_X1    g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(G120gat), .ZN(new_n463_));
  OR2_X1    g262(.A1(G127gat), .A2(G134gat), .ZN(new_n464_));
  INV_X1    g263(.A(G113gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G127gat), .A2(G134gat), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n464_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n465_), .B1(new_n464_), .B2(new_n466_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n463_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n469_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n471_), .A2(G120gat), .A3(new_n467_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G155gat), .A2(G162gat), .ZN(new_n474_));
  OR2_X1    g273(.A1(new_n474_), .A2(KEYINPUT1), .ZN(new_n475_));
  OR2_X1    g274(.A1(G155gat), .A2(G162gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(KEYINPUT1), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n475_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(G141gat), .A2(G148gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(KEYINPUT85), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G141gat), .A2(G148gat), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n478_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n476_), .A2(new_n474_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT2), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n481_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n481_), .A2(new_n485_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT86), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n481_), .A2(KEYINPUT86), .A3(new_n485_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n486_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n479_), .B(KEYINPUT3), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n484_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n473_), .B1(new_n483_), .B2(new_n493_), .ZN(new_n494_));
  AND3_X1   g293(.A1(new_n481_), .A2(KEYINPUT86), .A3(new_n485_), .ZN(new_n495_));
  AOI21_X1  g294(.A(KEYINPUT86), .B1(new_n481_), .B2(new_n485_), .ZN(new_n496_));
  OAI22_X1  g295(.A1(new_n495_), .A2(new_n496_), .B1(new_n485_), .B2(new_n481_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT3), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n479_), .B(new_n498_), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n476_), .B(new_n474_), .C1(new_n497_), .C2(new_n499_), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n500_), .A2(new_n472_), .A3(new_n470_), .A4(new_n482_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n494_), .A2(new_n501_), .A3(KEYINPUT4), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G225gat), .A2(G233gat), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT4), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n473_), .B(new_n504_), .C1(new_n483_), .C2(new_n493_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n502_), .A2(new_n503_), .A3(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n503_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n494_), .A2(new_n501_), .A3(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n462_), .A2(new_n506_), .A3(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT97), .ZN(new_n510_));
  OR2_X1    g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n509_), .A2(new_n510_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n502_), .A2(new_n507_), .A3(new_n505_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n460_), .A2(new_n461_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n494_), .A2(new_n501_), .A3(new_n503_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n513_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT33), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT33), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n513_), .A2(new_n518_), .A3(new_n514_), .A4(new_n515_), .ZN(new_n519_));
  AOI22_X1  g318(.A1(new_n511_), .A2(new_n512_), .B1(new_n517_), .B2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT96), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n452_), .A2(new_n521_), .A3(new_n453_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n455_), .A2(new_n520_), .A3(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n445_), .A2(new_n432_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT98), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n414_), .A2(KEYINPUT92), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT92), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n406_), .A2(new_n413_), .A3(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n530_), .A2(new_n427_), .A3(new_n394_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(new_n441_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(new_n431_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n445_), .A2(KEYINPUT98), .A3(new_n432_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n526_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n535_));
  AND2_X1   g334(.A1(new_n450_), .A2(KEYINPUT32), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT99), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n516_), .A2(new_n538_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n513_), .A2(KEYINPUT99), .A3(new_n514_), .A4(new_n515_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n513_), .A2(new_n515_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n542_), .A2(KEYINPUT100), .A3(new_n462_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(KEYINPUT100), .B1(new_n542_), .B2(new_n462_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n541_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  OR2_X1    g345(.A1(new_n446_), .A2(new_n536_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n537_), .A2(new_n546_), .A3(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n523_), .A2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n550_));
  XNOR2_X1  g349(.A(KEYINPUT88), .B(G22gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT29), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n500_), .A2(new_n553_), .A3(new_n482_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G78gat), .B(G106gat), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n555_), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n500_), .A2(new_n553_), .A3(new_n482_), .A4(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n552_), .B1(new_n556_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n556_), .A2(new_n552_), .A3(new_n558_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(KEYINPUT89), .A2(G233gat), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(KEYINPUT89), .A2(G233gat), .ZN(new_n565_));
  OAI21_X1  g364(.A(G228gat), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  AND3_X1   g365(.A1(new_n406_), .A2(new_n528_), .A3(new_n413_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n528_), .B1(new_n406_), .B2(new_n413_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(KEYINPUT29), .B1(new_n483_), .B2(new_n493_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n566_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n553_), .B1(new_n500_), .B2(new_n482_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n566_), .ZN(new_n573_));
  NOR3_X1   g372(.A1(new_n572_), .A2(new_n415_), .A3(new_n573_), .ZN(new_n574_));
  NOR3_X1   g373(.A1(new_n571_), .A2(new_n574_), .A3(G50gat), .ZN(new_n575_));
  INV_X1    g374(.A(G50gat), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n573_), .B1(new_n530_), .B2(new_n572_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n570_), .A2(new_n414_), .A3(new_n566_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n576_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n562_), .B1(new_n575_), .B2(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(G50gat), .B1(new_n571_), .B2(new_n574_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n577_), .A2(new_n576_), .A3(new_n578_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n581_), .A2(new_n582_), .A3(new_n560_), .A4(new_n561_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n580_), .A2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G15gat), .B(G71gat), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n585_), .B1(new_n470_), .B2(new_n472_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n470_), .A2(new_n472_), .A3(new_n585_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G227gat), .A2(G233gat), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n589_), .B(KEYINPUT30), .Z(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n587_), .A2(new_n588_), .A3(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n588_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n590_), .B1(new_n593_), .B2(new_n586_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(KEYINPUT84), .B(G43gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT31), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(G99gat), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT31), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n596_), .B(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(new_n287_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n440_), .A2(new_n598_), .A3(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n598_), .A2(new_n601_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n603_), .A2(new_n439_), .A3(new_n438_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n595_), .A2(new_n605_), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n602_), .A2(new_n592_), .A3(new_n594_), .A4(new_n604_), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n584_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n542_), .A2(new_n462_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT100), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  AOI22_X1  g411(.A1(new_n612_), .A2(new_n543_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n580_), .A2(new_n608_), .A3(new_n583_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n608_), .B1(new_n580_), .B2(new_n583_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n613_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n453_), .A2(KEYINPUT27), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n618_), .B1(new_n535_), .B2(new_n451_), .ZN(new_n619_));
  AOI21_X1  g418(.A(KEYINPUT27), .B1(new_n452_), .B2(new_n453_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  AOI22_X1  g420(.A1(new_n549_), .A2(new_n609_), .B1(new_n617_), .B2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(G230gat), .A2(G233gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT64), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n294_), .A2(new_n235_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n330_), .A2(new_n331_), .ZN(new_n627_));
  NOR3_X1   g426(.A1(new_n231_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n627_), .A2(new_n628_), .A3(new_n284_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n626_), .A2(KEYINPUT12), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT12), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n294_), .A2(new_n631_), .A3(new_n235_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n625_), .B1(new_n630_), .B2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n626_), .A2(new_n629_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n633_), .B1(new_n625_), .B2(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(G120gat), .B(G148gat), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT5), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(G176gat), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(G204gat), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n635_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n630_), .A2(new_n632_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(new_n624_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n634_), .A2(new_n625_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n643_), .A2(new_n644_), .A3(new_n639_), .ZN(new_n645_));
  XOR2_X1   g444(.A(KEYINPUT69), .B(KEYINPUT13), .Z(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n641_), .A2(new_n645_), .A3(new_n647_), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n643_), .A2(new_n644_), .A3(new_n639_), .ZN(new_n649_));
  OAI22_X1  g448(.A1(new_n640_), .A2(new_n649_), .B1(KEYINPUT69), .B2(KEYINPUT13), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n648_), .A2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(G229gat), .A2(G233gat), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n210_), .A2(new_n307_), .A3(new_n213_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n307_), .B1(new_n210_), .B2(new_n213_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n653_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(KEYINPUT80), .ZN(new_n658_));
  INV_X1    g457(.A(new_n214_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(new_n317_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n214_), .A2(new_n314_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n660_), .A2(new_n652_), .A3(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n654_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT80), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n663_), .A2(new_n664_), .A3(new_n653_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n658_), .A2(new_n662_), .A3(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(G113gat), .B(G141gat), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT81), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(new_n371_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(new_n399_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n666_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n670_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n658_), .A2(new_n665_), .A3(new_n662_), .A4(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n671_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n651_), .A2(new_n674_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n622_), .A2(new_n675_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n367_), .A2(new_n676_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n613_), .B(KEYINPUT101), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n677_), .A2(new_n203_), .A3(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT103), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT38), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n680_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n683_), .B1(KEYINPUT103), .B2(KEYINPUT38), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n349_), .A2(new_n352_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n686_), .A2(new_n247_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n676_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT102), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n688_), .B(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(G1gat), .B1(new_n690_), .B2(new_n613_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n680_), .A2(new_n681_), .A3(new_n682_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n684_), .A2(new_n691_), .A3(new_n692_), .ZN(G1324gat));
  OAI21_X1  g492(.A(G8gat), .B1(new_n688_), .B2(new_n621_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT39), .ZN(new_n695_));
  INV_X1    g494(.A(new_n621_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n677_), .A2(new_n202_), .A3(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT40), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n698_), .B(new_n699_), .ZN(G1325gat));
  INV_X1    g499(.A(G15gat), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n677_), .A2(new_n701_), .A3(new_n608_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n608_), .ZN(new_n703_));
  OAI21_X1  g502(.A(G15gat), .B1(new_n690_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT41), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n704_), .A2(new_n705_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n702_), .B1(new_n706_), .B2(new_n707_), .ZN(G1326gat));
  INV_X1    g507(.A(G22gat), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n677_), .A2(new_n709_), .A3(new_n584_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n584_), .ZN(new_n711_));
  OR2_X1    g510(.A1(new_n690_), .A2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT42), .ZN(new_n713_));
  AND3_X1   g512(.A1(new_n712_), .A2(new_n713_), .A3(G22gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n712_), .B2(G22gat), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n710_), .B1(new_n714_), .B2(new_n715_), .ZN(G1327gat));
  NAND2_X1  g515(.A1(new_n686_), .A2(new_n247_), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT106), .Z(new_n718_));
  NAND2_X1  g517(.A1(new_n676_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n720_), .A2(new_n298_), .A3(new_n546_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n675_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT44), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(KEYINPUT105), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n722_), .A2(new_n247_), .A3(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n609_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n727_), .B1(new_n523_), .B2(new_n548_), .ZN(new_n728_));
  NOR3_X1   g527(.A1(new_n616_), .A2(new_n620_), .A3(new_n619_), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n361_), .B(new_n365_), .C1(new_n728_), .C2(new_n729_), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n730_), .A2(KEYINPUT104), .A3(KEYINPUT43), .ZN(new_n731_));
  AOI21_X1  g530(.A(KEYINPUT43), .B1(new_n730_), .B2(KEYINPUT104), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n726_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n723_), .A2(KEYINPUT105), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n734_), .ZN(new_n736_));
  OAI211_X1 g535(.A(new_n736_), .B(new_n726_), .C1(new_n731_), .C2(new_n732_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n678_), .B1(new_n735_), .B2(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n721_), .B1(new_n738_), .B2(new_n298_), .ZN(G1328gat));
  INV_X1    g538(.A(KEYINPUT46), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n676_), .A2(new_n299_), .A3(new_n696_), .A4(new_n718_), .ZN(new_n741_));
  OR2_X1    g540(.A1(new_n741_), .A2(KEYINPUT107), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(KEYINPUT107), .ZN(new_n743_));
  AOI21_X1  g542(.A(KEYINPUT45), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n742_), .A2(KEYINPUT45), .A3(new_n743_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n735_), .A2(new_n737_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n299_), .B1(new_n748_), .B2(new_n696_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n740_), .B1(new_n747_), .B2(new_n749_), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n742_), .A2(KEYINPUT45), .A3(new_n743_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n751_), .A2(new_n744_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n621_), .B1(new_n735_), .B2(new_n737_), .ZN(new_n753_));
  OAI211_X1 g552(.A(new_n752_), .B(KEYINPUT46), .C1(new_n299_), .C2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n750_), .A2(new_n754_), .ZN(G1329gat));
  INV_X1    g554(.A(KEYINPUT47), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n356_), .A2(new_n358_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n350_), .B1(new_n757_), .B2(new_n352_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n354_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n365_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(KEYINPUT104), .B1(new_n622_), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT43), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n730_), .A2(KEYINPUT104), .A3(KEYINPUT43), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n736_), .B1(new_n765_), .B2(new_n726_), .ZN(new_n766_));
  AOI211_X1 g565(.A(new_n734_), .B(new_n725_), .C1(new_n763_), .C2(new_n764_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n608_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(G43gat), .ZN(new_n769_));
  INV_X1    g568(.A(G43gat), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n720_), .A2(new_n770_), .A3(new_n608_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n756_), .B1(new_n769_), .B2(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n703_), .B1(new_n735_), .B2(new_n737_), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n756_), .B(new_n771_), .C1(new_n773_), .C2(new_n770_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n772_), .A2(new_n775_), .ZN(G1330gat));
  NAND3_X1  g575(.A1(new_n720_), .A2(new_n576_), .A3(new_n584_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n711_), .B1(new_n735_), .B2(new_n737_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n777_), .B1(new_n778_), .B2(new_n576_), .ZN(G1331gat));
  INV_X1    g578(.A(new_n651_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n674_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n782_), .A2(new_n622_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n687_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT108), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT108), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n783_), .A2(new_n786_), .A3(new_n687_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n785_), .A2(new_n787_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(KEYINPUT109), .B(G57gat), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n788_), .A2(new_n546_), .A3(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n367_), .A2(new_n783_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n225_), .B1(new_n791_), .B2(new_n678_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT110), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n793_), .B(new_n794_), .ZN(G1332gat));
  NAND4_X1  g594(.A1(new_n367_), .A2(new_n226_), .A3(new_n696_), .A4(new_n783_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n785_), .A2(new_n696_), .A3(new_n787_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(G64gat), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT111), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT111), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n797_), .A2(new_n800_), .A3(G64gat), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n799_), .A2(KEYINPUT48), .A3(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(KEYINPUT48), .B1(new_n799_), .B2(new_n801_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n796_), .B1(new_n802_), .B2(new_n803_), .ZN(G1333gat));
  OR3_X1    g603(.A1(new_n791_), .A2(G71gat), .A3(new_n703_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n788_), .A2(new_n608_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(G71gat), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n807_), .A2(KEYINPUT49), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n807_), .A2(KEYINPUT49), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n805_), .B1(new_n808_), .B2(new_n809_), .ZN(G1334gat));
  OR3_X1    g609(.A1(new_n791_), .A2(G78gat), .A3(new_n711_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n788_), .A2(new_n584_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT50), .ZN(new_n813_));
  AND3_X1   g612(.A1(new_n812_), .A2(new_n813_), .A3(G78gat), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n813_), .B1(new_n812_), .B2(G78gat), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n811_), .B1(new_n814_), .B2(new_n815_), .ZN(G1335gat));
  INV_X1    g615(.A(KEYINPUT112), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n765_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n247_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n782_), .A2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n763_), .A2(KEYINPUT112), .A3(new_n764_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n818_), .A2(new_n820_), .A3(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n546_), .A2(new_n255_), .A3(new_n257_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n783_), .A2(new_n718_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(G85gat), .B1(new_n826_), .B2(new_n679_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n824_), .A2(new_n827_), .ZN(G1336gat));
  NAND3_X1  g627(.A1(new_n696_), .A2(new_n259_), .A3(new_n261_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n822_), .A2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(G92gat), .B1(new_n826_), .B2(new_n696_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n830_), .A2(new_n831_), .ZN(G1337gat));
  OAI21_X1  g631(.A(G99gat), .B1(new_n822_), .B2(new_n703_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n826_), .A2(new_n281_), .A3(new_n608_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT51), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT51), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n833_), .A2(new_n837_), .A3(new_n834_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n838_), .ZN(G1338gat));
  NAND3_X1  g638(.A1(new_n826_), .A2(new_n282_), .A3(new_n584_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n765_), .A2(new_n584_), .A3(new_n820_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT52), .ZN(new_n842_));
  AND3_X1   g641(.A1(new_n841_), .A2(new_n842_), .A3(G106gat), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n842_), .B1(new_n841_), .B2(G106gat), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n840_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(KEYINPUT53), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n847_), .B(new_n840_), .C1(new_n843_), .C2(new_n844_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n848_), .ZN(G1339gat));
  OAI21_X1  g648(.A(new_n685_), .B1(KEYINPUT117), .B2(KEYINPUT57), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n674_), .A2(new_n645_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT114), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT55), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n643_), .A2(new_n853_), .A3(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n630_), .A2(new_n625_), .A3(new_n632_), .ZN(new_n856_));
  OAI21_X1  g655(.A(KEYINPUT55), .B1(new_n633_), .B2(KEYINPUT114), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n855_), .A2(new_n856_), .A3(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n639_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT56), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n858_), .A2(KEYINPUT56), .A3(new_n859_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n852_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n640_), .A2(new_n649_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n660_), .A2(new_n653_), .A3(new_n661_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n663_), .A2(new_n652_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n866_), .A2(new_n867_), .A3(new_n670_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n673_), .A2(new_n868_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n865_), .A2(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n851_), .B1(new_n864_), .B2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT117), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT57), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n872_), .B1(KEYINPUT115), .B2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n871_), .A2(new_n875_), .ZN(new_n876_));
  AND3_X1   g675(.A1(new_n364_), .A2(KEYINPUT75), .A3(KEYINPUT37), .ZN(new_n877_));
  AOI22_X1  g676(.A1(new_n364_), .A2(KEYINPUT37), .B1(KEYINPUT75), .B2(new_n353_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT116), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n880_), .B1(new_n869_), .B2(new_n649_), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n645_), .A2(new_n673_), .A3(KEYINPUT116), .A4(new_n868_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  AND3_X1   g682(.A1(new_n858_), .A2(KEYINPUT56), .A3(new_n859_), .ZN(new_n884_));
  AOI21_X1  g683(.A(KEYINPUT56), .B1(new_n858_), .B2(new_n859_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n883_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT58), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n883_), .B(KEYINPUT58), .C1(new_n884_), .C2(new_n885_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n879_), .A2(new_n888_), .A3(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n852_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n891_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n870_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n894_), .A2(new_n874_), .A3(new_n851_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n876_), .A2(new_n890_), .A3(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n247_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n674_), .B1(new_n648_), .B2(new_n650_), .ZN(new_n898_));
  OAI211_X1 g697(.A(new_n898_), .B(new_n819_), .C1(new_n877_), .C2(new_n878_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(KEYINPUT113), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT113), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n366_), .A2(new_n901_), .A3(new_n898_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n900_), .A2(new_n902_), .A3(KEYINPUT54), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT54), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n899_), .A2(KEYINPUT113), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n901_), .B1(new_n366_), .B2(new_n898_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n904_), .B1(new_n905_), .B2(new_n906_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n897_), .A2(new_n903_), .A3(new_n907_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n696_), .A2(new_n678_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(new_n614_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(KEYINPUT118), .ZN(new_n911_));
  AND2_X1   g710(.A1(new_n908_), .A2(new_n911_), .ZN(new_n912_));
  AOI21_X1  g711(.A(G113gat), .B1(new_n912_), .B2(new_n674_), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT59), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n908_), .A2(new_n914_), .A3(new_n911_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n914_), .B1(new_n908_), .B2(new_n911_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n916_), .A2(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n674_), .A2(G113gat), .ZN(new_n919_));
  XOR2_X1   g718(.A(new_n919_), .B(KEYINPUT119), .Z(new_n920_));
  AOI21_X1  g719(.A(new_n913_), .B1(new_n918_), .B2(new_n920_), .ZN(G1340gat));
  XNOR2_X1  g720(.A(KEYINPUT120), .B(G120gat), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n780_), .A2(new_n922_), .ZN(new_n923_));
  INV_X1    g722(.A(KEYINPUT60), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(new_n924_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n651_), .B1(new_n912_), .B2(new_n925_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n912_), .A2(new_n924_), .A3(new_n925_), .ZN(new_n927_));
  AOI22_X1  g726(.A1(new_n918_), .A2(new_n926_), .B1(new_n927_), .B2(new_n922_), .ZN(G1341gat));
  AOI21_X1  g727(.A(G127gat), .B1(new_n912_), .B2(new_n819_), .ZN(new_n929_));
  AND2_X1   g728(.A1(new_n819_), .A2(G127gat), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n929_), .B1(new_n918_), .B2(new_n930_), .ZN(G1342gat));
  NAND2_X1  g730(.A1(new_n908_), .A2(new_n911_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(KEYINPUT59), .ZN(new_n933_));
  INV_X1    g732(.A(G134gat), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n760_), .A2(new_n934_), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n933_), .A2(new_n915_), .A3(new_n935_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n907_), .A2(new_n903_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n874_), .B1(new_n894_), .B2(new_n851_), .ZN(new_n938_));
  AOI211_X1 g737(.A(new_n875_), .B(new_n850_), .C1(new_n892_), .C2(new_n893_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n938_), .A2(new_n939_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n819_), .B1(new_n940_), .B2(new_n890_), .ZN(new_n941_));
  OAI211_X1 g740(.A(new_n686_), .B(new_n911_), .C1(new_n937_), .C2(new_n941_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n942_), .A2(new_n934_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n943_), .A2(KEYINPUT121), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT121), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n942_), .A2(new_n945_), .A3(new_n934_), .ZN(new_n946_));
  AND3_X1   g745(.A1(new_n936_), .A2(new_n944_), .A3(new_n946_), .ZN(G1343gat));
  NAND4_X1  g746(.A1(new_n908_), .A2(new_n674_), .A3(new_n615_), .A4(new_n909_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(G141gat), .ZN(G1344gat));
  NAND4_X1  g748(.A1(new_n908_), .A2(new_n780_), .A3(new_n615_), .A4(new_n909_), .ZN(new_n950_));
  XNOR2_X1  g749(.A(new_n950_), .B(G148gat), .ZN(G1345gat));
  NAND4_X1  g750(.A1(new_n908_), .A2(new_n615_), .A3(new_n819_), .A4(new_n909_), .ZN(new_n952_));
  XNOR2_X1  g751(.A(KEYINPUT61), .B(G155gat), .ZN(new_n953_));
  XNOR2_X1  g752(.A(new_n952_), .B(new_n953_), .ZN(G1346gat));
  AND2_X1   g753(.A1(new_n908_), .A2(new_n615_), .ZN(new_n955_));
  AND2_X1   g754(.A1(new_n955_), .A2(new_n909_), .ZN(new_n956_));
  NOR2_X1   g755(.A1(new_n760_), .A2(new_n346_), .ZN(new_n957_));
  NAND3_X1  g756(.A1(new_n955_), .A2(new_n686_), .A3(new_n909_), .ZN(new_n958_));
  AOI22_X1  g757(.A1(new_n956_), .A2(new_n957_), .B1(new_n958_), .B2(new_n346_), .ZN(G1347gat));
  NOR3_X1   g758(.A1(new_n679_), .A2(new_n703_), .A3(new_n621_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n960_), .A2(new_n674_), .ZN(new_n961_));
  XOR2_X1   g760(.A(new_n961_), .B(KEYINPUT122), .Z(new_n962_));
  NAND3_X1  g761(.A1(new_n908_), .A2(new_n711_), .A3(new_n962_), .ZN(new_n963_));
  INV_X1    g762(.A(KEYINPUT62), .ZN(new_n964_));
  AND3_X1   g763(.A1(new_n963_), .A2(new_n964_), .A3(G169gat), .ZN(new_n965_));
  AOI21_X1  g764(.A(new_n964_), .B1(new_n963_), .B2(G169gat), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n908_), .A2(new_n711_), .ZN(new_n967_));
  NAND3_X1  g766(.A1(new_n960_), .A2(new_n674_), .A3(new_n382_), .ZN(new_n968_));
  OAI22_X1  g767(.A1(new_n965_), .A2(new_n966_), .B1(new_n967_), .B2(new_n968_), .ZN(G1348gat));
  NAND4_X1  g768(.A1(new_n908_), .A2(new_n780_), .A3(new_n711_), .A4(new_n960_), .ZN(new_n970_));
  XNOR2_X1  g769(.A(new_n970_), .B(G176gat), .ZN(G1349gat));
  AND3_X1   g770(.A1(new_n908_), .A2(new_n711_), .A3(new_n960_), .ZN(new_n972_));
  INV_X1    g771(.A(KEYINPUT123), .ZN(new_n973_));
  NAND4_X1  g772(.A1(new_n972_), .A2(new_n973_), .A3(new_n416_), .A4(new_n819_), .ZN(new_n974_));
  NAND4_X1  g773(.A1(new_n908_), .A2(new_n711_), .A3(new_n819_), .A4(new_n960_), .ZN(new_n975_));
  INV_X1    g774(.A(G183gat), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n975_), .A2(new_n976_), .ZN(new_n977_));
  OAI21_X1  g776(.A(KEYINPUT123), .B1(new_n975_), .B2(new_n417_), .ZN(new_n978_));
  AND3_X1   g777(.A1(new_n974_), .A2(new_n977_), .A3(new_n978_), .ZN(G1350gat));
  NAND2_X1  g778(.A1(new_n972_), .A2(new_n879_), .ZN(new_n980_));
  NAND2_X1  g779(.A1(new_n980_), .A2(G190gat), .ZN(new_n981_));
  NAND3_X1  g780(.A1(new_n972_), .A2(new_n418_), .A3(new_n686_), .ZN(new_n982_));
  NAND2_X1  g781(.A1(new_n981_), .A2(new_n982_), .ZN(G1351gat));
  NAND2_X1  g782(.A1(new_n613_), .A2(new_n615_), .ZN(new_n984_));
  XOR2_X1   g783(.A(new_n984_), .B(KEYINPUT124), .Z(new_n985_));
  NAND3_X1  g784(.A1(new_n908_), .A2(new_n696_), .A3(new_n985_), .ZN(new_n986_));
  NOR2_X1   g785(.A1(new_n986_), .A2(new_n781_), .ZN(new_n987_));
  XNOR2_X1  g786(.A(KEYINPUT125), .B(G197gat), .ZN(new_n988_));
  XNOR2_X1  g787(.A(new_n987_), .B(new_n988_), .ZN(G1352gat));
  NOR2_X1   g788(.A1(new_n986_), .A2(new_n651_), .ZN(new_n990_));
  XNOR2_X1  g789(.A(KEYINPUT126), .B(G204gat), .ZN(new_n991_));
  INV_X1    g790(.A(new_n991_), .ZN(new_n992_));
  XNOR2_X1  g791(.A(new_n990_), .B(new_n992_), .ZN(G1353gat));
  NAND4_X1  g792(.A1(new_n908_), .A2(new_n696_), .A3(new_n819_), .A4(new_n985_), .ZN(new_n994_));
  NOR2_X1   g793(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n995_));
  AND2_X1   g794(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n996_));
  NOR3_X1   g795(.A1(new_n994_), .A2(new_n995_), .A3(new_n996_), .ZN(new_n997_));
  NAND2_X1  g796(.A1(new_n994_), .A2(new_n995_), .ZN(new_n998_));
  INV_X1    g797(.A(KEYINPUT127), .ZN(new_n999_));
  NAND2_X1  g798(.A1(new_n998_), .A2(new_n999_), .ZN(new_n1000_));
  NAND3_X1  g799(.A1(new_n994_), .A2(KEYINPUT127), .A3(new_n995_), .ZN(new_n1001_));
  AOI21_X1  g800(.A(new_n997_), .B1(new_n1000_), .B2(new_n1001_), .ZN(G1354gat));
  INV_X1    g801(.A(G218gat), .ZN(new_n1003_));
  NOR3_X1   g802(.A1(new_n986_), .A2(new_n1003_), .A3(new_n760_), .ZN(new_n1004_));
  INV_X1    g803(.A(new_n986_), .ZN(new_n1005_));
  NAND2_X1  g804(.A1(new_n1005_), .A2(new_n686_), .ZN(new_n1006_));
  AOI21_X1  g805(.A(new_n1004_), .B1(new_n1003_), .B2(new_n1006_), .ZN(G1355gat));
endmodule


