//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 0 0 1 1 0 1 1 1 0 1 1 0 0 1 1 1 0 1 0 1 1 1 1 0 0 0 0 0 1 0 1 1 0 1 0 0 1 0 0 0 1 1 0 0 0 1 1 1 0 0 0 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n651_, new_n652_, new_n653_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n763_, new_n764_,
    new_n765_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n774_, new_n775_, new_n776_, new_n778_, new_n779_,
    new_n780_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n887_,
    new_n888_, new_n889_, new_n891_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n914_, new_n915_, new_n917_,
    new_n918_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n937_, new_n938_,
    new_n939_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n952_,
    new_n953_, new_n954_;
  NOR2_X1   g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  AND2_X1   g001(.A1(G183gat), .A2(G190gat), .ZN(new_n203_));
  AOI21_X1  g002(.A(new_n202_), .B1(new_n203_), .B2(KEYINPUT23), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G183gat), .A2(G190gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n204_), .A2(new_n207_), .ZN(new_n208_));
  OR2_X1    g007(.A1(KEYINPUT79), .A2(G176gat), .ZN(new_n209_));
  INV_X1    g008(.A(G169gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT22), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT22), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(G169gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(KEYINPUT79), .A2(G176gat), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n209_), .A2(new_n211_), .A3(new_n213_), .A4(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n208_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT25), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT77), .B1(new_n218_), .B2(G183gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT77), .ZN(new_n220_));
  INV_X1    g019(.A(G183gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n220_), .A2(new_n221_), .A3(KEYINPUT25), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n218_), .A2(G183gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n219_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT26), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT78), .ZN(new_n226_));
  INV_X1    g025(.A(G190gat), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n225_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(KEYINPUT78), .A2(KEYINPUT26), .A3(G190gat), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n224_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n205_), .A2(KEYINPUT23), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n206_), .A2(G183gat), .A3(G190gat), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT24), .ZN(new_n233_));
  NOR2_X1   g032(.A1(G169gat), .A2(G176gat), .ZN(new_n234_));
  AOI22_X1  g033(.A1(new_n231_), .A2(new_n232_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n234_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n236_), .A2(KEYINPUT24), .A3(new_n216_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n235_), .A2(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n217_), .B1(new_n230_), .B2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT30), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G227gat), .A2(G233gat), .ZN(new_n241_));
  INV_X1    g040(.A(G15gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(G71gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(G99gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n240_), .B(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(G134gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(G127gat), .ZN(new_n248_));
  INV_X1    g047(.A(G127gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(G134gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(G120gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(G113gat), .ZN(new_n253_));
  INV_X1    g052(.A(G113gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(G120gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n251_), .A2(new_n256_), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n248_), .A2(new_n250_), .A3(new_n253_), .A4(new_n255_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n246_), .A2(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT80), .B(G43gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT31), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  OR2_X1    g063(.A1(new_n240_), .A2(new_n245_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n240_), .A2(new_n245_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n259_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  OR3_X1    g066(.A1(new_n261_), .A2(new_n264_), .A3(new_n267_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n264_), .B1(new_n261_), .B2(new_n267_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT91), .B(KEYINPUT27), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT86), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n221_), .A2(KEYINPUT25), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n227_), .A2(KEYINPUT26), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n225_), .A2(G190gat), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n274_), .A2(new_n223_), .A3(new_n275_), .A4(new_n276_), .ZN(new_n277_));
  AND2_X1   g076(.A1(new_n235_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT84), .ZN(new_n279_));
  AND3_X1   g078(.A1(new_n216_), .A2(new_n279_), .A3(KEYINPUT24), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n279_), .B1(new_n216_), .B2(KEYINPUT24), .ZN(new_n281_));
  OR3_X1    g080(.A1(new_n280_), .A2(new_n281_), .A3(new_n234_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT85), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n212_), .A2(G169gat), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n210_), .A2(KEYINPUT22), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n283_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  AND2_X1   g085(.A1(new_n209_), .A2(new_n214_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n211_), .A2(new_n213_), .A3(KEYINPUT85), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n286_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  AOI22_X1  g088(.A1(new_n204_), .A2(new_n207_), .B1(G169gat), .B2(G176gat), .ZN(new_n290_));
  AOI22_X1  g089(.A1(new_n278_), .A2(new_n282_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  XOR2_X1   g090(.A(G211gat), .B(G218gat), .Z(new_n292_));
  NOR2_X1   g091(.A1(G197gat), .A2(G204gat), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G197gat), .A2(G204gat), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n292_), .A2(KEYINPUT21), .A3(new_n294_), .A4(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n294_), .A2(KEYINPUT21), .A3(new_n295_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT21), .ZN(new_n298_));
  AND2_X1   g097(.A1(G197gat), .A2(G204gat), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n298_), .B1(new_n299_), .B2(new_n293_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G211gat), .B(G218gat), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n297_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  AND2_X1   g101(.A1(new_n296_), .A2(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n273_), .B1(new_n291_), .B2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT20), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n231_), .A2(new_n232_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n234_), .A2(new_n233_), .ZN(new_n307_));
  AND3_X1   g106(.A1(new_n237_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n228_), .A2(new_n229_), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n309_), .A2(new_n222_), .A3(new_n223_), .A4(new_n219_), .ZN(new_n310_));
  AOI22_X1  g109(.A1(new_n308_), .A2(new_n310_), .B1(new_n290_), .B2(new_n215_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n305_), .B1(new_n311_), .B2(new_n303_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n296_), .A2(new_n302_), .ZN(new_n313_));
  AND2_X1   g112(.A1(new_n289_), .A2(new_n290_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n235_), .A2(new_n277_), .ZN(new_n315_));
  NOR3_X1   g114(.A1(new_n280_), .A2(new_n281_), .A3(new_n234_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  OAI211_X1 g116(.A(KEYINPUT86), .B(new_n313_), .C1(new_n314_), .C2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n304_), .A2(new_n312_), .A3(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G226gat), .A2(G233gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT19), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  AOI211_X1 g121(.A(new_n305_), .B(new_n321_), .C1(new_n239_), .C2(new_n313_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n291_), .A2(new_n303_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(KEYINPUT87), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT87), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n291_), .A2(new_n326_), .A3(new_n303_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n323_), .A2(new_n325_), .A3(new_n327_), .ZN(new_n328_));
  XOR2_X1   g127(.A(G8gat), .B(G36gat), .Z(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT88), .B(KEYINPUT18), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G64gat), .B(G92gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  AND3_X1   g132(.A1(new_n322_), .A2(new_n328_), .A3(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n333_), .B1(new_n322_), .B2(new_n328_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n272_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G1gat), .B(G29gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(G85gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT0), .B(G57gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G225gat), .A2(G233gat), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT81), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT3), .ZN(new_n345_));
  INV_X1    g144(.A(G141gat), .ZN(new_n346_));
  INV_X1    g145(.A(G148gat), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n344_), .A2(new_n345_), .A3(new_n346_), .A4(new_n347_), .ZN(new_n348_));
  OAI22_X1  g147(.A1(KEYINPUT81), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G141gat), .A2(G148gat), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT2), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n353_));
  NAND4_X1  g152(.A1(new_n348_), .A2(new_n349_), .A3(new_n352_), .A4(new_n353_), .ZN(new_n354_));
  OR2_X1    g153(.A1(G155gat), .A2(G162gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G155gat), .A2(G162gat), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n354_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n346_), .A2(new_n347_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n360_));
  AND3_X1   g159(.A1(new_n359_), .A2(new_n360_), .A3(new_n350_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT1), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n355_), .A2(new_n362_), .A3(new_n356_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n361_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n358_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(new_n260_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n343_), .B1(new_n366_), .B2(KEYINPUT4), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT90), .ZN(new_n369_));
  AND3_X1   g168(.A1(new_n358_), .A2(new_n259_), .A3(new_n364_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n259_), .B1(new_n364_), .B2(new_n358_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n369_), .B1(new_n372_), .B2(KEYINPUT4), .ZN(new_n373_));
  AOI22_X1  g172(.A1(new_n354_), .A2(new_n357_), .B1(new_n361_), .B2(new_n363_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(new_n259_), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n366_), .A2(new_n369_), .A3(new_n375_), .A4(KEYINPUT4), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n368_), .B1(new_n373_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n372_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n379_), .A2(new_n343_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n341_), .B1(new_n378_), .B2(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n366_), .A2(KEYINPUT4), .A3(new_n375_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(KEYINPUT90), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n367_), .B1(new_n384_), .B2(new_n376_), .ZN(new_n385_));
  NOR3_X1   g184(.A1(new_n385_), .A2(new_n340_), .A3(new_n380_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n382_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G228gat), .A2(G233gat), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT82), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT29), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n391_), .B1(new_n358_), .B2(new_n364_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n390_), .B1(new_n392_), .B2(new_n303_), .ZN(new_n393_));
  OAI221_X1 g192(.A(new_n313_), .B1(new_n389_), .B2(new_n388_), .C1(new_n374_), .C2(new_n391_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G78gat), .B(G106gat), .ZN(new_n396_));
  AOI21_X1  g195(.A(KEYINPUT83), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n374_), .A2(new_n391_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G22gat), .B(G50gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT28), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n398_), .B(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n396_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n402_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n403_));
  AND3_X1   g202(.A1(new_n393_), .A2(new_n394_), .A3(new_n402_), .ZN(new_n404_));
  OAI22_X1  g203(.A1(new_n397_), .A2(new_n401_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n403_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n401_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n393_), .A2(new_n394_), .A3(new_n402_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n406_), .A2(new_n407_), .A3(KEYINPUT83), .A4(new_n408_), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n405_), .A2(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(KEYINPUT20), .B1(new_n311_), .B2(new_n303_), .ZN(new_n411_));
  NOR3_X1   g210(.A1(new_n314_), .A2(new_n317_), .A3(new_n313_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n321_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n413_), .B1(new_n319_), .B2(new_n321_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n333_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n322_), .A2(new_n328_), .A3(new_n333_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n416_), .A2(new_n417_), .A3(KEYINPUT27), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n336_), .A2(new_n387_), .A3(new_n410_), .A4(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT92), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n378_), .A2(new_n341_), .A3(new_n381_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n340_), .B1(new_n385_), .B2(new_n380_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n405_), .A2(new_n409_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT92), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n425_), .A2(new_n426_), .A3(new_n336_), .A4(new_n418_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n420_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n421_), .A2(KEYINPUT33), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT33), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n378_), .A2(new_n381_), .A3(new_n430_), .A4(new_n341_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n429_), .A2(new_n431_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n366_), .A2(KEYINPUT4), .ZN(new_n433_));
  AOI211_X1 g232(.A(new_n343_), .B(new_n433_), .C1(new_n384_), .C2(new_n376_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n340_), .B1(new_n379_), .B2(new_n342_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT89), .B1(new_n334_), .B2(new_n335_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n322_), .A2(new_n328_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(new_n415_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT89), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n440_), .A2(new_n441_), .A3(new_n417_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n432_), .A2(new_n437_), .A3(new_n438_), .A4(new_n442_), .ZN(new_n443_));
  AND2_X1   g242(.A1(new_n333_), .A2(KEYINPUT32), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n414_), .A2(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n445_), .B1(new_n439_), .B2(new_n444_), .ZN(new_n446_));
  OR2_X1    g245(.A1(new_n387_), .A2(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n410_), .B1(new_n443_), .B2(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n270_), .B1(new_n428_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n270_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n336_), .A2(new_n424_), .A3(new_n418_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT93), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n451_), .A2(KEYINPUT93), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n450_), .B(new_n387_), .C1(new_n453_), .C2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n449_), .A2(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G15gat), .B(G22gat), .ZN(new_n457_));
  INV_X1    g256(.A(G1gat), .ZN(new_n458_));
  INV_X1    g257(.A(G8gat), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT14), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT71), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n457_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  AND2_X1   g261(.A1(new_n460_), .A2(new_n461_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G1gat), .B(G8gat), .ZN(new_n464_));
  OR3_X1    g263(.A1(new_n462_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n464_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n466_));
  AND2_X1   g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G29gat), .B(G36gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(KEYINPUT69), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G43gat), .B(G50gat), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  OR2_X1    g271(.A1(new_n468_), .A2(KEYINPUT69), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n468_), .A2(KEYINPUT69), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n473_), .A2(new_n474_), .A3(new_n470_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n472_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n467_), .A2(new_n476_), .ZN(new_n477_));
  AND2_X1   g276(.A1(new_n472_), .A2(new_n475_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n465_), .A2(new_n466_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n481_), .A2(G229gat), .A3(G233gat), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT15), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n476_), .A2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n472_), .A2(KEYINPUT15), .A3(new_n475_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n484_), .A2(new_n479_), .A3(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G229gat), .A2(G233gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(KEYINPUT76), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n486_), .A2(new_n477_), .A3(new_n488_), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n482_), .A2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G113gat), .B(G141gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G169gat), .B(G197gat), .ZN(new_n492_));
  XOR2_X1   g291(.A(new_n491_), .B(new_n492_), .Z(new_n493_));
  OR2_X1    g292(.A1(new_n490_), .A2(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n482_), .A2(new_n489_), .A3(new_n493_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n456_), .A2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT94), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT12), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT9), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n500_), .A2(G85gat), .A3(G92gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(KEYINPUT10), .B(G99gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G85gat), .B(G92gat), .ZN(new_n503_));
  OAI221_X1 g302(.A(new_n501_), .B1(new_n502_), .B2(G106gat), .C1(new_n500_), .C2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G99gat), .A2(G106gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT6), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT6), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n507_), .A2(G99gat), .A3(G106gat), .ZN(new_n508_));
  AND3_X1   g307(.A1(new_n506_), .A2(new_n508_), .A3(KEYINPUT65), .ZN(new_n509_));
  AOI21_X1  g308(.A(KEYINPUT65), .B1(new_n506_), .B2(new_n508_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n504_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n506_), .A2(new_n508_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT66), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(G99gat), .A2(G106gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT7), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n506_), .A2(new_n508_), .A3(KEYINPUT66), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n515_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n503_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(KEYINPUT8), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n517_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n503_), .A2(KEYINPUT8), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n512_), .B1(new_n522_), .B2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G57gat), .B(G64gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G71gat), .B(G78gat), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n527_), .A2(new_n528_), .A3(KEYINPUT11), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(KEYINPUT11), .ZN(new_n530_));
  INV_X1    g329(.A(new_n528_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n527_), .A2(KEYINPUT11), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n529_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT67), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n499_), .B1(new_n526_), .B2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G230gat), .A2(G233gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT64), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n526_), .A2(new_n536_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n525_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT8), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n542_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n543_));
  OAI22_X1  g342(.A1(new_n541_), .A2(new_n543_), .B1(new_n511_), .B2(new_n504_), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n534_), .A2(new_n499_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(new_n546_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n537_), .A2(new_n539_), .A3(new_n540_), .A4(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT68), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n540_), .A2(new_n547_), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n551_), .A2(KEYINPUT68), .A3(new_n539_), .A4(new_n537_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n539_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n540_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n526_), .A2(new_n536_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n553_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n550_), .A2(new_n552_), .A3(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G120gat), .B(G148gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT5), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G176gat), .B(G204gat), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n559_), .B(new_n560_), .Z(new_n561_));
  NAND2_X1  g360(.A1(new_n557_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n561_), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n550_), .A2(new_n552_), .A3(new_n556_), .A4(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT13), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G183gat), .B(G211gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT73), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G127gat), .B(G155gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n571_));
  XOR2_X1   g370(.A(new_n570_), .B(new_n571_), .Z(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(KEYINPUT17), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(KEYINPUT74), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n570_), .B(new_n571_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT17), .ZN(new_n576_));
  OR3_X1    g375(.A1(new_n575_), .A2(KEYINPUT74), .A3(new_n576_), .ZN(new_n577_));
  AND2_X1   g376(.A1(G231gat), .A2(G233gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n479_), .B(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(new_n534_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n574_), .A2(new_n577_), .A3(new_n580_), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n579_), .A2(new_n536_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n579_), .A2(new_n536_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n575_), .A2(new_n576_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n573_), .A2(new_n582_), .A3(new_n583_), .A4(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n581_), .A2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT75), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n544_), .A2(new_n485_), .A3(new_n484_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n526_), .A2(new_n476_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G232gat), .A2(G233gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT34), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT35), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n589_), .A2(new_n590_), .A3(new_n595_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n593_), .A2(new_n594_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n597_), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n589_), .A2(new_n590_), .A3(new_n599_), .A4(new_n595_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT70), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  XOR2_X1   g402(.A(G190gat), .B(G218gat), .Z(new_n604_));
  XNOR2_X1  g403(.A(G134gat), .B(G162gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(KEYINPUT36), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n601_), .A2(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n607_), .A2(KEYINPUT36), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n603_), .A2(new_n610_), .A3(new_n612_), .ZN(new_n613_));
  OAI211_X1 g412(.A(new_n601_), .B(new_n602_), .C1(new_n611_), .C2(new_n609_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT37), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n613_), .A2(KEYINPUT37), .A3(new_n614_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  AND3_X1   g418(.A1(new_n566_), .A2(new_n588_), .A3(new_n619_), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n498_), .A2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n621_), .A2(new_n458_), .A3(new_n423_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT38), .ZN(new_n623_));
  OR2_X1    g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n566_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n496_), .ZN(new_n626_));
  NOR3_X1   g425(.A1(new_n625_), .A2(new_n626_), .A3(new_n587_), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n627_), .A2(KEYINPUT95), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n268_), .A2(new_n269_), .A3(new_n387_), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n451_), .A2(KEYINPUT93), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n629_), .B1(new_n630_), .B2(new_n452_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n387_), .A2(new_n446_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n438_), .A2(new_n442_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n436_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n632_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  OAI211_X1 g434(.A(new_n420_), .B(new_n427_), .C1(new_n635_), .C2(new_n410_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n631_), .B1(new_n636_), .B2(new_n270_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n637_), .A2(new_n615_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n627_), .A2(KEYINPUT95), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n628_), .A2(new_n638_), .A3(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(G1gat), .B1(new_n640_), .B2(new_n387_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n622_), .A2(new_n623_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n624_), .A2(new_n641_), .A3(new_n642_), .ZN(G1324gat));
  AND2_X1   g442(.A1(new_n336_), .A2(new_n418_), .ZN(new_n644_));
  OAI21_X1  g443(.A(G8gat), .B1(new_n640_), .B2(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT39), .ZN(new_n646_));
  INV_X1    g445(.A(new_n644_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n621_), .A2(new_n459_), .A3(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n649_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g449(.A(G15gat), .B1(new_n640_), .B2(new_n270_), .ZN(new_n651_));
  XOR2_X1   g450(.A(new_n651_), .B(KEYINPUT41), .Z(new_n652_));
  NAND3_X1  g451(.A1(new_n621_), .A2(new_n242_), .A3(new_n450_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1326gat));
  NOR2_X1   g453(.A1(new_n424_), .A2(G22gat), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT97), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n621_), .A2(new_n656_), .ZN(new_n657_));
  OAI21_X1  g456(.A(G22gat), .B1(new_n640_), .B2(new_n424_), .ZN(new_n658_));
  XOR2_X1   g457(.A(KEYINPUT96), .B(KEYINPUT42), .Z(new_n659_));
  AND2_X1   g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n658_), .A2(new_n659_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n657_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT98), .Z(G1327gat));
  XNOR2_X1  g462(.A(KEYINPUT103), .B(KEYINPUT44), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n625_), .A2(new_n626_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(new_n587_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT101), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT43), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n617_), .A2(new_n668_), .A3(new_n618_), .ZN(new_n669_));
  AOI211_X1 g468(.A(new_n667_), .B(new_n669_), .C1(new_n449_), .C2(new_n455_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n669_), .ZN(new_n671_));
  AOI21_X1  g470(.A(KEYINPUT101), .B1(new_n456_), .B2(new_n671_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n670_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n619_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n674_), .B1(new_n637_), .B2(KEYINPUT99), .ZN(new_n675_));
  AND3_X1   g474(.A1(new_n449_), .A2(KEYINPUT99), .A3(new_n455_), .ZN(new_n676_));
  OAI21_X1  g475(.A(KEYINPUT43), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT100), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n673_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT99), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n619_), .B1(new_n456_), .B2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n637_), .A2(KEYINPUT99), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n668_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(KEYINPUT100), .ZN(new_n684_));
  AOI211_X1 g483(.A(KEYINPUT102), .B(new_n666_), .C1(new_n679_), .C2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT102), .ZN(new_n686_));
  AOI21_X1  g485(.A(KEYINPUT99), .B1(new_n449_), .B2(new_n455_), .ZN(new_n687_));
  NOR3_X1   g486(.A1(new_n676_), .A2(new_n687_), .A3(new_n619_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n678_), .B1(new_n688_), .B2(new_n668_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n667_), .B1(new_n637_), .B2(new_n669_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n456_), .A2(KEYINPUT101), .A3(new_n671_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n689_), .A2(new_n684_), .A3(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n666_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n686_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n664_), .B1(new_n685_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT104), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n693_), .A2(KEYINPUT44), .A3(new_n694_), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n696_), .A2(new_n697_), .A3(new_n423_), .A4(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n664_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n692_), .B1(new_n683_), .B2(KEYINPUT100), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n688_), .A2(new_n678_), .A3(new_n668_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n694_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(KEYINPUT102), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n693_), .A2(new_n686_), .A3(new_n694_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n700_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n698_), .A2(new_n423_), .ZN(new_n707_));
  OAI21_X1  g506(.A(KEYINPUT104), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n699_), .A2(new_n708_), .A3(G29gat), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n587_), .A2(new_n615_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n625_), .A2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n498_), .A2(new_n711_), .ZN(new_n712_));
  OR3_X1    g511(.A1(new_n712_), .A2(G29gat), .A3(new_n387_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n709_), .A2(new_n713_), .ZN(G1328gat));
  INV_X1    g513(.A(KEYINPUT46), .ZN(new_n715_));
  INV_X1    g514(.A(G36gat), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n698_), .A2(new_n647_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n716_), .B1(new_n696_), .B2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n712_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n720_), .A2(new_n716_), .A3(new_n647_), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT45), .Z(new_n722_));
  OAI21_X1  g521(.A(new_n715_), .B1(new_n719_), .B2(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(G36gat), .B1(new_n706_), .B2(new_n717_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n721_), .B(KEYINPUT45), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n724_), .A2(KEYINPUT46), .A3(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n723_), .A2(new_n726_), .ZN(G1329gat));
  AND3_X1   g526(.A1(new_n693_), .A2(KEYINPUT44), .A3(new_n694_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n450_), .A2(G43gat), .ZN(new_n729_));
  NOR3_X1   g528(.A1(new_n706_), .A2(new_n728_), .A3(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(G43gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n731_), .B1(new_n712_), .B2(new_n270_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT105), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(KEYINPUT47), .B1(new_n730_), .B2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT47), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n696_), .A2(new_n698_), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n736_), .B(new_n733_), .C1(new_n737_), .C2(new_n729_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n735_), .A2(new_n738_), .ZN(G1330gat));
  AOI21_X1  g538(.A(G50gat), .B1(new_n720_), .B2(new_n410_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n737_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n410_), .A2(G50gat), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n740_), .B1(new_n741_), .B2(new_n742_), .ZN(G1331gat));
  NOR2_X1   g542(.A1(new_n566_), .A2(new_n496_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n638_), .A2(new_n588_), .A3(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(G57gat), .B1(new_n745_), .B2(new_n387_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n637_), .A2(new_n496_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n587_), .B1(new_n618_), .B2(new_n617_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n747_), .A2(new_n625_), .A3(new_n748_), .ZN(new_n749_));
  OR2_X1    g548(.A1(new_n387_), .A2(G57gat), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n746_), .B1(new_n749_), .B2(new_n750_), .ZN(G1332gat));
  OAI21_X1  g550(.A(G64gat), .B1(new_n745_), .B2(new_n644_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT48), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n644_), .A2(G64gat), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT106), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n753_), .B1(new_n749_), .B2(new_n755_), .ZN(G1333gat));
  OAI21_X1  g555(.A(G71gat), .B1(new_n745_), .B2(new_n270_), .ZN(new_n757_));
  XOR2_X1   g556(.A(KEYINPUT107), .B(KEYINPUT49), .Z(new_n758_));
  XNOR2_X1  g557(.A(new_n757_), .B(new_n758_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n270_), .A2(G71gat), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT108), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n759_), .B1(new_n749_), .B2(new_n761_), .ZN(G1334gat));
  OAI21_X1  g561(.A(G78gat), .B1(new_n745_), .B2(new_n424_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT50), .ZN(new_n764_));
  OR2_X1    g563(.A1(new_n424_), .A2(G78gat), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n764_), .B1(new_n749_), .B2(new_n765_), .ZN(G1335gat));
  INV_X1    g565(.A(G85gat), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n744_), .A2(new_n587_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n768_), .B1(new_n679_), .B2(new_n684_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n767_), .B1(new_n769_), .B2(new_n423_), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n747_), .A2(new_n625_), .A3(new_n587_), .A4(new_n615_), .ZN(new_n771_));
  NOR3_X1   g570(.A1(new_n771_), .A2(G85gat), .A3(new_n387_), .ZN(new_n772_));
  OR2_X1    g571(.A1(new_n770_), .A2(new_n772_), .ZN(G1336gat));
  INV_X1    g572(.A(G92gat), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n774_), .B1(new_n769_), .B2(new_n647_), .ZN(new_n775_));
  NOR3_X1   g574(.A1(new_n771_), .A2(G92gat), .A3(new_n644_), .ZN(new_n776_));
  OR2_X1    g575(.A1(new_n775_), .A2(new_n776_), .ZN(G1337gat));
  NOR3_X1   g576(.A1(new_n771_), .A2(new_n270_), .A3(new_n502_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n769_), .A2(new_n450_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n778_), .B1(new_n779_), .B2(G99gat), .ZN(new_n780_));
  XOR2_X1   g579(.A(new_n780_), .B(KEYINPUT51), .Z(G1338gat));
  OR3_X1    g580(.A1(new_n771_), .A2(G106gat), .A3(new_n424_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n768_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n693_), .A2(new_n410_), .A3(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n785_));
  AND3_X1   g584(.A1(new_n784_), .A2(new_n785_), .A3(G106gat), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n785_), .B1(new_n784_), .B2(G106gat), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n782_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT53), .ZN(G1339gat));
  AOI21_X1  g588(.A(new_n488_), .B1(new_n467_), .B2(new_n476_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n493_), .B1(new_n790_), .B2(new_n486_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n481_), .A2(new_n488_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT110), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n791_), .A2(new_n792_), .A3(KEYINPUT110), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n795_), .A2(new_n495_), .A3(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT111), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT111), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n795_), .A2(new_n799_), .A3(new_n495_), .A4(new_n796_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n798_), .A2(new_n800_), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n801_), .A2(new_n564_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n548_), .A2(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n539_), .B1(new_n551_), .B2(new_n537_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n550_), .A2(new_n552_), .A3(new_n803_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(KEYINPUT56), .B1(new_n808_), .B2(new_n561_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT56), .ZN(new_n810_));
  AOI211_X1 g609(.A(new_n810_), .B(new_n563_), .C1(new_n806_), .C2(new_n807_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n802_), .B1(new_n809_), .B2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT58), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n802_), .B(KEYINPUT58), .C1(new_n809_), .C2(new_n811_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n814_), .A2(new_n674_), .A3(new_n815_), .ZN(new_n816_));
  AND2_X1   g615(.A1(new_n496_), .A2(new_n564_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n817_), .B1(new_n809_), .B2(new_n811_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n801_), .A2(new_n565_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n615_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(KEYINPUT112), .A2(KEYINPUT57), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n821_), .ZN(new_n823_));
  AOI211_X1 g622(.A(new_n615_), .B(new_n823_), .C1(new_n818_), .C2(new_n819_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n816_), .B1(new_n822_), .B2(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n588_), .B1(new_n825_), .B2(KEYINPUT113), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT113), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n816_), .B(new_n827_), .C1(new_n822_), .C2(new_n824_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n620_), .A2(KEYINPUT109), .A3(new_n830_), .A4(new_n626_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n748_), .A2(new_n566_), .A3(new_n830_), .A4(new_n626_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT109), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n748_), .A2(new_n626_), .A3(new_n566_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT54), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n831_), .A2(new_n834_), .A3(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n829_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT114), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n453_), .A2(new_n454_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n450_), .A2(new_n423_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n838_), .A2(new_n839_), .A3(new_n842_), .ZN(new_n843_));
  AND3_X1   g642(.A1(new_n831_), .A2(new_n834_), .A3(new_n836_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n844_), .B1(new_n826_), .B2(new_n828_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n842_), .ZN(new_n846_));
  OAI21_X1  g645(.A(KEYINPUT114), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n843_), .A2(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(G113gat), .B1(new_n848_), .B2(new_n496_), .ZN(new_n849_));
  OAI21_X1  g648(.A(KEYINPUT59), .B1(new_n845_), .B2(new_n846_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n825_), .A2(new_n587_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT116), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n825_), .A2(KEYINPUT116), .A3(new_n587_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(new_n837_), .A3(new_n854_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(KEYINPUT115), .B(KEYINPUT59), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n846_), .A2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n850_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n496_), .A2(G113gat), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(KEYINPUT117), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n849_), .B1(new_n860_), .B2(new_n862_), .ZN(G1340gat));
  XNOR2_X1  g662(.A(KEYINPUT118), .B(G120gat), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n864_), .B1(new_n566_), .B2(KEYINPUT60), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n864_), .A2(KEYINPUT60), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(KEYINPUT119), .B2(new_n866_), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n848_), .B(new_n867_), .C1(KEYINPUT119), .C2(new_n865_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n859_), .A2(new_n566_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n868_), .B1(new_n869_), .B2(new_n864_), .ZN(G1341gat));
  NAND3_X1  g669(.A1(new_n843_), .A2(new_n588_), .A3(new_n847_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n249_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT120), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n871_), .A2(KEYINPUT120), .A3(new_n249_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n587_), .A2(new_n249_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(KEYINPUT121), .ZN(new_n877_));
  AOI22_X1  g676(.A1(new_n874_), .A2(new_n875_), .B1(new_n860_), .B2(new_n877_), .ZN(G1342gat));
  NAND3_X1  g677(.A1(new_n850_), .A2(new_n674_), .A3(new_n858_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(G134gat), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n843_), .A2(new_n847_), .A3(new_n247_), .A4(new_n615_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT122), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n880_), .A2(KEYINPUT122), .A3(new_n881_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(G1343gat));
  NOR4_X1   g685(.A1(new_n450_), .A2(new_n647_), .A3(new_n424_), .A4(new_n387_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n838_), .A2(new_n887_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n888_), .A2(new_n626_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(new_n346_), .ZN(G1344gat));
  NOR2_X1   g689(.A1(new_n888_), .A2(new_n566_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(new_n347_), .ZN(G1345gat));
  OR3_X1    g691(.A1(new_n888_), .A2(KEYINPUT123), .A3(new_n587_), .ZN(new_n893_));
  OAI21_X1  g692(.A(KEYINPUT123), .B1(new_n888_), .B2(new_n587_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(KEYINPUT61), .B(G155gat), .ZN(new_n895_));
  AND3_X1   g694(.A1(new_n893_), .A2(new_n894_), .A3(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n895_), .B1(new_n893_), .B2(new_n894_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n896_), .A2(new_n897_), .ZN(G1346gat));
  OAI21_X1  g697(.A(G162gat), .B1(new_n888_), .B2(new_n619_), .ZN(new_n899_));
  INV_X1    g698(.A(G162gat), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n615_), .A2(new_n900_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n899_), .B1(new_n888_), .B2(new_n901_), .ZN(G1347gat));
  NOR2_X1   g701(.A1(new_n629_), .A2(new_n644_), .ZN(new_n903_));
  AND3_X1   g702(.A1(new_n855_), .A2(new_n424_), .A3(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n496_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(G169gat), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT62), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n905_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n909_));
  AND2_X1   g708(.A1(new_n286_), .A2(new_n288_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  OAI211_X1 g710(.A(new_n908_), .B(new_n909_), .C1(new_n911_), .C2(new_n905_), .ZN(G1348gat));
  NAND2_X1  g711(.A1(new_n904_), .A2(new_n625_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n845_), .A2(new_n410_), .ZN(new_n914_));
  AND3_X1   g713(.A1(new_n625_), .A2(G176gat), .A3(new_n903_), .ZN(new_n915_));
  AOI22_X1  g714(.A1(new_n913_), .A2(new_n287_), .B1(new_n914_), .B2(new_n915_), .ZN(G1349gat));
  NAND3_X1  g715(.A1(new_n914_), .A2(new_n588_), .A3(new_n903_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n587_), .B1(new_n274_), .B2(new_n223_), .ZN(new_n918_));
  AOI22_X1  g717(.A1(new_n917_), .A2(new_n221_), .B1(new_n904_), .B2(new_n918_), .ZN(G1350gat));
  NAND2_X1  g718(.A1(new_n275_), .A2(new_n276_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n920_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n904_), .A2(new_n921_), .A3(new_n615_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n922_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n227_), .B1(new_n904_), .B2(new_n674_), .ZN(new_n924_));
  OAI21_X1  g723(.A(KEYINPUT124), .B1(new_n923_), .B2(new_n924_), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT124), .ZN(new_n926_));
  AND2_X1   g725(.A1(new_n904_), .A2(new_n674_), .ZN(new_n927_));
  OAI211_X1 g726(.A(new_n926_), .B(new_n922_), .C1(new_n927_), .C2(new_n227_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n925_), .A2(new_n928_), .ZN(G1351gat));
  NAND2_X1  g728(.A1(new_n270_), .A2(new_n425_), .ZN(new_n930_));
  INV_X1    g729(.A(new_n930_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n931_), .A2(KEYINPUT125), .ZN(new_n932_));
  AND2_X1   g731(.A1(new_n931_), .A2(KEYINPUT125), .ZN(new_n933_));
  NOR4_X1   g732(.A1(new_n845_), .A2(new_n644_), .A3(new_n932_), .A4(new_n933_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(new_n496_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g735(.A1(new_n934_), .A2(new_n625_), .ZN(new_n937_));
  INV_X1    g736(.A(G204gat), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n938_), .A2(KEYINPUT126), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n937_), .B(new_n939_), .ZN(G1353gat));
  INV_X1    g739(.A(KEYINPUT63), .ZN(new_n941_));
  INV_X1    g740(.A(G211gat), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n941_), .A2(new_n942_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n944_));
  AND4_X1   g743(.A1(new_n588_), .A2(new_n934_), .A3(new_n943_), .A4(new_n944_), .ZN(new_n945_));
  INV_X1    g744(.A(KEYINPUT127), .ZN(new_n946_));
  AND2_X1   g745(.A1(new_n934_), .A2(new_n588_), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n946_), .B1(new_n947_), .B2(new_n943_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n934_), .A2(new_n588_), .ZN(new_n949_));
  NAND4_X1  g748(.A1(new_n949_), .A2(KEYINPUT127), .A3(new_n941_), .A4(new_n942_), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n945_), .B1(new_n948_), .B2(new_n950_), .ZN(G1354gat));
  INV_X1    g750(.A(G218gat), .ZN(new_n952_));
  NAND3_X1  g751(.A1(new_n934_), .A2(new_n952_), .A3(new_n615_), .ZN(new_n953_));
  AND2_X1   g752(.A1(new_n934_), .A2(new_n674_), .ZN(new_n954_));
  OAI21_X1  g753(.A(new_n953_), .B1(new_n954_), .B2(new_n952_), .ZN(G1355gat));
endmodule


