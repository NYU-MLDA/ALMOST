//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 0 0 1 0 0 0 0 0 1 0 1 0 1 1 1 0 1 1 0 1 1 0 0 1 1 1 1 1 0 0 0 0 1 1 1 0 1 0 1 0 0 1 1 1 0 0 1 1 0 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n614_, new_n615_, new_n616_, new_n617_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n673_, new_n674_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n836_, new_n837_, new_n839_, new_n840_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n867_, new_n868_, new_n870_,
    new_n871_, new_n872_, new_n874_, new_n875_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n887_;
  INV_X1    g000(.A(KEYINPUT81), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G232gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT34), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT35), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT75), .ZN(new_n206_));
  XOR2_X1   g005(.A(G85gat), .B(G92gat), .Z(new_n207_));
  INV_X1    g006(.A(KEYINPUT68), .ZN(new_n208_));
  OAI221_X1 g007(.A(new_n208_), .B1(KEYINPUT69), .B2(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n209_));
  NOR2_X1   g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(KEYINPUT69), .A2(KEYINPUT7), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n210_), .B1(new_n211_), .B2(KEYINPUT68), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n209_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G99gat), .A2(G106gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT6), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n216_), .B(new_n217_), .C1(new_n208_), .C2(KEYINPUT7), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n207_), .B1(new_n213_), .B2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT8), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT8), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n221_), .B(new_n207_), .C1(new_n213_), .C2(new_n218_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n216_), .A2(new_n217_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT10), .B(G99gat), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT64), .B1(new_n225_), .B2(G106gat), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT64), .ZN(new_n227_));
  INV_X1    g026(.A(G106gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT10), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n229_), .A2(G99gat), .ZN(new_n230_));
  INV_X1    g029(.A(G99gat), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n231_), .A2(KEYINPUT10), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n227_), .B(new_n228_), .C1(new_n230_), .C2(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n224_), .B1(new_n226_), .B2(new_n233_), .ZN(new_n234_));
  OR2_X1    g033(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n235_));
  OR2_X1    g034(.A1(KEYINPUT66), .A2(G92gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(KEYINPUT66), .A2(G92gat), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .A4(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT9), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  AND3_X1   g040(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n242_));
  NOR2_X1   g041(.A1(G85gat), .A2(G92gat), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n241_), .A2(new_n244_), .ZN(new_n245_));
  AND3_X1   g044(.A1(new_n234_), .A2(KEYINPUT67), .A3(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(KEYINPUT67), .B1(new_n234_), .B2(new_n245_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n223_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G29gat), .B(G36gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G43gat), .B(G50gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  OAI22_X1  g051(.A1(new_n248_), .A2(new_n252_), .B1(KEYINPUT35), .B2(new_n204_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n251_), .B(KEYINPUT15), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n248_), .A2(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n206_), .B1(new_n253_), .B2(new_n255_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n205_), .A2(KEYINPUT75), .ZN(new_n257_));
  OR2_X1    g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n257_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n258_), .A2(KEYINPUT36), .A3(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G134gat), .B(G162gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(G218gat), .ZN(new_n262_));
  XOR2_X1   g061(.A(KEYINPUT76), .B(G190gat), .Z(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n260_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT36), .ZN(new_n266_));
  OR2_X1    g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT77), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n258_), .A2(new_n269_), .A3(new_n259_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n268_), .A2(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n265_), .A2(new_n270_), .A3(new_n267_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n272_), .A2(KEYINPUT78), .A3(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT37), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n272_), .A2(KEYINPUT78), .A3(KEYINPUT37), .A4(new_n273_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT74), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT71), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G57gat), .B(G64gat), .ZN(new_n282_));
  OR2_X1    g081(.A1(new_n282_), .A2(KEYINPUT11), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(KEYINPUT11), .ZN(new_n284_));
  XOR2_X1   g083(.A(G71gat), .B(G78gat), .Z(new_n285_));
  NAND3_X1  g084(.A1(new_n283_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  OR2_X1    g085(.A1(new_n284_), .A2(new_n285_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n288_), .B(new_n223_), .C1(new_n246_), .C2(new_n247_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT70), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G230gat), .A2(G233gat), .ZN(new_n291_));
  AND3_X1   g090(.A1(new_n289_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n290_), .B1(new_n289_), .B2(new_n291_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT12), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT67), .ZN(new_n296_));
  INV_X1    g095(.A(new_n224_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n233_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n231_), .A2(KEYINPUT10), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n229_), .A2(G99gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n227_), .B1(new_n301_), .B2(new_n228_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n297_), .B1(new_n298_), .B2(new_n302_), .ZN(new_n303_));
  AOI211_X1 g102(.A(new_n243_), .B(new_n242_), .C1(new_n239_), .C2(new_n240_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n296_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n234_), .A2(new_n245_), .A3(KEYINPUT67), .ZN(new_n306_));
  AOI22_X1  g105(.A1(new_n305_), .A2(new_n306_), .B1(new_n220_), .B2(new_n222_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n295_), .B1(new_n307_), .B2(new_n288_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n288_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n248_), .A2(KEYINPUT12), .A3(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n281_), .B1(new_n294_), .B2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n289_), .A2(new_n291_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT70), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n289_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  AND3_X1   g115(.A1(new_n248_), .A2(KEYINPUT12), .A3(new_n309_), .ZN(new_n317_));
  AOI21_X1  g116(.A(KEYINPUT12), .B1(new_n248_), .B2(new_n309_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n316_), .A2(new_n319_), .A3(KEYINPUT71), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n312_), .A2(new_n320_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n307_), .A2(new_n288_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n289_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n321_), .B1(new_n291_), .B2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT73), .B(G120gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G176gat), .B(G204gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(G148gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n328_), .B(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n325_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n325_), .A2(new_n331_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n280_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n325_), .A2(new_n331_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n336_), .A2(KEYINPUT74), .A3(new_n332_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n335_), .A2(new_n337_), .A3(KEYINPUT13), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT13), .ZN(new_n339_));
  NOR3_X1   g138(.A1(new_n333_), .A2(new_n334_), .A3(new_n280_), .ZN(new_n340_));
  AOI21_X1  g139(.A(KEYINPUT74), .B1(new_n336_), .B2(new_n332_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n339_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G231gat), .A2(G233gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n288_), .B(new_n343_), .ZN(new_n344_));
  XOR2_X1   g143(.A(G15gat), .B(G22gat), .Z(new_n345_));
  XOR2_X1   g144(.A(KEYINPUT79), .B(G1gat), .Z(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(G8gat), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n345_), .B1(new_n347_), .B2(KEYINPUT14), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G1gat), .B(G8gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n344_), .B(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT80), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G127gat), .B(G155gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(G211gat), .ZN(new_n354_));
  XOR2_X1   g153(.A(KEYINPUT16), .B(G183gat), .Z(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT17), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  XOR2_X1   g157(.A(new_n352_), .B(new_n358_), .Z(new_n359_));
  INV_X1    g158(.A(new_n351_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n360_), .A2(new_n357_), .A3(new_n356_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n279_), .A2(new_n338_), .A3(new_n342_), .A4(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G57gat), .B(G85gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT101), .B(KEYINPUT0), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G1gat), .B(G29gat), .ZN(new_n367_));
  XOR2_X1   g166(.A(new_n366_), .B(new_n367_), .Z(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  AND2_X1   g168(.A1(G155gat), .A2(G162gat), .ZN(new_n370_));
  INV_X1    g169(.A(G141gat), .ZN(new_n371_));
  INV_X1    g170(.A(G148gat), .ZN(new_n372_));
  AOI22_X1  g171(.A1(new_n370_), .A2(KEYINPUT1), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G155gat), .B(G162gat), .ZN(new_n374_));
  OAI221_X1 g173(.A(new_n373_), .B1(new_n371_), .B2(new_n372_), .C1(KEYINPUT1), .C2(new_n374_), .ZN(new_n375_));
  OR3_X1    g174(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT2), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n377_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n379_));
  OAI21_X1  g178(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n376_), .A2(new_n378_), .A3(new_n379_), .A4(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n374_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n375_), .A2(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G127gat), .B(G134gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(KEYINPUT91), .ZN(new_n386_));
  XOR2_X1   g185(.A(G113gat), .B(G120gat), .Z(new_n387_));
  NOR2_X1   g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n388_), .A2(KEYINPUT92), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n386_), .A2(new_n387_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n386_), .A2(KEYINPUT92), .A3(new_n387_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n384_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n393_), .A2(KEYINPUT4), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT99), .ZN(new_n395_));
  OR2_X1    g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n386_), .A2(new_n387_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n384_), .B1(new_n397_), .B2(new_n388_), .ZN(new_n398_));
  OR2_X1    g197(.A1(new_n398_), .A2(KEYINPUT100), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n393_), .A2(new_n395_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n398_), .A2(KEYINPUT100), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n396_), .A2(new_n399_), .A3(new_n400_), .A4(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n394_), .B1(new_n402_), .B2(KEYINPUT4), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G225gat), .A2(G233gat), .ZN(new_n404_));
  OR2_X1    g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n402_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(new_n404_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n369_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n407_), .B(new_n369_), .C1(new_n403_), .C2(new_n404_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n408_), .A2(new_n410_), .ZN(new_n411_));
  XOR2_X1   g210(.A(G78gat), .B(G106gat), .Z(new_n412_));
  INV_X1    g211(.A(G204gat), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n413_), .A2(KEYINPUT94), .A3(G197gat), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT94), .ZN(new_n415_));
  INV_X1    g214(.A(G197gat), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n415_), .B1(new_n416_), .B2(G204gat), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n416_), .A2(G204gat), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n414_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  OR2_X1    g218(.A1(new_n419_), .A2(KEYINPUT21), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(KEYINPUT95), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n413_), .A2(G197gat), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT21), .B1(new_n418_), .B2(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G211gat), .B(G218gat), .ZN(new_n424_));
  XOR2_X1   g223(.A(new_n424_), .B(KEYINPUT96), .Z(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n421_), .A2(new_n423_), .A3(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n425_), .A2(KEYINPUT21), .A3(new_n419_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT29), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n429_), .B1(new_n430_), .B2(new_n384_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(KEYINPUT93), .A2(G233gat), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(KEYINPUT93), .A2(G233gat), .ZN(new_n435_));
  OAI21_X1  g234(.A(G228gat), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  OR2_X1    g235(.A1(new_n432_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n432_), .A2(new_n436_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n412_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n437_), .A2(new_n438_), .A3(new_n412_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n384_), .A2(new_n430_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(KEYINPUT28), .B(G22gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(G50gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n443_), .B(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n446_), .B1(new_n439_), .B2(KEYINPUT97), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n442_), .A2(new_n447_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n440_), .A2(KEYINPUT97), .A3(new_n441_), .A4(new_n446_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(KEYINPUT88), .B(G176gat), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT87), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT22), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n451_), .B1(new_n452_), .B2(G169gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(KEYINPUT22), .B(G169gat), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n450_), .B(new_n453_), .C1(new_n454_), .C2(new_n451_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G169gat), .A2(G176gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G183gat), .A2(G190gat), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT23), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n457_), .B(KEYINPUT86), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n459_), .B1(new_n460_), .B2(new_n458_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(G183gat), .A2(G190gat), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n455_), .B(new_n456_), .C1(new_n461_), .C2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n460_), .A2(new_n458_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n464_), .B1(new_n458_), .B2(new_n457_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n456_), .A2(KEYINPUT24), .ZN(new_n466_));
  NOR2_X1   g265(.A1(G169gat), .A2(G176gat), .ZN(new_n467_));
  MUX2_X1   g266(.A(new_n466_), .B(KEYINPUT24), .S(new_n467_), .Z(new_n468_));
  INV_X1    g267(.A(G190gat), .ZN(new_n469_));
  OR3_X1    g268(.A1(new_n469_), .A2(KEYINPUT85), .A3(KEYINPUT26), .ZN(new_n470_));
  XNOR2_X1  g269(.A(KEYINPUT25), .B(G183gat), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT26), .B1(new_n469_), .B2(KEYINPUT85), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n470_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n468_), .A2(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n463_), .B1(new_n465_), .B2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT89), .B(KEYINPUT30), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT90), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G15gat), .B(G43gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G227gat), .A2(G233gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G71gat), .B(G99gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n479_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT31), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT31), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n479_), .A2(new_n487_), .A3(new_n484_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n489_), .A2(new_n392_), .A3(new_n391_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n477_), .A2(new_n478_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n391_), .A2(new_n392_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n486_), .A2(new_n492_), .A3(new_n488_), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n490_), .A2(new_n491_), .A3(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n491_), .B1(new_n490_), .B2(new_n493_), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n448_), .B(new_n449_), .C1(new_n494_), .C2(new_n495_), .ZN(new_n496_));
  OR2_X1    g295(.A1(new_n429_), .A2(new_n475_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G226gat), .A2(G233gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT19), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n456_), .B1(new_n465_), .B2(new_n462_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n500_), .B1(new_n450_), .B2(new_n454_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n471_), .ZN(new_n502_));
  XOR2_X1   g301(.A(KEYINPUT26), .B(G190gat), .Z(new_n503_));
  OAI21_X1  g302(.A(new_n468_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n504_), .A2(new_n461_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n429_), .B1(new_n501_), .B2(new_n505_), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n497_), .A2(KEYINPUT20), .A3(new_n499_), .A4(new_n506_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n501_), .A2(new_n505_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n508_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n429_), .A2(new_n475_), .ZN(new_n510_));
  AND3_X1   g309(.A1(new_n509_), .A2(KEYINPUT20), .A3(new_n510_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n507_), .B1(new_n511_), .B2(new_n499_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G8gat), .B(G36gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(G92gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(KEYINPUT18), .B(G64gat), .ZN(new_n515_));
  XOR2_X1   g314(.A(new_n514_), .B(new_n515_), .Z(new_n516_));
  NAND2_X1  g315(.A1(new_n512_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT98), .ZN(new_n518_));
  INV_X1    g317(.A(new_n516_), .ZN(new_n519_));
  OAI211_X1 g318(.A(new_n507_), .B(new_n519_), .C1(new_n511_), .C2(new_n499_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n517_), .A2(new_n518_), .A3(new_n520_), .ZN(new_n521_));
  XOR2_X1   g320(.A(KEYINPUT104), .B(KEYINPUT27), .Z(new_n522_));
  NAND3_X1  g321(.A1(new_n512_), .A2(KEYINPUT98), .A3(new_n516_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n521_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n497_), .A2(KEYINPUT20), .A3(new_n506_), .ZN(new_n525_));
  MUX2_X1   g324(.A(new_n525_), .B(new_n511_), .S(new_n499_), .Z(new_n526_));
  OAI211_X1 g325(.A(new_n517_), .B(KEYINPUT27), .C1(new_n526_), .C2(new_n516_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n524_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT105), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT105), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n524_), .A2(new_n530_), .A3(new_n527_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n496_), .B1(new_n529_), .B2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n448_), .A2(new_n449_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n494_), .A2(new_n495_), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n533_), .A2(new_n534_), .A3(new_n524_), .A4(new_n527_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n411_), .B1(new_n532_), .B2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n516_), .A2(KEYINPUT32), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n512_), .A2(new_n538_), .ZN(new_n539_));
  OAI221_X1 g338(.A(new_n539_), .B1(new_n526_), .B2(new_n538_), .C1(new_n408_), .C2(new_n410_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(KEYINPUT102), .A2(KEYINPUT33), .ZN(new_n541_));
  NAND2_X1  g340(.A1(KEYINPUT102), .A2(KEYINPUT33), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n541_), .B1(new_n409_), .B2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n521_), .A2(new_n523_), .ZN(new_n544_));
  OAI211_X1 g343(.A(new_n543_), .B(new_n544_), .C1(new_n409_), .C2(new_n542_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n404_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n406_), .A2(new_n546_), .ZN(new_n547_));
  OAI211_X1 g346(.A(new_n547_), .B(new_n368_), .C1(new_n403_), .C2(new_n546_), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n548_), .B(KEYINPUT103), .Z(new_n549_));
  OAI21_X1  g348(.A(new_n540_), .B1(new_n545_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n533_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n550_), .A2(new_n551_), .A3(new_n534_), .ZN(new_n552_));
  AOI22_X1  g351(.A1(new_n202_), .A2(new_n363_), .B1(new_n537_), .B2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n350_), .A2(new_n251_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n349_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n348_), .B(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(new_n254_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G229gat), .A2(G233gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT82), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n554_), .A2(new_n557_), .A3(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT83), .ZN(new_n561_));
  OR2_X1    g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n556_), .A2(new_n252_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n554_), .A2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n564_), .A2(G229gat), .A3(G233gat), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n560_), .A2(new_n561_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G113gat), .B(G141gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G169gat), .B(G197gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n562_), .A2(new_n565_), .A3(new_n566_), .A4(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT84), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n562_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(new_n569_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n572_), .B(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n342_), .A2(new_n338_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n362_), .ZN(new_n578_));
  NOR3_X1   g377(.A1(new_n577_), .A2(new_n278_), .A3(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n576_), .B1(new_n579_), .B2(KEYINPUT81), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n553_), .A2(new_n580_), .ZN(new_n581_));
  NOR3_X1   g380(.A1(new_n581_), .A2(new_n411_), .A3(new_n346_), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n582_), .B(KEYINPUT38), .Z(new_n583_));
  NAND2_X1  g382(.A1(new_n537_), .A2(new_n552_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n272_), .A2(new_n273_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n584_), .A2(new_n585_), .A3(new_n362_), .ZN(new_n586_));
  NOR3_X1   g385(.A1(new_n586_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(G1gat), .B1(new_n588_), .B2(new_n411_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n583_), .A2(new_n589_), .ZN(G1324gat));
  NAND2_X1  g389(.A1(new_n529_), .A2(new_n531_), .ZN(new_n591_));
  NOR4_X1   g390(.A1(new_n586_), .A2(new_n576_), .A3(new_n577_), .A4(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT39), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n594_), .A2(KEYINPUT106), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(KEYINPUT106), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n593_), .A2(G8gat), .A3(new_n595_), .A4(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(G8gat), .ZN(new_n598_));
  INV_X1    g397(.A(new_n591_), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n553_), .A2(new_n598_), .A3(new_n580_), .A4(new_n599_), .ZN(new_n600_));
  OAI211_X1 g399(.A(KEYINPUT106), .B(new_n594_), .C1(new_n592_), .C2(new_n598_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n597_), .A2(new_n600_), .A3(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT40), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n597_), .A2(new_n601_), .A3(KEYINPUT40), .A4(new_n600_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(G1325gat));
  INV_X1    g405(.A(G15gat), .ZN(new_n607_));
  INV_X1    g406(.A(new_n534_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n607_), .B1(new_n587_), .B2(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT41), .ZN(new_n610_));
  NOR3_X1   g409(.A1(new_n581_), .A2(G15gat), .A3(new_n534_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT107), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(G1326gat));
  OR3_X1    g412(.A1(new_n581_), .A2(G22gat), .A3(new_n551_), .ZN(new_n614_));
  OAI21_X1  g413(.A(G22gat), .B1(new_n588_), .B2(new_n551_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n615_), .A2(KEYINPUT42), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n615_), .A2(KEYINPUT42), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n614_), .B1(new_n616_), .B2(new_n617_), .ZN(G1327gat));
  AOI21_X1  g417(.A(new_n585_), .B1(new_n537_), .B2(new_n552_), .ZN(new_n619_));
  NOR3_X1   g418(.A1(new_n577_), .A2(new_n576_), .A3(new_n362_), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n411_), .ZN(new_n622_));
  AOI21_X1  g421(.A(G29gat), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n279_), .A2(KEYINPUT43), .ZN(new_n624_));
  INV_X1    g423(.A(new_n496_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n531_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n530_), .B1(new_n524_), .B2(new_n527_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n625_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n622_), .B1(new_n628_), .B2(new_n535_), .ZN(new_n629_));
  AND3_X1   g428(.A1(new_n550_), .A2(new_n551_), .A3(new_n534_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n624_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n278_), .A2(KEYINPUT108), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT108), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n276_), .A2(new_n633_), .A3(new_n277_), .ZN(new_n634_));
  AOI22_X1  g433(.A1(new_n537_), .A2(new_n552_), .B1(new_n632_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT43), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n631_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(new_n620_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT44), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  AND3_X1   g439(.A1(new_n640_), .A2(G29gat), .A3(new_n622_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n637_), .A2(KEYINPUT44), .A3(new_n620_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n623_), .B1(new_n641_), .B2(new_n642_), .ZN(G1328gat));
  NAND3_X1  g442(.A1(new_n640_), .A2(new_n599_), .A3(new_n642_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(G36gat), .ZN(new_n645_));
  INV_X1    g444(.A(G36gat), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n591_), .B(KEYINPUT109), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n619_), .A2(new_n646_), .A3(new_n647_), .A4(new_n620_), .ZN(new_n648_));
  OR2_X1    g447(.A1(new_n648_), .A2(KEYINPUT110), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(KEYINPUT110), .ZN(new_n650_));
  XOR2_X1   g449(.A(KEYINPUT111), .B(KEYINPUT45), .Z(new_n651_));
  NAND3_X1  g450(.A1(new_n649_), .A2(new_n650_), .A3(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n651_), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n648_), .A2(KEYINPUT110), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n648_), .A2(KEYINPUT110), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n653_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n645_), .A2(KEYINPUT46), .A3(new_n652_), .A4(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT46), .ZN(new_n658_));
  AOI21_X1  g457(.A(KEYINPUT44), .B1(new_n637_), .B2(new_n620_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n659_), .A2(new_n591_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n646_), .B1(new_n660_), .B2(new_n642_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n656_), .A2(new_n652_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n658_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n657_), .A2(new_n663_), .ZN(G1329gat));
  AND2_X1   g463(.A1(new_n621_), .A2(new_n608_), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n665_), .A2(G43gat), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n642_), .A2(G43gat), .A3(new_n608_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n666_), .B1(new_n659_), .B2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(KEYINPUT47), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT47), .ZN(new_n670_));
  OAI211_X1 g469(.A(new_n666_), .B(new_n670_), .C1(new_n659_), .C2(new_n667_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(G1330gat));
  AOI21_X1  g471(.A(G50gat), .B1(new_n621_), .B2(new_n533_), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n640_), .A2(G50gat), .A3(new_n533_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n673_), .B1(new_n674_), .B2(new_n642_), .ZN(G1331gat));
  NOR2_X1   g474(.A1(new_n278_), .A2(new_n578_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n575_), .B1(new_n342_), .B2(new_n338_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n584_), .A2(new_n676_), .A3(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(G57gat), .B1(new_n679_), .B2(new_n622_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n586_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n681_), .A2(new_n677_), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n622_), .A2(G57gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n680_), .B1(new_n682_), .B2(new_n683_), .ZN(G1332gat));
  INV_X1    g483(.A(KEYINPUT48), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n682_), .A2(new_n647_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n685_), .B1(new_n686_), .B2(G64gat), .ZN(new_n687_));
  INV_X1    g486(.A(G64gat), .ZN(new_n688_));
  AOI211_X1 g487(.A(KEYINPUT48), .B(new_n688_), .C1(new_n682_), .C2(new_n647_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n647_), .A2(new_n688_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT112), .ZN(new_n691_));
  OAI22_X1  g490(.A1(new_n687_), .A2(new_n689_), .B1(new_n678_), .B2(new_n691_), .ZN(G1333gat));
  NOR2_X1   g491(.A1(new_n534_), .A2(G71gat), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT113), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n679_), .A2(new_n694_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n681_), .A2(new_n608_), .A3(new_n677_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT49), .ZN(new_n697_));
  AND3_X1   g496(.A1(new_n696_), .A2(new_n697_), .A3(G71gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n697_), .B1(new_n696_), .B2(G71gat), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n695_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT114), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  OAI211_X1 g501(.A(KEYINPUT114), .B(new_n695_), .C1(new_n698_), .C2(new_n699_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1334gat));
  OR3_X1    g503(.A1(new_n678_), .A2(G78gat), .A3(new_n551_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n682_), .A2(new_n533_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(G78gat), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n707_), .A2(KEYINPUT50), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n707_), .A2(KEYINPUT50), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n705_), .B1(new_n708_), .B2(new_n709_), .ZN(G1335gat));
  NAND2_X1  g509(.A1(new_n677_), .A2(new_n578_), .ZN(new_n711_));
  AOI211_X1 g510(.A(new_n585_), .B(new_n711_), .C1(new_n537_), .C2(new_n552_), .ZN(new_n712_));
  AOI21_X1  g511(.A(G85gat), .B1(new_n712_), .B2(new_n622_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT115), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n711_), .B(KEYINPUT116), .Z(new_n715_));
  AND2_X1   g514(.A1(new_n715_), .A2(new_n637_), .ZN(new_n716_));
  NAND4_X1  g515(.A1(new_n716_), .A2(new_n622_), .A3(new_n235_), .A4(new_n237_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n714_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT117), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n714_), .A2(KEYINPUT117), .A3(new_n717_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1336gat));
  AOI21_X1  g521(.A(G92gat), .B1(new_n712_), .B2(new_n599_), .ZN(new_n723_));
  AND3_X1   g522(.A1(new_n647_), .A2(new_n236_), .A3(new_n238_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n723_), .B1(new_n716_), .B2(new_n724_), .ZN(G1337gat));
  NAND3_X1  g524(.A1(new_n712_), .A2(new_n301_), .A3(new_n608_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n716_), .A2(new_n608_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n726_), .B1(new_n727_), .B2(new_n231_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT51), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n729_), .A2(KEYINPUT118), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(new_n731_));
  OAI221_X1 g530(.A(new_n726_), .B1(KEYINPUT118), .B2(new_n729_), .C1(new_n727_), .C2(new_n231_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(G1338gat));
  NAND3_X1  g532(.A1(new_n712_), .A2(new_n228_), .A3(new_n533_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n715_), .A2(new_n637_), .A3(new_n533_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT52), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n735_), .A2(new_n736_), .A3(G106gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n735_), .B2(G106gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n734_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(KEYINPUT53), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT53), .ZN(new_n741_));
  OAI211_X1 g540(.A(new_n741_), .B(new_n734_), .C1(new_n737_), .C2(new_n738_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(G1339gat));
  INV_X1    g542(.A(KEYINPUT55), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n294_), .A2(new_n281_), .A3(new_n311_), .ZN(new_n745_));
  AOI21_X1  g544(.A(KEYINPUT71), .B1(new_n316_), .B2(new_n319_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n744_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(KEYINPUT119), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n294_), .A2(new_n744_), .A3(new_n311_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n291_), .B1(new_n319_), .B2(new_n289_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT119), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n321_), .A2(new_n752_), .A3(new_n744_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n748_), .A2(new_n751_), .A3(new_n753_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(KEYINPUT120), .A2(KEYINPUT56), .ZN(new_n755_));
  AND3_X1   g554(.A1(new_n754_), .A2(new_n331_), .A3(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n754_), .B2(new_n331_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n336_), .A2(new_n575_), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n756_), .A2(new_n757_), .A3(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n564_), .A2(new_n559_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n554_), .A2(new_n557_), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n760_), .B(new_n569_), .C1(new_n761_), .C2(new_n559_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n571_), .A2(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n763_), .B1(new_n335_), .B2(new_n337_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n585_), .B1(new_n759_), .B2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT57), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT58), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n754_), .A2(new_n331_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT56), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n336_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n754_), .A2(new_n331_), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n571_), .B(new_n762_), .C1(new_n772_), .C2(KEYINPUT56), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n768_), .B1(new_n771_), .B2(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n763_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n334_), .B1(new_n772_), .B2(KEYINPUT56), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(KEYINPUT58), .A3(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n774_), .A2(new_n278_), .A3(new_n777_), .ZN(new_n778_));
  OAI211_X1 g577(.A(KEYINPUT57), .B(new_n585_), .C1(new_n759_), .C2(new_n764_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n767_), .A2(new_n778_), .A3(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT121), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n767_), .A2(new_n778_), .A3(KEYINPUT121), .A4(new_n779_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n782_), .A2(new_n578_), .A3(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT54), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n785_), .B1(new_n363_), .B2(new_n575_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n579_), .A2(KEYINPUT54), .A3(new_n576_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n784_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n532_), .A2(new_n622_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n790_), .A2(new_n575_), .A3(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(G113gat), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n576_), .A2(new_n794_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n791_), .A2(KEYINPUT59), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n780_), .A2(new_n578_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n797_), .B1(new_n798_), .B2(new_n788_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n791_), .B1(new_n784_), .B2(new_n789_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT59), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n796_), .B(new_n799_), .C1(new_n800_), .C2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n795_), .A2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(KEYINPUT122), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT122), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n795_), .A2(new_n802_), .A3(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n806_), .ZN(G1340gat));
  OAI211_X1 g606(.A(new_n577_), .B(new_n799_), .C1(new_n800_), .C2(new_n801_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n790_), .A2(new_n792_), .ZN(new_n809_));
  INV_X1    g608(.A(G120gat), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT60), .B1(new_n577_), .B2(new_n810_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n809_), .A2(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(G120gat), .B1(new_n808_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n812_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n813_), .B1(KEYINPUT60), .B2(new_n814_), .ZN(G1341gat));
  NAND3_X1  g614(.A1(new_n788_), .A2(new_n362_), .A3(new_n792_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT123), .ZN(new_n817_));
  INV_X1    g616(.A(G127gat), .ZN(new_n818_));
  AND3_X1   g617(.A1(new_n816_), .A2(new_n817_), .A3(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n817_), .B1(new_n816_), .B2(new_n818_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n799_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n821_), .B1(new_n809_), .B2(KEYINPUT59), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n578_), .A2(new_n818_), .ZN(new_n823_));
  AOI211_X1 g622(.A(new_n819_), .B(new_n820_), .C1(new_n822_), .C2(new_n823_), .ZN(G1342gat));
  INV_X1    g623(.A(new_n585_), .ZN(new_n825_));
  AOI21_X1  g624(.A(G134gat), .B1(new_n800_), .B2(new_n825_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(KEYINPUT124), .B(G134gat), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n279_), .A2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n826_), .B1(new_n822_), .B2(new_n828_), .ZN(G1343gat));
  NOR2_X1   g628(.A1(new_n551_), .A2(new_n608_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n831_), .B1(new_n784_), .B2(new_n789_), .ZN(new_n832_));
  XOR2_X1   g631(.A(new_n591_), .B(KEYINPUT109), .Z(new_n833_));
  NAND4_X1  g632(.A1(new_n832_), .A2(new_n622_), .A3(new_n575_), .A4(new_n833_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(G141gat), .ZN(G1344gat));
  NAND4_X1  g634(.A1(new_n832_), .A2(new_n622_), .A3(new_n577_), .A4(new_n833_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(KEYINPUT125), .B(G148gat), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n836_), .B(new_n837_), .ZN(G1345gat));
  NAND4_X1  g637(.A1(new_n832_), .A2(new_n622_), .A3(new_n362_), .A4(new_n833_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(KEYINPUT61), .B(G155gat), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n839_), .B(new_n840_), .ZN(G1346gat));
  NAND2_X1  g640(.A1(new_n790_), .A2(new_n830_), .ZN(new_n842_));
  NOR3_X1   g641(.A1(new_n842_), .A2(new_n411_), .A3(new_n647_), .ZN(new_n843_));
  INV_X1    g642(.A(G162gat), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n844_), .B1(new_n632_), .B2(new_n634_), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n832_), .A2(new_n622_), .A3(new_n825_), .A4(new_n833_), .ZN(new_n846_));
  AOI22_X1  g645(.A1(new_n843_), .A2(new_n845_), .B1(new_n844_), .B2(new_n846_), .ZN(G1347gat));
  NOR2_X1   g646(.A1(new_n798_), .A2(new_n788_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n833_), .A2(new_n622_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n625_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n848_), .A2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n575_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(G169gat), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT62), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n851_), .A2(new_n575_), .A3(new_n454_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n852_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n855_), .A2(new_n856_), .A3(new_n857_), .ZN(G1348gat));
  NAND2_X1  g657(.A1(new_n851_), .A2(new_n577_), .ZN(new_n859_));
  AND2_X1   g658(.A1(new_n859_), .A2(new_n450_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n850_), .B1(new_n784_), .B2(new_n789_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n861_), .A2(G176gat), .A3(new_n577_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT126), .ZN(new_n863_));
  AND2_X1   g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n862_), .A2(new_n863_), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n860_), .A2(new_n864_), .A3(new_n865_), .ZN(G1349gat));
  AOI21_X1  g665(.A(G183gat), .B1(new_n861_), .B2(new_n362_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n578_), .A2(new_n471_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n867_), .B1(new_n851_), .B2(new_n868_), .ZN(G1350gat));
  INV_X1    g668(.A(new_n851_), .ZN(new_n870_));
  OAI21_X1  g669(.A(G190gat), .B1(new_n870_), .B2(new_n279_), .ZN(new_n871_));
  OR2_X1    g670(.A1(new_n585_), .A2(new_n503_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n871_), .B1(new_n870_), .B2(new_n872_), .ZN(G1351gat));
  INV_X1    g672(.A(new_n849_), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n842_), .A2(new_n576_), .A3(new_n874_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(new_n416_), .ZN(G1352gat));
  NAND3_X1  g675(.A1(new_n832_), .A2(new_n577_), .A3(new_n849_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(G204gat), .ZN(G1353gat));
  NOR3_X1   g677(.A1(new_n842_), .A2(new_n578_), .A3(new_n874_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n880_));
  AND2_X1   g679(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n879_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n882_), .B1(new_n879_), .B2(new_n880_), .ZN(G1354gat));
  NOR2_X1   g682(.A1(new_n842_), .A2(new_n874_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n825_), .ZN(new_n885_));
  INV_X1    g684(.A(G218gat), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n279_), .A2(new_n886_), .ZN(new_n887_));
  AOI22_X1  g686(.A1(new_n885_), .A2(new_n886_), .B1(new_n884_), .B2(new_n887_), .ZN(G1355gat));
endmodule


