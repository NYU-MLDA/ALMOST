//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 1 0 0 0 1 0 1 1 0 0 1 1 0 1 0 0 0 0 0 1 0 0 0 0 1 1 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 1 0 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n707_, new_n708_, new_n709_,
    new_n711_, new_n712_, new_n713_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n855_, new_n856_, new_n857_,
    new_n859_, new_n860_, new_n861_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n896_, new_n898_, new_n899_, new_n900_,
    new_n901_, new_n903_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n918_;
  INV_X1    g000(.A(KEYINPUT12), .ZN(new_n202_));
  INV_X1    g001(.A(G85gat), .ZN(new_n203_));
  INV_X1    g002(.A(G92gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G85gat), .A2(G92gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n205_), .A2(KEYINPUT9), .A3(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT10), .B(G99gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n207_), .B1(new_n208_), .B2(G106gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT6), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT9), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n213_), .A2(G85gat), .A3(G92gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n212_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT64), .B1(new_n209_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n216_), .ZN(new_n218_));
  INV_X1    g017(.A(G106gat), .ZN(new_n219_));
  INV_X1    g018(.A(G99gat), .ZN(new_n220_));
  AND2_X1   g019(.A1(new_n220_), .A2(KEYINPUT10), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n220_), .A2(KEYINPUT10), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n219_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT64), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n218_), .A2(new_n223_), .A3(new_n224_), .A4(new_n207_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n217_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT7), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n227_), .A2(new_n220_), .A3(new_n219_), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n228_), .A2(new_n212_), .A3(new_n215_), .A4(new_n229_), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n205_), .A2(new_n206_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(KEYINPUT65), .A2(KEYINPUT8), .ZN(new_n232_));
  AND3_X1   g031(.A1(new_n230_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n232_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n226_), .A2(new_n235_), .ZN(new_n236_));
  OR2_X1    g035(.A1(G71gat), .A2(G78gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G71gat), .A2(G78gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G57gat), .A2(G64gat), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(G57gat), .A2(G64gat), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT11), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(G57gat), .ZN(new_n244_));
  INV_X1    g043(.A(G64gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT11), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n246_), .A2(new_n247_), .A3(new_n240_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n239_), .B1(new_n243_), .B2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n246_), .A2(new_n240_), .ZN(new_n250_));
  AOI22_X1  g049(.A1(new_n250_), .A2(KEYINPUT11), .B1(new_n237_), .B2(new_n238_), .ZN(new_n251_));
  OAI21_X1  g050(.A(KEYINPUT66), .B1(new_n249_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n239_), .ZN(new_n253_));
  NOR3_X1   g052(.A1(new_n241_), .A2(new_n242_), .A3(KEYINPUT11), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n247_), .B1(new_n246_), .B2(new_n240_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n253_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT66), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n243_), .A2(new_n239_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n256_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n252_), .A2(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n202_), .B1(new_n236_), .B2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G230gat), .A2(G233gat), .ZN(new_n262_));
  AND2_X1   g061(.A1(new_n217_), .A2(new_n225_), .ZN(new_n263_));
  OR2_X1    g062(.A1(new_n233_), .A2(new_n234_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n263_), .A2(new_n260_), .A3(new_n264_), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n217_), .B(new_n225_), .C1(new_n234_), .C2(new_n233_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n202_), .B1(new_n256_), .B2(new_n258_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n261_), .A2(new_n262_), .A3(new_n265_), .A4(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT67), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  AND2_X1   g070(.A1(new_n265_), .A2(new_n268_), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n272_), .A2(KEYINPUT67), .A3(new_n262_), .A4(new_n261_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n262_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n265_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n236_), .A2(new_n260_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n275_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n274_), .A2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G120gat), .B(G148gat), .ZN(new_n280_));
  INV_X1    g079(.A(G204gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT5), .ZN(new_n283_));
  INV_X1    g082(.A(G176gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n279_), .A2(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n274_), .A2(new_n278_), .A3(new_n285_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT13), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n287_), .B(new_n288_), .C1(KEYINPUT68), .C2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n287_), .A2(new_n288_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT68), .B(KEYINPUT13), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n290_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G29gat), .B(G36gat), .ZN(new_n295_));
  INV_X1    g094(.A(G43gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(G50gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n295_), .B(G43gat), .ZN(new_n299_));
  INV_X1    g098(.A(G50gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n298_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT15), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n298_), .A2(new_n301_), .A3(KEYINPUT15), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G15gat), .B(G22gat), .ZN(new_n307_));
  INV_X1    g106(.A(G1gat), .ZN(new_n308_));
  INV_X1    g107(.A(G8gat), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT14), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n307_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G1gat), .B(G8gat), .ZN(new_n312_));
  XOR2_X1   g111(.A(new_n311_), .B(new_n312_), .Z(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n306_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G229gat), .A2(G233gat), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n314_), .A2(new_n302_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n315_), .A2(new_n316_), .A3(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n302_), .B(new_n314_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n316_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n319_), .A2(new_n322_), .ZN(new_n323_));
  OR2_X1    g122(.A1(new_n323_), .A2(KEYINPUT72), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G113gat), .B(G141gat), .ZN(new_n325_));
  INV_X1    g124(.A(G169gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(G197gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n323_), .A2(KEYINPUT72), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n324_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n329_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n319_), .A2(new_n322_), .A3(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT73), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n319_), .A2(new_n322_), .A3(KEYINPUT73), .A4(new_n332_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n331_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n294_), .A2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G127gat), .B(G134gat), .ZN(new_n340_));
  INV_X1    g139(.A(G113gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(G120gat), .ZN(new_n343_));
  AND2_X1   g142(.A1(G155gat), .A2(G162gat), .ZN(new_n344_));
  NOR2_X1   g143(.A1(G155gat), .A2(G162gat), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(G141gat), .A2(G148gat), .ZN(new_n347_));
  XOR2_X1   g146(.A(new_n347_), .B(KEYINPUT3), .Z(new_n348_));
  NAND2_X1  g147(.A1(G141gat), .A2(G148gat), .ZN(new_n349_));
  XOR2_X1   g148(.A(new_n349_), .B(KEYINPUT2), .Z(new_n350_));
  OAI21_X1  g149(.A(new_n346_), .B1(new_n348_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT1), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n347_), .B1(new_n346_), .B2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n344_), .A2(KEYINPUT1), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n353_), .A2(new_n354_), .A3(new_n349_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n351_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n343_), .A2(new_n356_), .ZN(new_n357_));
  OR2_X1    g156(.A1(new_n357_), .A2(KEYINPUT4), .ZN(new_n358_));
  INV_X1    g157(.A(G120gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n342_), .B(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n360_), .A2(new_n355_), .A3(new_n351_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n361_), .A2(new_n357_), .A3(KEYINPUT4), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n358_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G225gat), .A2(G233gat), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT93), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n361_), .A2(new_n357_), .A3(new_n364_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT95), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT93), .ZN(new_n368_));
  INV_X1    g167(.A(new_n364_), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n358_), .A2(new_n362_), .A3(new_n368_), .A4(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n365_), .A2(new_n367_), .A3(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G1gat), .B(G29gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G57gat), .B(G85gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n372_), .B(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n375_));
  XOR2_X1   g174(.A(new_n374_), .B(new_n375_), .Z(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n371_), .A2(new_n377_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n365_), .A2(new_n367_), .A3(new_n376_), .A4(new_n370_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT27), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G211gat), .B(G218gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G197gat), .B(G204gat), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT21), .ZN(new_n385_));
  NOR3_X1   g184(.A1(new_n383_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n328_), .A2(G204gat), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n385_), .B1(new_n388_), .B2(KEYINPUT84), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(new_n384_), .ZN(new_n390_));
  AOI21_X1  g189(.A(KEYINPUT85), .B1(new_n390_), .B2(new_n383_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n389_), .A2(new_n384_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT84), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n281_), .A2(G197gat), .ZN(new_n394_));
  AND4_X1   g193(.A1(new_n393_), .A2(new_n388_), .A3(new_n394_), .A4(KEYINPUT21), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n383_), .B1(new_n392_), .B2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT85), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n387_), .B1(new_n391_), .B2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT76), .B(KEYINPUT23), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G183gat), .A2(G190gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n402_), .B1(KEYINPUT23), .B2(new_n401_), .ZN(new_n403_));
  INV_X1    g202(.A(G183gat), .ZN(new_n404_));
  INV_X1    g203(.A(G190gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  AND2_X1   g205(.A1(new_n403_), .A2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(KEYINPUT22), .B(G169gat), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT91), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n408_), .B(new_n409_), .ZN(new_n410_));
  XOR2_X1   g209(.A(KEYINPUT80), .B(G176gat), .Z(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G169gat), .A2(G176gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT92), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT92), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n412_), .A2(new_n416_), .A3(new_n413_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n407_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n418_));
  XOR2_X1   g217(.A(KEYINPUT89), .B(KEYINPUT24), .Z(new_n419_));
  NAND2_X1  g218(.A1(new_n326_), .A2(new_n284_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(new_n413_), .ZN(new_n421_));
  OR2_X1    g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n401_), .A2(KEYINPUT23), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n423_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(KEYINPUT25), .B(G183gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(KEYINPUT26), .B(G190gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n419_), .A2(new_n326_), .A3(new_n284_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n422_), .A2(new_n424_), .A3(new_n427_), .A4(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(KEYINPUT90), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n399_), .B1(new_n418_), .B2(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n403_), .B1(KEYINPUT24), .B2(new_n420_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(KEYINPUT77), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n420_), .A2(KEYINPUT24), .A3(new_n413_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(KEYINPUT74), .B(G190gat), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT26), .ZN(new_n436_));
  XOR2_X1   g235(.A(KEYINPUT75), .B(KEYINPUT26), .Z(new_n437_));
  OAI221_X1 g236(.A(new_n425_), .B1(new_n435_), .B2(new_n436_), .C1(new_n437_), .C2(new_n405_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT77), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n403_), .B(new_n439_), .C1(KEYINPUT24), .C2(new_n420_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n433_), .A2(new_n434_), .A3(new_n438_), .A4(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n424_), .B1(G183gat), .B2(new_n435_), .ZN(new_n442_));
  AND2_X1   g241(.A1(KEYINPUT78), .A2(G169gat), .ZN(new_n443_));
  NOR2_X1   g242(.A1(KEYINPUT78), .A2(G169gat), .ZN(new_n444_));
  OAI21_X1  g243(.A(KEYINPUT22), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n445_), .B(KEYINPUT79), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n411_), .B1(KEYINPUT22), .B2(new_n326_), .ZN(new_n447_));
  OAI211_X1 g246(.A(new_n442_), .B(new_n413_), .C1(new_n446_), .C2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n441_), .A2(new_n448_), .ZN(new_n449_));
  OAI211_X1 g248(.A(new_n431_), .B(KEYINPUT20), .C1(new_n399_), .C2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G226gat), .A2(G233gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(KEYINPUT19), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n452_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT20), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n455_), .B1(new_n449_), .B2(new_n399_), .ZN(new_n456_));
  OR2_X1    g255(.A1(new_n418_), .A2(new_n430_), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n454_), .B(new_n456_), .C1(new_n457_), .C2(new_n399_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(KEYINPUT18), .B(G64gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(G92gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G8gat), .B(G36gat), .ZN(new_n461_));
  XOR2_X1   g260(.A(new_n460_), .B(new_n461_), .Z(new_n462_));
  AND3_X1   g261(.A1(new_n453_), .A2(new_n458_), .A3(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n462_), .B1(new_n453_), .B2(new_n458_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n382_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n462_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n450_), .A2(new_n452_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n390_), .A2(KEYINPUT85), .A3(new_n383_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n396_), .A2(new_n397_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n386_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT86), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  AOI211_X1 g271(.A(KEYINPUT86), .B(new_n386_), .C1(new_n468_), .C2(new_n469_), .ZN(new_n473_));
  AND2_X1   g272(.A1(new_n415_), .A2(new_n417_), .ZN(new_n474_));
  OAI221_X1 g273(.A(new_n429_), .B1(new_n472_), .B2(new_n473_), .C1(new_n407_), .C2(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n454_), .B1(new_n475_), .B2(new_n456_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n466_), .B1(new_n467_), .B2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n453_), .A2(new_n458_), .A3(new_n462_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n477_), .A2(KEYINPUT27), .A3(new_n478_), .ZN(new_n479_));
  AND2_X1   g278(.A1(new_n465_), .A2(new_n479_), .ZN(new_n480_));
  XOR2_X1   g279(.A(G78gat), .B(G106gat), .Z(new_n481_));
  NAND2_X1  g280(.A1(new_n399_), .A2(KEYINPUT86), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT29), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n483_), .B1(new_n351_), .B2(new_n355_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n470_), .A2(new_n471_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n482_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G228gat), .A2(G233gat), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n488_), .B(KEYINPUT83), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NOR3_X1   g291(.A1(new_n470_), .A2(new_n484_), .A3(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n481_), .B1(new_n490_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n481_), .ZN(new_n496_));
  AOI211_X1 g295(.A(new_n496_), .B(new_n493_), .C1(new_n487_), .C2(new_n489_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT87), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n356_), .A2(KEYINPUT29), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G22gat), .B(G50gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT28), .ZN(new_n501_));
  AND2_X1   g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n499_), .A2(new_n501_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n498_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  NOR3_X1   g303(.A1(new_n495_), .A2(new_n497_), .A3(new_n504_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n472_), .A2(new_n473_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n488_), .B1(new_n506_), .B2(new_n485_), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n496_), .B(new_n504_), .C1(new_n507_), .C2(new_n493_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n502_), .A2(new_n503_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n490_), .A2(new_n481_), .A3(new_n494_), .A4(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  OAI21_X1  g310(.A(KEYINPUT88), .B1(new_n505_), .B2(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n496_), .B1(new_n507_), .B2(new_n493_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n490_), .A2(new_n481_), .A3(new_n494_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n504_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n513_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT88), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n516_), .A2(new_n517_), .A3(new_n510_), .A4(new_n508_), .ZN(new_n518_));
  AND3_X1   g317(.A1(new_n441_), .A2(KEYINPUT81), .A3(new_n448_), .ZN(new_n519_));
  AOI21_X1  g318(.A(KEYINPUT81), .B1(new_n441_), .B2(new_n448_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G227gat), .A2(G233gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT30), .ZN(new_n522_));
  XOR2_X1   g321(.A(G15gat), .B(G43gat), .Z(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  XOR2_X1   g323(.A(G71gat), .B(G99gat), .Z(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  OR3_X1    g326(.A1(new_n519_), .A2(new_n520_), .A3(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT82), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n527_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n528_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n360_), .B(KEYINPUT31), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n531_), .A2(new_n533_), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n528_), .A2(new_n529_), .A3(new_n530_), .A4(new_n532_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n512_), .A2(new_n518_), .A3(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n536_), .B1(new_n512_), .B2(new_n518_), .ZN(new_n538_));
  OAI211_X1 g337(.A(new_n381_), .B(new_n480_), .C1(new_n537_), .C2(new_n538_), .ZN(new_n539_));
  OAI211_X1 g338(.A(KEYINPUT32), .B(new_n462_), .C1(new_n467_), .C2(new_n476_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n462_), .A2(KEYINPUT32), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n453_), .A2(new_n458_), .A3(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n380_), .A2(new_n540_), .A3(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n453_), .A2(new_n458_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(new_n466_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n377_), .B1(new_n363_), .B2(new_n369_), .ZN(new_n546_));
  AND3_X1   g345(.A1(new_n361_), .A2(new_n357_), .A3(new_n369_), .ZN(new_n547_));
  OAI211_X1 g346(.A(new_n545_), .B(new_n478_), .C1(new_n546_), .C2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT33), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n379_), .B(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n543_), .B1(new_n548_), .B2(new_n550_), .ZN(new_n551_));
  AND2_X1   g350(.A1(new_n512_), .A2(new_n518_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n536_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n551_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n339_), .B1(new_n539_), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G231gat), .A2(G233gat), .ZN(new_n556_));
  XOR2_X1   g355(.A(new_n313_), .B(new_n556_), .Z(new_n557_));
  AND2_X1   g356(.A1(new_n252_), .A2(new_n259_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(KEYINPUT16), .B(G183gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(G211gat), .ZN(new_n561_));
  XOR2_X1   g360(.A(G127gat), .B(G155gat), .Z(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT17), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n563_), .A2(new_n564_), .ZN(new_n566_));
  NOR3_X1   g365(.A1(new_n559_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT71), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n256_), .A2(new_n258_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n557_), .B(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(new_n565_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n568_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n306_), .A2(new_n266_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(G232gat), .A2(G233gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT34), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(KEYINPUT35), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n575_), .A2(KEYINPUT35), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n266_), .A2(new_n302_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n573_), .A2(new_n576_), .A3(new_n577_), .A4(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n236_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n581_));
  OAI211_X1 g380(.A(KEYINPUT35), .B(new_n575_), .C1(new_n581_), .C2(new_n578_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n580_), .A2(new_n582_), .A3(KEYINPUT69), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G190gat), .B(G218gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(G134gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(G162gat), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n586_), .A2(KEYINPUT36), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n583_), .A2(new_n588_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n580_), .A2(new_n582_), .A3(KEYINPUT69), .A4(new_n587_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n580_), .A2(new_n582_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n592_), .A2(KEYINPUT36), .A3(new_n586_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n572_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n555_), .A2(new_n595_), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n596_), .B(KEYINPUT97), .Z(new_n597_));
  OAI21_X1  g396(.A(G1gat), .B1(new_n597_), .B2(new_n381_), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n598_), .B(KEYINPUT98), .Z(new_n599_));
  INV_X1    g398(.A(KEYINPUT70), .ZN(new_n600_));
  AND3_X1   g399(.A1(new_n591_), .A2(new_n600_), .A3(new_n593_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n600_), .B1(new_n591_), .B2(new_n593_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT37), .ZN(new_n603_));
  OR3_X1    g402(.A1(new_n601_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n603_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n572_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n555_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT38), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(KEYINPUT96), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n607_), .A2(new_n308_), .A3(new_n380_), .A4(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n608_), .A2(KEYINPUT96), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n599_), .A2(new_n612_), .ZN(G1324gat));
  INV_X1    g412(.A(new_n480_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n555_), .A2(new_n614_), .A3(new_n595_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(G8gat), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n616_), .A2(KEYINPUT39), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n616_), .A2(KEYINPUT39), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT99), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n607_), .A2(new_n309_), .A3(new_n614_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n619_), .A2(new_n620_), .A3(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT40), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n620_), .B1(new_n619_), .B2(new_n621_), .ZN(new_n625_));
  OR3_X1    g424(.A1(new_n623_), .A2(new_n624_), .A3(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n624_), .B1(new_n623_), .B2(new_n625_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(G1325gat));
  OAI21_X1  g427(.A(G15gat), .B1(new_n597_), .B2(new_n553_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n629_), .A2(KEYINPUT100), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n629_), .A2(KEYINPUT100), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT41), .ZN(new_n632_));
  OR3_X1    g431(.A1(new_n630_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(G15gat), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n607_), .A2(new_n634_), .A3(new_n536_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n632_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n633_), .A2(new_n635_), .A3(new_n636_), .ZN(G1326gat));
  OAI21_X1  g436(.A(G22gat), .B1(new_n597_), .B2(new_n552_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT42), .ZN(new_n639_));
  INV_X1    g438(.A(G22gat), .ZN(new_n640_));
  INV_X1    g439(.A(new_n552_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n607_), .A2(new_n640_), .A3(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n639_), .A2(new_n642_), .ZN(G1327gat));
  INV_X1    g442(.A(new_n572_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n339_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n539_), .A2(new_n554_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n604_), .A2(new_n605_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(KEYINPUT43), .B1(new_n649_), .B2(KEYINPUT101), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n647_), .B1(new_n539_), .B2(new_n554_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT101), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT43), .ZN(new_n653_));
  NOR3_X1   g452(.A1(new_n651_), .A2(new_n652_), .A3(new_n653_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n645_), .B1(new_n650_), .B2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT44), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  OAI211_X1 g456(.A(KEYINPUT44), .B(new_n645_), .C1(new_n650_), .C2(new_n654_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n657_), .A2(new_n380_), .A3(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(KEYINPUT102), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT102), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n657_), .A2(new_n661_), .A3(new_n380_), .A4(new_n658_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n660_), .A2(G29gat), .A3(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT103), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n660_), .A2(KEYINPUT103), .A3(G29gat), .A4(new_n662_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n572_), .A2(new_n594_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT104), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n555_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  OR3_X1    g470(.A1(new_n671_), .A2(G29gat), .A3(new_n381_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n667_), .A2(new_n672_), .ZN(G1328gat));
  INV_X1    g472(.A(KEYINPUT105), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT46), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n671_), .A2(G36gat), .A3(new_n480_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT45), .Z(new_n677_));
  NAND2_X1  g476(.A1(new_n657_), .A2(new_n658_), .ZN(new_n678_));
  OAI21_X1  g477(.A(G36gat), .B1(new_n678_), .B2(new_n480_), .ZN(new_n679_));
  AOI211_X1 g478(.A(new_n674_), .B(new_n675_), .C1(new_n677_), .C2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n674_), .A2(new_n675_), .ZN(new_n682_));
  AND4_X1   g481(.A1(new_n681_), .A2(new_n677_), .A3(new_n682_), .A4(new_n679_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n680_), .A2(new_n683_), .ZN(G1329gat));
  OAI21_X1  g483(.A(G43gat), .B1(new_n678_), .B2(new_n553_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n536_), .A2(new_n296_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n685_), .B1(new_n671_), .B2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT47), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n687_), .B(new_n688_), .ZN(G1330gat));
  OAI21_X1  g488(.A(G50gat), .B1(new_n678_), .B2(new_n552_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n670_), .A2(new_n300_), .A3(new_n641_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1331gat));
  INV_X1    g491(.A(new_n294_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n338_), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n646_), .A2(new_n693_), .A3(new_n694_), .A4(new_n595_), .ZN(new_n695_));
  NOR3_X1   g494(.A1(new_n695_), .A2(new_n244_), .A3(new_n381_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n338_), .B1(new_n539_), .B2(new_n554_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT106), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n698_), .A2(new_n693_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n699_), .A2(new_n380_), .A3(new_n606_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n696_), .B1(new_n700_), .B2(new_n244_), .ZN(G1332gat));
  OAI21_X1  g500(.A(G64gat), .B1(new_n695_), .B2(new_n480_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT48), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n699_), .A2(new_n606_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n614_), .A2(new_n245_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n703_), .B1(new_n704_), .B2(new_n705_), .ZN(G1333gat));
  OAI21_X1  g505(.A(G71gat), .B1(new_n695_), .B2(new_n553_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT49), .ZN(new_n708_));
  OR2_X1    g507(.A1(new_n553_), .A2(G71gat), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n708_), .B1(new_n704_), .B2(new_n709_), .ZN(G1334gat));
  OAI21_X1  g509(.A(G78gat), .B1(new_n695_), .B2(new_n552_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT50), .ZN(new_n712_));
  OR2_X1    g511(.A1(new_n552_), .A2(G78gat), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n712_), .B1(new_n704_), .B2(new_n713_), .ZN(G1335gat));
  OR2_X1    g513(.A1(new_n650_), .A2(new_n654_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n644_), .A2(new_n294_), .A3(new_n338_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  NOR3_X1   g516(.A1(new_n717_), .A2(new_n203_), .A3(new_n381_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n699_), .A2(new_n669_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(new_n380_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n718_), .B1(new_n720_), .B2(new_n203_), .ZN(G1336gat));
  NAND2_X1  g520(.A1(new_n699_), .A2(new_n669_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n204_), .B1(new_n722_), .B2(new_n480_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT107), .ZN(new_n724_));
  NOR3_X1   g523(.A1(new_n717_), .A2(new_n204_), .A3(new_n480_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n724_), .A2(new_n725_), .ZN(G1337gat));
  OAI21_X1  g525(.A(G99gat), .B1(new_n717_), .B2(new_n553_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n536_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n727_), .B1(new_n722_), .B2(new_n728_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g529(.A1(new_n719_), .A2(new_n219_), .A3(new_n641_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n715_), .A2(new_n641_), .A3(new_n716_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT52), .ZN(new_n733_));
  AND3_X1   g532(.A1(new_n732_), .A2(new_n733_), .A3(G106gat), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n732_), .B2(G106gat), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n731_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g536(.A1(new_n480_), .A2(new_n380_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n537_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT57), .ZN(new_n742_));
  XOR2_X1   g541(.A(KEYINPUT109), .B(KEYINPUT55), .Z(new_n743_));
  NAND2_X1  g542(.A1(new_n265_), .A2(new_n268_), .ZN(new_n744_));
  AOI21_X1  g543(.A(KEYINPUT12), .B1(new_n558_), .B2(new_n266_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(KEYINPUT67), .B1(new_n746_), .B2(new_n262_), .ZN(new_n747_));
  NOR4_X1   g546(.A1(new_n744_), .A2(new_n745_), .A3(new_n270_), .A4(new_n275_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n743_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT110), .ZN(new_n750_));
  OAI22_X1  g549(.A1(new_n744_), .A2(new_n745_), .B1(new_n750_), .B2(new_n262_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n262_), .A2(new_n750_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n261_), .A2(new_n265_), .A3(new_n268_), .A4(new_n752_), .ZN(new_n753_));
  OR2_X1    g552(.A1(new_n275_), .A2(KEYINPUT55), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n751_), .A2(new_n753_), .A3(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n749_), .A2(KEYINPUT111), .A3(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT111), .ZN(new_n757_));
  INV_X1    g556(.A(new_n743_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n758_), .B1(new_n271_), .B2(new_n273_), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n751_), .A2(new_n753_), .A3(new_n754_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n757_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n756_), .A2(new_n761_), .A3(KEYINPUT56), .A4(new_n286_), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n338_), .B(new_n288_), .C1(new_n762_), .C2(KEYINPUT112), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n756_), .A2(new_n761_), .A3(new_n286_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT56), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n767_), .A2(KEYINPUT112), .A3(new_n762_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT113), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n315_), .A2(new_n769_), .A3(new_n318_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n313_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n771_));
  OAI21_X1  g570(.A(KEYINPUT113), .B1(new_n771_), .B2(new_n317_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n770_), .A2(new_n321_), .A3(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n320_), .A2(new_n316_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  AOI22_X1  g574(.A1(new_n775_), .A2(new_n329_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n776_));
  AOI22_X1  g575(.A1(new_n764_), .A2(new_n768_), .B1(new_n291_), .B2(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n742_), .B1(new_n777_), .B2(new_n594_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n291_), .A2(new_n776_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n768_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n779_), .B1(new_n780_), .B2(new_n763_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n594_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n781_), .A2(KEYINPUT57), .A3(new_n782_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n778_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT115), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n767_), .A2(new_n762_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n776_), .A2(new_n288_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n789_), .A2(KEYINPUT114), .A3(KEYINPUT58), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT58), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n787_), .B1(new_n767_), .B2(new_n762_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n791_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  AOI211_X1 g593(.A(new_n785_), .B(new_n647_), .C1(new_n790_), .C2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n790_), .A2(new_n794_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n648_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(new_n785_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n784_), .A2(new_n796_), .A3(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n572_), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n647_), .A2(new_n294_), .A3(new_n694_), .A4(new_n644_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT108), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT108), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n606_), .A2(new_n804_), .A3(new_n294_), .A4(new_n694_), .ZN(new_n805_));
  AND3_X1   g604(.A1(new_n803_), .A2(KEYINPUT54), .A3(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT54), .B1(new_n803_), .B2(new_n805_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n741_), .B1(new_n801_), .B2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(G113gat), .B1(new_n809_), .B2(new_n338_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT59), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n740_), .A2(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n798_), .A2(new_n778_), .A3(new_n783_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n572_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n812_), .B1(new_n808_), .B2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n816_), .B1(new_n809_), .B2(new_n811_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n817_), .B1(KEYINPUT116), .B2(new_n341_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT116), .ZN(new_n819_));
  OAI21_X1  g618(.A(G113gat), .B1(new_n694_), .B2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n810_), .B1(new_n818_), .B2(new_n820_), .ZN(G1340gat));
  AOI21_X1  g620(.A(KEYINPUT115), .B1(new_n797_), .B2(new_n648_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n822_), .A2(new_n795_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n644_), .B1(new_n823_), .B2(new_n784_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n803_), .A2(new_n805_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n803_), .A2(KEYINPUT54), .A3(new_n805_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n740_), .B1(new_n824_), .B2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n815_), .B1(new_n830_), .B2(KEYINPUT59), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n359_), .B1(new_n831_), .B2(new_n693_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT60), .ZN(new_n833_));
  AOI21_X1  g632(.A(G120gat), .B1(new_n693_), .B2(new_n833_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n359_), .A2(KEYINPUT60), .ZN(new_n835_));
  NOR3_X1   g634(.A1(new_n830_), .A2(new_n834_), .A3(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(KEYINPUT117), .B1(new_n832_), .B2(new_n836_), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n816_), .B(new_n693_), .C1(new_n809_), .C2(new_n811_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(G120gat), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n840_));
  INV_X1    g639(.A(new_n836_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n839_), .A2(new_n840_), .A3(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n837_), .A2(new_n842_), .ZN(G1341gat));
  INV_X1    g642(.A(G127gat), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n844_), .B1(new_n830_), .B2(new_n572_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT118), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n845_), .B(new_n846_), .ZN(new_n847_));
  NOR3_X1   g646(.A1(new_n817_), .A2(new_n844_), .A3(new_n572_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n847_), .A2(new_n848_), .ZN(G1342gat));
  AOI21_X1  g648(.A(G134gat), .B1(new_n809_), .B2(new_n594_), .ZN(new_n850_));
  XOR2_X1   g649(.A(KEYINPUT119), .B(G134gat), .Z(new_n851_));
  NAND2_X1  g650(.A1(new_n648_), .A2(new_n851_), .ZN(new_n852_));
  XOR2_X1   g651(.A(new_n852_), .B(KEYINPUT120), .Z(new_n853_));
  AOI21_X1  g652(.A(new_n850_), .B1(new_n831_), .B2(new_n853_), .ZN(G1343gat));
  INV_X1    g653(.A(new_n538_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n855_), .B1(new_n801_), .B2(new_n808_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n856_), .A2(new_n380_), .A3(new_n338_), .A4(new_n480_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g657(.A(new_n856_), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n859_), .A2(new_n294_), .A3(new_n738_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(KEYINPUT121), .B(G148gat), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n860_), .B(new_n861_), .ZN(G1345gat));
  NOR3_X1   g661(.A1(new_n859_), .A2(new_n572_), .A3(new_n738_), .ZN(new_n863_));
  XOR2_X1   g662(.A(KEYINPUT61), .B(G155gat), .Z(new_n864_));
  XNOR2_X1  g663(.A(new_n863_), .B(new_n864_), .ZN(G1346gat));
  NOR2_X1   g664(.A1(new_n859_), .A2(new_n738_), .ZN(new_n866_));
  AOI21_X1  g665(.A(G162gat), .B1(new_n866_), .B2(new_n594_), .ZN(new_n867_));
  AND2_X1   g666(.A1(new_n648_), .A2(G162gat), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n867_), .B1(new_n866_), .B2(new_n868_), .ZN(G1347gat));
  NOR2_X1   g668(.A1(new_n480_), .A2(new_n380_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n871_), .A2(new_n739_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n873_), .B1(new_n808_), .B2(new_n814_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n875_), .A2(new_n694_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n876_), .A2(new_n326_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(KEYINPUT62), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT62), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n879_), .B1(new_n876_), .B2(new_n410_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n878_), .B1(new_n880_), .B2(new_n877_), .ZN(G1348gat));
  INV_X1    g680(.A(new_n411_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n882_), .B1(new_n874_), .B2(new_n693_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(KEYINPUT122), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n871_), .A2(new_n553_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n824_), .A2(new_n829_), .ZN(new_n887_));
  OAI21_X1  g686(.A(KEYINPUT123), .B1(new_n887_), .B2(new_n641_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n801_), .A2(new_n808_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT123), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n889_), .A2(new_n890_), .A3(new_n552_), .ZN(new_n891_));
  AOI211_X1 g690(.A(new_n284_), .B(new_n886_), .C1(new_n888_), .C2(new_n891_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n884_), .B1(new_n892_), .B2(new_n693_), .ZN(G1349gat));
  NOR3_X1   g692(.A1(new_n875_), .A2(new_n425_), .A3(new_n572_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n888_), .A2(new_n891_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n895_), .A2(new_n644_), .A3(new_n885_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n894_), .B1(new_n896_), .B2(new_n404_), .ZN(G1350gat));
  NAND3_X1  g696(.A1(new_n874_), .A2(new_n426_), .A3(new_n594_), .ZN(new_n898_));
  OAI21_X1  g697(.A(G190gat), .B1(new_n875_), .B2(new_n647_), .ZN(new_n899_));
  AND2_X1   g698(.A1(new_n899_), .A2(KEYINPUT124), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n899_), .A2(KEYINPUT124), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n898_), .B1(new_n900_), .B2(new_n901_), .ZN(G1351gat));
  NAND3_X1  g701(.A1(new_n856_), .A2(new_n338_), .A3(new_n870_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g703(.A1(new_n856_), .A2(new_n693_), .A3(new_n870_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(G204gat), .ZN(G1353gat));
  NAND4_X1  g705(.A1(new_n889_), .A2(new_n538_), .A3(new_n644_), .A4(new_n870_), .ZN(new_n907_));
  OR2_X1    g706(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT125), .ZN(new_n910_));
  XNOR2_X1  g709(.A(KEYINPUT63), .B(G211gat), .ZN(new_n911_));
  NAND4_X1  g710(.A1(new_n856_), .A2(new_n644_), .A3(new_n870_), .A4(new_n911_), .ZN(new_n912_));
  AND3_X1   g711(.A1(new_n909_), .A2(new_n910_), .A3(new_n912_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n910_), .B1(new_n909_), .B2(new_n912_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n913_), .A2(new_n914_), .ZN(G1354gat));
  XNOR2_X1  g714(.A(KEYINPUT126), .B(G218gat), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n859_), .A2(new_n871_), .A3(new_n916_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n856_), .A2(new_n594_), .A3(new_n870_), .ZN(new_n918_));
  AOI22_X1  g717(.A1(new_n917_), .A2(new_n648_), .B1(new_n918_), .B2(new_n916_), .ZN(G1355gat));
endmodule


