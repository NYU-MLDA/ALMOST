//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 1 0 0 1 0 1 1 1 1 0 0 0 1 0 1 0 0 1 1 0 1 0 0 1 0 0 0 1 0 1 1 0 0 0 1 0 0 1 0 1 1 0 1 1 0 1 0 1 1 1 0 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n736_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n759_, new_n760_, new_n761_, new_n762_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n786_, new_n787_, new_n789_, new_n790_, new_n791_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n893_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n934_, new_n935_, new_n937_,
    new_n938_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n954_, new_n955_, new_n956_;
  INV_X1    g000(.A(KEYINPUT99), .ZN(new_n202_));
  XOR2_X1   g001(.A(G8gat), .B(G36gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT18), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G64gat), .B(G92gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G226gat), .A2(G233gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT19), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT20), .ZN(new_n211_));
  NOR2_X1   g010(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(G169gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT23), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n214_), .B1(G183gat), .B2(G190gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G183gat), .A2(G190gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT82), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(KEYINPUT82), .A2(G183gat), .A3(G190gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n215_), .B1(new_n220_), .B2(new_n214_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(G183gat), .A2(G190gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n213_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  AOI21_X1  g022(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n224_), .B1(new_n220_), .B2(KEYINPUT23), .ZN(new_n225_));
  NOR3_X1   g024(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT25), .B(G183gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT26), .B(G190gat), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n226_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G169gat), .A2(G176gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT24), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT95), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(G169gat), .ZN(new_n234_));
  INV_X1    g033(.A(G176gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n230_), .A2(KEYINPUT95), .A3(KEYINPUT24), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n233_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n225_), .A2(new_n229_), .A3(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n223_), .A2(new_n239_), .ZN(new_n240_));
  OR2_X1    g039(.A1(G197gat), .A2(G204gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G197gat), .A2(G204gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT21), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n241_), .A2(KEYINPUT21), .A3(new_n242_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G211gat), .B(G218gat), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n245_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  OR2_X1    g047(.A1(new_n246_), .A2(new_n247_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n240_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT96), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n240_), .A2(KEYINPUT96), .A3(new_n250_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n211_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT78), .B(G183gat), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n225_), .B1(G190gat), .B2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(new_n213_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n250_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n236_), .A2(KEYINPUT24), .A3(new_n230_), .ZN(new_n260_));
  AND2_X1   g059(.A1(KEYINPUT79), .A2(KEYINPUT26), .ZN(new_n261_));
  NOR2_X1   g060(.A1(KEYINPUT79), .A2(KEYINPUT26), .ZN(new_n262_));
  OAI21_X1  g061(.A(G190gat), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT80), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT80), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n265_), .B(G190gat), .C1(new_n261_), .C2(new_n262_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(G190gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT26), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT25), .ZN(new_n270_));
  OR2_X1    g069(.A1(KEYINPUT78), .A2(G183gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(KEYINPUT78), .A2(G183gat), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n270_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n269_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  OAI211_X1 g074(.A(KEYINPUT81), .B(new_n260_), .C1(new_n267_), .C2(new_n275_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n221_), .A2(new_n226_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n256_), .A2(KEYINPUT25), .ZN(new_n279_));
  INV_X1    g078(.A(new_n274_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n281_), .A2(new_n269_), .A3(new_n264_), .A4(new_n266_), .ZN(new_n282_));
  AOI21_X1  g081(.A(KEYINPUT81), .B1(new_n282_), .B2(new_n260_), .ZN(new_n283_));
  OAI211_X1 g082(.A(new_n258_), .B(new_n259_), .C1(new_n278_), .C2(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n210_), .B1(new_n255_), .B2(new_n284_), .ZN(new_n285_));
  OAI211_X1 g084(.A(KEYINPUT20), .B(new_n210_), .C1(new_n240_), .C2(new_n250_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n258_), .B1(new_n278_), .B2(new_n283_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n286_), .B1(new_n287_), .B2(new_n250_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n207_), .B1(new_n285_), .B2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n284_), .ZN(new_n290_));
  AOI221_X4 g089(.A(new_n252_), .B1(new_n248_), .B2(new_n249_), .C1(new_n223_), .C2(new_n239_), .ZN(new_n291_));
  AOI21_X1  g090(.A(KEYINPUT96), .B1(new_n240_), .B2(new_n250_), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT20), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n209_), .B1(new_n290_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n288_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n294_), .A2(new_n206_), .A3(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT97), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G155gat), .A2(G162gat), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(G155gat), .A2(G162gat), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT88), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT3), .ZN(new_n303_));
  INV_X1    g102(.A(G141gat), .ZN(new_n304_));
  INV_X1    g103(.A(G148gat), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n303_), .A2(new_n304_), .A3(new_n305_), .A4(KEYINPUT87), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT87), .ZN(new_n307_));
  OAI22_X1  g106(.A1(new_n307_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n308_));
  AND2_X1   g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G141gat), .A2(G148gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT2), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT2), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n312_), .A2(G141gat), .A3(G148gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n311_), .A2(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n302_), .B1(new_n309_), .B2(new_n314_), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n314_), .A2(new_n302_), .A3(new_n308_), .A4(new_n306_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n301_), .B1(new_n315_), .B2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G113gat), .B(G120gat), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(G134gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(G127gat), .ZN(new_n322_));
  INV_X1    g121(.A(G127gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(G134gat), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n322_), .A2(new_n324_), .A3(KEYINPUT83), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(KEYINPUT83), .B1(new_n322_), .B2(new_n324_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n320_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n322_), .A2(new_n324_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT83), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n331_), .A2(new_n325_), .A3(new_n319_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n328_), .A2(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n300_), .B1(KEYINPUT1), .B2(new_n298_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n334_), .B1(KEYINPUT1), .B2(new_n298_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(G141gat), .A2(G148gat), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n335_), .A2(new_n310_), .A3(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n318_), .A2(new_n333_), .A3(new_n338_), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n328_), .A2(new_n332_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n301_), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n311_), .A2(new_n313_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n306_), .A2(new_n308_), .ZN(new_n343_));
  OAI21_X1  g142(.A(KEYINPUT88), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n341_), .B1(new_n344_), .B2(new_n316_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n338_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n340_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  AND3_X1   g146(.A1(new_n339_), .A2(new_n347_), .A3(KEYINPUT4), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT4), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n340_), .B(new_n349_), .C1(new_n345_), .C2(new_n346_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G225gat), .A2(G233gat), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n297_), .B1(new_n348_), .B2(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n339_), .A2(new_n347_), .A3(new_n351_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n339_), .A2(new_n347_), .A3(KEYINPUT4), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n356_), .A2(KEYINPUT97), .A3(new_n352_), .A4(new_n350_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G1gat), .B(G29gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(G85gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT0), .B(G57gat), .ZN(new_n360_));
  XOR2_X1   g159(.A(new_n359_), .B(new_n360_), .Z(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT33), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n354_), .A2(new_n355_), .A3(new_n357_), .A4(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n339_), .A2(new_n347_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT98), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n339_), .A2(new_n347_), .A3(KEYINPUT98), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n368_), .A2(new_n352_), .A3(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n356_), .A2(new_n351_), .A3(new_n350_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n370_), .A2(new_n371_), .A3(new_n362_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n289_), .A2(new_n296_), .A3(new_n365_), .A4(new_n372_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n354_), .A2(new_n355_), .A3(new_n361_), .A4(new_n357_), .ZN(new_n374_));
  AND2_X1   g173(.A1(new_n374_), .A2(new_n363_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n202_), .B1(new_n373_), .B2(new_n375_), .ZN(new_n376_));
  NOR3_X1   g175(.A1(new_n285_), .A2(new_n207_), .A3(new_n288_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n206_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n365_), .A2(new_n372_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n374_), .A2(new_n363_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n379_), .A2(new_n380_), .A3(KEYINPUT99), .A4(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n206_), .A2(KEYINPUT32), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n260_), .B1(new_n267_), .B2(new_n275_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT81), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n386_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n259_), .B1(new_n387_), .B2(new_n258_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT92), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n250_), .B(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT20), .B1(new_n390_), .B2(new_n240_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n209_), .B1(new_n388_), .B2(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n255_), .A2(new_n210_), .A3(new_n284_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n383_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n284_), .B(KEYINPUT20), .C1(new_n292_), .C2(new_n291_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n288_), .B1(new_n395_), .B2(new_n209_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n394_), .B1(new_n396_), .B2(new_n383_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n354_), .A2(new_n355_), .A3(new_n357_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(new_n362_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n374_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n397_), .A2(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n376_), .A2(new_n382_), .A3(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(KEYINPUT29), .B1(new_n345_), .B2(new_n346_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G228gat), .A2(G233gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(KEYINPUT90), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n250_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(KEYINPUT91), .B1(new_n403_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n403_), .A2(KEYINPUT91), .A3(new_n407_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n405_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n390_), .A2(new_n403_), .ZN(new_n412_));
  AOI22_X1  g211(.A1(new_n409_), .A2(new_n410_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G78gat), .B(G106gat), .ZN(new_n414_));
  XOR2_X1   g213(.A(new_n414_), .B(KEYINPUT93), .Z(new_n415_));
  NAND2_X1  g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n412_), .A2(new_n411_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n410_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n417_), .B1(new_n418_), .B2(new_n408_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n415_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n416_), .A2(new_n421_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n345_), .A2(new_n346_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT29), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(KEYINPUT28), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT28), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n423_), .A2(new_n427_), .A3(new_n424_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G22gat), .B(G50gat), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n426_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n429_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n427_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n432_));
  NOR4_X1   g231(.A1(new_n345_), .A2(new_n346_), .A3(KEYINPUT28), .A4(KEYINPUT29), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n431_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n430_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT89), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n430_), .A2(KEYINPUT89), .A3(new_n434_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n415_), .A2(KEYINPUT94), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n435_), .B1(new_n413_), .B2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n419_), .A2(new_n440_), .ZN(new_n443_));
  AOI22_X1  g242(.A1(new_n422_), .A2(new_n439_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n402_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT27), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n446_), .B1(new_n396_), .B2(new_n206_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n392_), .A2(new_n393_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(new_n207_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT100), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT100), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n447_), .A2(new_n452_), .A3(new_n449_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n451_), .A2(new_n453_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n444_), .A2(new_n400_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(KEYINPUT101), .B(KEYINPUT27), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n456_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n454_), .A2(new_n455_), .A3(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n445_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G227gat), .A2(G233gat), .ZN(new_n460_));
  INV_X1    g259(.A(G15gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n460_), .B(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(G43gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G71gat), .B(G99gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  OAI211_X1 g265(.A(KEYINPUT30), .B(new_n258_), .C1(new_n278_), .C2(new_n283_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(KEYINPUT30), .B1(new_n387_), .B2(new_n258_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n466_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT31), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n333_), .B(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT30), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n287_), .A2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n474_), .A2(new_n467_), .A3(new_n465_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n470_), .A2(new_n472_), .A3(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT85), .ZN(new_n477_));
  AND2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n470_), .A2(KEYINPUT85), .A3(new_n472_), .A4(new_n475_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT84), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n470_), .A2(new_n475_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n472_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n481_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  AOI211_X1 g283(.A(KEYINPUT84), .B(new_n472_), .C1(new_n470_), .C2(new_n475_), .ZN(new_n485_));
  OAI22_X1  g284(.A1(new_n478_), .A2(new_n480_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT86), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n474_), .A2(new_n467_), .A3(new_n465_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n465_), .B1(new_n474_), .B2(new_n467_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n483_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT84), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n482_), .A2(new_n481_), .A3(new_n483_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n476_), .A2(new_n477_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(new_n479_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n494_), .A2(KEYINPUT86), .A3(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n488_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n459_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n400_), .ZN(new_n501_));
  AND3_X1   g300(.A1(new_n494_), .A2(KEYINPUT86), .A3(new_n496_), .ZN(new_n502_));
  AOI21_X1  g301(.A(KEYINPUT86), .B1(new_n494_), .B2(new_n496_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n501_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT102), .ZN(new_n505_));
  INV_X1    g304(.A(new_n453_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n452_), .B1(new_n447_), .B2(new_n449_), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n444_), .B(new_n457_), .C1(new_n506_), .C2(new_n507_), .ZN(new_n508_));
  NOR3_X1   g307(.A1(new_n504_), .A2(new_n505_), .A3(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n400_), .B1(new_n488_), .B2(new_n497_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n508_), .ZN(new_n511_));
  AOI21_X1  g310(.A(KEYINPUT102), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n500_), .B1(new_n509_), .B2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(KEYINPUT65), .B(KEYINPUT6), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G99gat), .A2(G106gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(G85gat), .ZN(new_n517_));
  INV_X1    g316(.A(G92gat), .ZN(new_n518_));
  NOR3_X1   g317(.A1(new_n517_), .A2(new_n518_), .A3(KEYINPUT9), .ZN(new_n519_));
  XOR2_X1   g318(.A(G85gat), .B(G92gat), .Z(new_n520_));
  AOI21_X1  g319(.A(new_n519_), .B1(new_n520_), .B2(KEYINPUT9), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT10), .B(G99gat), .ZN(new_n522_));
  XOR2_X1   g321(.A(KEYINPUT64), .B(G106gat), .Z(new_n523_));
  OAI211_X1 g322(.A(new_n516_), .B(new_n521_), .C1(new_n522_), .C2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n525_));
  INV_X1    g324(.A(G99gat), .ZN(new_n526_));
  INV_X1    g325(.A(G106gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n516_), .A2(new_n525_), .A3(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT8), .ZN(new_n532_));
  AND3_X1   g331(.A1(new_n531_), .A2(new_n532_), .A3(new_n520_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n532_), .B1(new_n531_), .B2(new_n520_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n524_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G29gat), .B(G36gat), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT71), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G43gat), .B(G50gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  OR2_X1    g340(.A1(new_n535_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n540_), .B(KEYINPUT15), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(new_n535_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G232gat), .A2(G233gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT34), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n542_), .B(new_n544_), .C1(KEYINPUT35), .C2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n546_), .A2(KEYINPUT35), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n547_), .A2(KEYINPUT35), .A3(new_n546_), .ZN(new_n551_));
  XOR2_X1   g350(.A(G190gat), .B(G218gat), .Z(new_n552_));
  XNOR2_X1  g351(.A(G134gat), .B(G162gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT36), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT72), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n550_), .A2(new_n551_), .A3(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT73), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT37), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n554_), .B(KEYINPUT36), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n563_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n564_));
  NOR3_X1   g363(.A1(new_n560_), .A2(new_n561_), .A3(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n558_), .A2(new_n559_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n550_), .A2(new_n551_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n563_), .B1(new_n568_), .B2(KEYINPUT74), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n569_), .B1(KEYINPUT74), .B2(new_n568_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n570_), .A2(new_n558_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n567_), .B1(new_n571_), .B2(KEYINPUT37), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G57gat), .B(G64gat), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n573_), .A2(KEYINPUT11), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(KEYINPUT11), .ZN(new_n575_));
  XOR2_X1   g374(.A(G71gat), .B(G78gat), .Z(new_n576_));
  NAND3_X1  g375(.A1(new_n574_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n575_), .A2(new_n576_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G231gat), .A2(G233gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G15gat), .B(G22gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(KEYINPUT75), .B(G1gat), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n583_), .A2(G8gat), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT14), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n582_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G1gat), .B(G8gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n581_), .B(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  XOR2_X1   g389(.A(G127gat), .B(G155gat), .Z(new_n591_));
  XNOR2_X1  g390(.A(G183gat), .B(G211gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  XOR2_X1   g392(.A(KEYINPUT76), .B(KEYINPUT16), .Z(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n595_), .A2(KEYINPUT17), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n595_), .A2(KEYINPUT17), .ZN(new_n597_));
  NOR3_X1   g396(.A1(new_n590_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(KEYINPUT77), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n590_), .A2(new_n596_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n598_), .A2(KEYINPUT77), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n572_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n543_), .A2(new_n588_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(G229gat), .A2(G233gat), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n588_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n608_), .B1(new_n609_), .B2(new_n540_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n540_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n541_), .A2(new_n588_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  AOI22_X1  g412(.A1(new_n606_), .A2(new_n610_), .B1(new_n613_), .B2(new_n608_), .ZN(new_n614_));
  XOR2_X1   g413(.A(G113gat), .B(G141gat), .Z(new_n615_));
  XNOR2_X1  g414(.A(G169gat), .B(G197gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n614_), .B(new_n617_), .ZN(new_n618_));
  XOR2_X1   g417(.A(G120gat), .B(G148gat), .Z(new_n619_));
  XNOR2_X1  g418(.A(G176gat), .B(G204gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(G230gat), .A2(G233gat), .ZN(new_n625_));
  INV_X1    g424(.A(new_n579_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n535_), .A2(new_n626_), .ZN(new_n627_));
  OAI211_X1 g426(.A(new_n579_), .B(new_n524_), .C1(new_n533_), .C2(new_n534_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n625_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n629_), .A2(KEYINPUT67), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n627_), .A2(new_n628_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n625_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n631_), .A2(KEYINPUT67), .A3(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n630_), .A2(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(KEYINPUT68), .B1(new_n535_), .B2(new_n626_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT12), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n628_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  AOI211_X1 g436(.A(KEYINPUT68), .B(KEYINPUT12), .C1(new_n535_), .C2(new_n626_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n637_), .A2(new_n632_), .A3(new_n638_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n624_), .B1(new_n634_), .B2(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n637_), .A2(new_n638_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(new_n625_), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n642_), .A2(new_n633_), .A3(new_n630_), .A4(new_n623_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n640_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT70), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n644_), .B1(new_n645_), .B2(KEYINPUT13), .ZN(new_n646_));
  XOR2_X1   g445(.A(KEYINPUT70), .B(KEYINPUT13), .Z(new_n647_));
  NAND3_X1  g446(.A1(new_n640_), .A2(new_n643_), .A3(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  AND4_X1   g448(.A1(new_n513_), .A2(new_n605_), .A3(new_n618_), .A4(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n501_), .A2(new_n583_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n652_), .A2(KEYINPUT38), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(KEYINPUT38), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n498_), .B1(new_n445_), .B2(new_n458_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n505_), .B1(new_n504_), .B2(new_n508_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n510_), .A2(new_n511_), .A3(KEYINPUT102), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n655_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n658_), .A2(new_n571_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n649_), .A2(new_n618_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n660_), .A2(new_n604_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n659_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(G1gat), .B1(new_n663_), .B2(new_n501_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n653_), .A2(new_n654_), .A3(new_n664_), .ZN(G1324gat));
  NAND2_X1  g464(.A1(new_n454_), .A2(new_n457_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n662_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(G8gat), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n668_), .B1(KEYINPUT103), .B2(KEYINPUT39), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(KEYINPUT103), .A2(KEYINPUT39), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n670_), .B(new_n671_), .Z(new_n672_));
  NAND3_X1  g471(.A1(new_n650_), .A2(new_n668_), .A3(new_n666_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n674_), .B(KEYINPUT40), .Z(G1325gat));
  AOI21_X1  g474(.A(new_n461_), .B1(new_n662_), .B2(new_n498_), .ZN(new_n676_));
  XOR2_X1   g475(.A(KEYINPUT104), .B(KEYINPUT41), .Z(new_n677_));
  OR2_X1    g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n650_), .A2(new_n461_), .A3(new_n498_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n676_), .A2(new_n677_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n678_), .A2(new_n679_), .A3(new_n680_), .ZN(G1326gat));
  INV_X1    g480(.A(G22gat), .ZN(new_n682_));
  INV_X1    g481(.A(new_n444_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n682_), .B1(new_n662_), .B2(new_n683_), .ZN(new_n684_));
  XOR2_X1   g483(.A(new_n684_), .B(KEYINPUT42), .Z(new_n685_));
  NAND3_X1  g484(.A1(new_n650_), .A2(new_n682_), .A3(new_n683_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(G1327gat));
  NOR2_X1   g486(.A1(new_n660_), .A2(new_n603_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT43), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n689_), .B1(new_n513_), .B2(new_n572_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n570_), .A2(new_n558_), .ZN(new_n691_));
  AOI22_X1  g490(.A1(new_n691_), .A2(new_n561_), .B1(new_n566_), .B2(new_n565_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n658_), .A2(KEYINPUT43), .A3(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n688_), .B1(new_n690_), .B2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  OAI211_X1 g495(.A(KEYINPUT44), .B(new_n688_), .C1(new_n690_), .C2(new_n693_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  OAI21_X1  g497(.A(G29gat), .B1(new_n698_), .B2(new_n501_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n571_), .A2(new_n604_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT105), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n701_), .A2(new_n513_), .A3(new_n618_), .A4(new_n649_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT106), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n702_), .B(new_n703_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n501_), .A2(G29gat), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT107), .Z(new_n706_));
  OAI21_X1  g505(.A(new_n699_), .B1(new_n704_), .B2(new_n706_), .ZN(G1328gat));
  XNOR2_X1  g506(.A(new_n666_), .B(KEYINPUT110), .ZN(new_n708_));
  INV_X1    g507(.A(G36gat), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(KEYINPUT45), .B1(new_n704_), .B2(new_n710_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n702_), .B(KEYINPUT106), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT45), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n712_), .A2(new_n713_), .A3(new_n709_), .A4(new_n708_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT46), .ZN(new_n715_));
  AOI22_X1  g514(.A1(new_n711_), .A2(new_n714_), .B1(KEYINPUT111), .B2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT109), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT108), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n696_), .A2(new_n718_), .A3(new_n697_), .A4(new_n666_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n719_), .A2(G36gat), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n696_), .A2(new_n666_), .A3(new_n697_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(KEYINPUT108), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n717_), .B1(new_n720_), .B2(new_n722_), .ZN(new_n723_));
  AND4_X1   g522(.A1(new_n717_), .A2(new_n722_), .A3(G36gat), .A4(new_n719_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n716_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n715_), .A2(KEYINPUT111), .ZN(new_n726_));
  XOR2_X1   g525(.A(new_n726_), .B(KEYINPUT112), .Z(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n725_), .A2(new_n728_), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n716_), .B(new_n727_), .C1(new_n723_), .C2(new_n724_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1329gat));
  OAI21_X1  g530(.A(G43gat), .B1(new_n698_), .B2(new_n499_), .ZN(new_n732_));
  OR2_X1    g531(.A1(new_n499_), .A2(G43gat), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n704_), .B2(new_n733_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g534(.A(G50gat), .B1(new_n712_), .B2(new_n683_), .ZN(new_n736_));
  INV_X1    g535(.A(G50gat), .ZN(new_n737_));
  NOR3_X1   g536(.A1(new_n698_), .A2(new_n737_), .A3(new_n444_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n736_), .A2(new_n738_), .ZN(G1331gat));
  NOR2_X1   g538(.A1(new_n658_), .A2(new_n618_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n649_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n740_), .A2(new_n605_), .A3(new_n741_), .ZN(new_n742_));
  XOR2_X1   g541(.A(new_n742_), .B(KEYINPUT113), .Z(new_n743_));
  INV_X1    g542(.A(G57gat), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n743_), .A2(new_n744_), .A3(new_n400_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n618_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n741_), .A2(new_n746_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n747_), .A2(new_n604_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n659_), .A2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  OAI21_X1  g549(.A(G57gat), .B1(new_n750_), .B2(new_n501_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n745_), .A2(new_n751_), .ZN(G1332gat));
  INV_X1    g551(.A(G64gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n749_), .B2(new_n708_), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT48), .Z(new_n755_));
  NAND3_X1  g554(.A1(new_n743_), .A2(new_n753_), .A3(new_n708_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  XOR2_X1   g556(.A(new_n757_), .B(KEYINPUT114), .Z(G1333gat));
  INV_X1    g557(.A(G71gat), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n759_), .B1(new_n749_), .B2(new_n498_), .ZN(new_n760_));
  XOR2_X1   g559(.A(new_n760_), .B(KEYINPUT49), .Z(new_n761_));
  NAND3_X1  g560(.A1(new_n743_), .A2(new_n759_), .A3(new_n498_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(G1334gat));
  NAND2_X1  g562(.A1(new_n749_), .A2(new_n683_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(G78gat), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT115), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT115), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n764_), .A2(new_n767_), .A3(G78gat), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT50), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(G78gat), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n743_), .A2(new_n772_), .A3(new_n683_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n766_), .A2(KEYINPUT50), .A3(new_n768_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n771_), .A2(new_n773_), .A3(new_n774_), .ZN(new_n775_));
  XOR2_X1   g574(.A(new_n775_), .B(KEYINPUT116), .Z(G1335gat));
  AND2_X1   g575(.A1(new_n701_), .A2(new_n741_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(new_n740_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n779_), .A2(new_n517_), .A3(new_n400_), .ZN(new_n780_));
  OAI21_X1  g579(.A(KEYINPUT43), .B1(new_n658_), .B2(new_n692_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n513_), .A2(new_n689_), .A3(new_n572_), .ZN(new_n782_));
  AOI211_X1 g581(.A(new_n603_), .B(new_n747_), .C1(new_n781_), .C2(new_n782_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n783_), .A2(new_n400_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n780_), .B1(new_n517_), .B2(new_n784_), .ZN(G1336gat));
  NAND3_X1  g584(.A1(new_n779_), .A2(new_n518_), .A3(new_n666_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n783_), .A2(new_n708_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n786_), .B1(new_n787_), .B2(new_n518_), .ZN(G1337gat));
  AOI21_X1  g587(.A(new_n526_), .B1(new_n783_), .B2(new_n498_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n499_), .A2(new_n522_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n789_), .B1(new_n779_), .B2(new_n790_), .ZN(new_n791_));
  XOR2_X1   g590(.A(new_n791_), .B(KEYINPUT51), .Z(G1338gat));
  AOI21_X1  g591(.A(new_n527_), .B1(new_n783_), .B2(new_n683_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT52), .ZN(new_n794_));
  NOR3_X1   g593(.A1(new_n778_), .A2(new_n444_), .A3(new_n523_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  XOR2_X1   g595(.A(KEYINPUT117), .B(KEYINPUT53), .Z(new_n797_));
  XNOR2_X1  g596(.A(new_n796_), .B(new_n797_), .ZN(G1339gat));
  NAND3_X1  g597(.A1(new_n605_), .A2(new_n746_), .A3(new_n649_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT54), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n799_), .B(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n643_), .A2(new_n618_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT56), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n632_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(KEYINPUT55), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(new_n642_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n641_), .A2(KEYINPUT55), .A3(new_n625_), .ZN(new_n807_));
  AOI211_X1 g606(.A(new_n803_), .B(new_n623_), .C1(new_n806_), .C2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT118), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n802_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n639_), .B1(KEYINPUT55), .B2(new_n804_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n807_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n624_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n803_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n806_), .A2(new_n807_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n815_), .A2(KEYINPUT56), .A3(new_n624_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n814_), .A2(KEYINPUT118), .A3(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n810_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT119), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n810_), .A2(new_n817_), .A3(KEYINPUT119), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n606_), .A2(new_n611_), .A3(new_n608_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n617_), .B1(new_n613_), .B2(new_n607_), .ZN(new_n823_));
  AOI22_X1  g622(.A1(new_n614_), .A2(new_n617_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n644_), .A2(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n820_), .A2(new_n821_), .A3(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n691_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT120), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT57), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n827_), .A2(new_n828_), .A3(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n825_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n831_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n571_), .B1(new_n832_), .B2(new_n821_), .ZN(new_n833_));
  OAI21_X1  g632(.A(KEYINPUT120), .B1(new_n833_), .B2(KEYINPUT57), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n643_), .A2(new_n824_), .ZN(new_n835_));
  AOI21_X1  g634(.A(KEYINPUT56), .B1(new_n815_), .B2(new_n624_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n835_), .B1(new_n836_), .B2(KEYINPUT121), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT121), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n814_), .A2(new_n838_), .A3(new_n816_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT58), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n837_), .A2(KEYINPUT58), .A3(new_n839_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n842_), .A2(new_n843_), .A3(new_n572_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(KEYINPUT122), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT122), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n842_), .A2(new_n843_), .A3(new_n572_), .A4(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n833_), .A2(KEYINPUT57), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n830_), .A2(new_n834_), .A3(new_n848_), .A4(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n801_), .B1(new_n850_), .B2(new_n604_), .ZN(new_n851_));
  NOR3_X1   g650(.A1(new_n499_), .A2(new_n501_), .A3(new_n508_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(KEYINPUT59), .B1(new_n851_), .B2(new_n853_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n853_), .A2(KEYINPUT59), .ZN(new_n855_));
  AOI211_X1 g654(.A(new_n829_), .B(new_n571_), .C1(new_n832_), .C2(new_n821_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n844_), .B1(new_n833_), .B2(KEYINPUT57), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT123), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n856_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  OAI211_X1 g658(.A(KEYINPUT123), .B(new_n844_), .C1(new_n833_), .C2(KEYINPUT57), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n603_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n855_), .B1(new_n861_), .B2(new_n801_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n854_), .A2(new_n862_), .ZN(new_n863_));
  OAI21_X1  g662(.A(G113gat), .B1(new_n863_), .B2(new_n746_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n850_), .A2(new_n604_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n801_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n852_), .ZN(new_n868_));
  OR2_X1    g667(.A1(new_n746_), .A2(G113gat), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n864_), .B1(new_n868_), .B2(new_n869_), .ZN(G1340gat));
  OAI21_X1  g669(.A(G120gat), .B1(new_n863_), .B2(new_n649_), .ZN(new_n871_));
  INV_X1    g670(.A(G120gat), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n872_), .B1(new_n649_), .B2(KEYINPUT60), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n873_), .B1(KEYINPUT60), .B2(new_n872_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n871_), .B1(new_n868_), .B2(new_n874_), .ZN(G1341gat));
  OAI21_X1  g674(.A(G127gat), .B1(new_n863_), .B2(new_n604_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n851_), .A2(new_n853_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n877_), .A2(new_n323_), .A3(new_n603_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n878_), .ZN(G1342gat));
  INV_X1    g678(.A(KEYINPUT124), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n692_), .A2(new_n321_), .ZN(new_n881_));
  AND3_X1   g680(.A1(new_n854_), .A2(new_n862_), .A3(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(G134gat), .B1(new_n877_), .B2(new_n571_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n880_), .B1(new_n882_), .B2(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n321_), .B1(new_n868_), .B2(new_n691_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n881_), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n885_), .B(KEYINPUT124), .C1(new_n863_), .C2(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n884_), .A2(new_n887_), .ZN(G1343gat));
  NOR3_X1   g687(.A1(new_n851_), .A2(new_n498_), .A3(new_n444_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n708_), .A2(new_n501_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n889_), .A2(new_n618_), .A3(new_n890_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g691(.A1(new_n889_), .A2(new_n741_), .A3(new_n890_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g693(.A1(new_n889_), .A2(new_n603_), .A3(new_n890_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(KEYINPUT61), .B(G155gat), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n895_), .B(new_n896_), .ZN(G1346gat));
  INV_X1    g696(.A(G162gat), .ZN(new_n898_));
  NAND4_X1  g697(.A1(new_n889_), .A2(new_n898_), .A3(new_n571_), .A4(new_n890_), .ZN(new_n899_));
  AND3_X1   g698(.A1(new_n889_), .A2(new_n572_), .A3(new_n890_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n899_), .B1(new_n900_), .B2(new_n898_), .ZN(G1347gat));
  NAND2_X1  g700(.A1(new_n708_), .A2(new_n501_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n902_), .A2(new_n499_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n903_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n904_), .A2(new_n683_), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n618_), .B(new_n905_), .C1(new_n861_), .C2(new_n801_), .ZN(new_n906_));
  OAI211_X1 g705(.A(KEYINPUT62), .B(new_n234_), .C1(new_n906_), .C2(KEYINPUT22), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT62), .ZN(new_n908_));
  AOI21_X1  g707(.A(KEYINPUT57), .B1(new_n826_), .B2(new_n691_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n844_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n858_), .B1(new_n909_), .B2(new_n910_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n911_), .A2(new_n849_), .A3(new_n860_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n801_), .B1(new_n912_), .B2(new_n604_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n905_), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n913_), .A2(new_n746_), .A3(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT22), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n908_), .B1(new_n915_), .B2(new_n916_), .ZN(new_n917_));
  OAI21_X1  g716(.A(G169gat), .B1(new_n906_), .B2(KEYINPUT62), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n907_), .B1(new_n917_), .B2(new_n918_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n919_), .ZN(G1348gat));
  NOR2_X1   g719(.A1(new_n913_), .A2(new_n914_), .ZN(new_n921_));
  AOI21_X1  g720(.A(G176gat), .B1(new_n921_), .B2(new_n741_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n851_), .A2(new_n683_), .ZN(new_n923_));
  NOR3_X1   g722(.A1(new_n904_), .A2(new_n235_), .A3(new_n649_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n922_), .B1(new_n923_), .B2(new_n924_), .ZN(G1349gat));
  NAND3_X1  g724(.A1(new_n923_), .A2(new_n603_), .A3(new_n903_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n926_), .A2(new_n271_), .A3(new_n272_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT125), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n604_), .A2(new_n227_), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n921_), .A2(new_n928_), .A3(new_n929_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n921_), .A2(new_n929_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n931_), .A2(KEYINPUT125), .ZN(new_n932_));
  AND3_X1   g731(.A1(new_n927_), .A2(new_n930_), .A3(new_n932_), .ZN(G1350gat));
  NAND3_X1  g732(.A1(new_n921_), .A2(new_n228_), .A3(new_n571_), .ZN(new_n934_));
  NOR3_X1   g733(.A1(new_n913_), .A2(new_n692_), .A3(new_n914_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n934_), .B1(new_n268_), .B2(new_n935_), .ZN(G1351gat));
  NOR4_X1   g735(.A1(new_n851_), .A2(new_n498_), .A3(new_n444_), .A4(new_n902_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n937_), .A2(new_n618_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g738(.A(KEYINPUT126), .ZN(new_n940_));
  AND2_X1   g739(.A1(new_n940_), .A2(G204gat), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n940_), .A2(G204gat), .ZN(new_n942_));
  OAI211_X1 g741(.A(new_n937_), .B(new_n741_), .C1(new_n941_), .C2(new_n942_), .ZN(new_n943_));
  INV_X1    g742(.A(new_n937_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n944_), .A2(new_n649_), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n943_), .B1(new_n945_), .B2(new_n942_), .ZN(G1353gat));
  INV_X1    g745(.A(KEYINPUT63), .ZN(new_n947_));
  INV_X1    g746(.A(G211gat), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n603_), .B1(new_n947_), .B2(new_n948_), .ZN(new_n949_));
  XOR2_X1   g748(.A(new_n949_), .B(KEYINPUT127), .Z(new_n950_));
  NAND2_X1  g749(.A1(new_n937_), .A2(new_n950_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n947_), .A2(new_n948_), .ZN(new_n952_));
  XNOR2_X1  g751(.A(new_n951_), .B(new_n952_), .ZN(G1354gat));
  OAI21_X1  g752(.A(G218gat), .B1(new_n944_), .B2(new_n692_), .ZN(new_n954_));
  INV_X1    g753(.A(G218gat), .ZN(new_n955_));
  NAND3_X1  g754(.A1(new_n937_), .A2(new_n955_), .A3(new_n571_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n954_), .A2(new_n956_), .ZN(G1355gat));
endmodule


